magic
tech sky130B
magscale 1 2
timestamp 1716986954
<< metal1 >>
rect 485038 700272 485044 700324
rect 485096 700312 485102 700324
rect 527174 700312 527180 700324
rect 485096 700284 527180 700312
rect 485096 700272 485102 700284
rect 527174 700272 527180 700284
rect 527232 700272 527238 700324
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 87598 683176 87604 683188
rect 3476 683148 87604 683176
rect 3476 683136 3482 683148
rect 87598 683136 87604 683148
rect 87656 683136 87662 683188
rect 487798 657500 487804 657552
rect 487856 657540 487862 657552
rect 534902 657540 534908 657552
rect 487856 657512 534908 657540
rect 487856 657500 487862 657512
rect 534902 657500 534908 657512
rect 534960 657500 534966 657552
rect 487890 657432 487896 657484
rect 487948 657472 487954 657484
rect 537662 657472 537668 657484
rect 487948 657444 537668 657472
rect 487948 657432 487954 657444
rect 537662 657432 537668 657444
rect 537720 657432 537726 657484
rect 486878 657364 486884 657416
rect 486936 657404 486942 657416
rect 496262 657404 496268 657416
rect 486936 657376 496268 657404
rect 486936 657364 486942 657376
rect 496262 657364 496268 657376
rect 496320 657364 496326 657416
rect 503162 657364 503168 657416
rect 503220 657404 503226 657416
rect 580442 657404 580448 657416
rect 503220 657376 580448 657404
rect 503220 657364 503226 657376
rect 580442 657364 580448 657376
rect 580500 657364 580506 657416
rect 487154 657296 487160 657348
rect 487212 657336 487218 657348
rect 497642 657336 497648 657348
rect 487212 657308 497648 657336
rect 487212 657296 487218 657308
rect 497642 657296 497648 657308
rect 497700 657296 497706 657348
rect 505094 657296 505100 657348
rect 505152 657336 505158 657348
rect 530762 657336 530768 657348
rect 505152 657308 530768 657336
rect 505152 657296 505158 657308
rect 530762 657296 530768 657308
rect 530820 657296 530826 657348
rect 490374 657228 490380 657280
rect 490432 657268 490438 657280
rect 529382 657268 529388 657280
rect 490432 657240 529388 657268
rect 490432 657228 490438 657240
rect 529382 657228 529388 657240
rect 529440 657228 529446 657280
rect 490466 657160 490472 657212
rect 490524 657200 490530 657212
rect 533522 657200 533528 657212
rect 490524 657172 533528 657200
rect 490524 657160 490530 657172
rect 533522 657160 533528 657172
rect 533580 657160 533586 657212
rect 489178 657092 489184 657144
rect 489236 657132 489242 657144
rect 532142 657132 532148 657144
rect 489236 657104 532148 657132
rect 489236 657092 489242 657104
rect 532142 657092 532148 657104
rect 532200 657092 532206 657144
rect 488442 657024 488448 657076
rect 488500 657064 488506 657076
rect 494882 657064 494888 657076
rect 488500 657036 494888 657064
rect 488500 657024 488506 657036
rect 494882 657024 494888 657036
rect 494940 657024 494946 657076
rect 487062 656956 487068 657008
rect 487120 656996 487126 657008
rect 493502 656996 493508 657008
rect 487120 656968 493508 656996
rect 487120 656956 487126 656968
rect 493502 656956 493508 656968
rect 493560 656956 493566 657008
rect 486970 656888 486976 656940
rect 487028 656928 487034 656940
rect 492122 656928 492128 656940
rect 487028 656900 492128 656928
rect 487028 656888 487034 656900
rect 492122 656888 492128 656900
rect 492180 656888 492186 656940
rect 494698 656888 494704 656940
rect 494756 656928 494762 656940
rect 504542 656928 504548 656940
rect 494756 656900 504548 656928
rect 494756 656888 494762 656900
rect 504542 656888 504548 656900
rect 504600 656888 504606 656940
rect 514754 656888 514760 656940
rect 514812 656928 514818 656940
rect 526622 656928 526628 656940
rect 514812 656900 526628 656928
rect 514812 656888 514818 656900
rect 526622 656888 526628 656900
rect 526680 656888 526686 656940
rect 224954 656140 224960 656192
rect 225012 656180 225018 656192
rect 503162 656180 503168 656192
rect 225012 656152 503168 656180
rect 225012 656140 225018 656152
rect 503162 656140 503168 656152
rect 503220 656140 503226 656192
rect 504542 655732 504548 655784
rect 504600 655772 504606 655784
rect 580626 655772 580632 655784
rect 504600 655744 580632 655772
rect 504600 655732 504606 655744
rect 580626 655732 580632 655744
rect 580684 655732 580690 655784
rect 500402 655664 500408 655716
rect 500460 655704 500466 655716
rect 577498 655704 577504 655716
rect 500460 655676 577504 655704
rect 500460 655664 500466 655676
rect 577498 655664 577504 655676
rect 577556 655664 577562 655716
rect 489270 655596 489276 655648
rect 489328 655636 489334 655648
rect 499022 655636 499028 655648
rect 489328 655608 499028 655636
rect 489328 655596 489334 655608
rect 499022 655596 499028 655608
rect 499080 655596 499086 655648
rect 501782 655596 501788 655648
rect 501840 655636 501846 655648
rect 580350 655636 580356 655648
rect 501840 655608 580356 655636
rect 501840 655596 501846 655608
rect 580350 655596 580356 655608
rect 580408 655596 580414 655648
rect 237650 655528 237656 655580
rect 237708 655568 237714 655580
rect 528002 655568 528008 655580
rect 237708 655540 528008 655568
rect 237708 655528 237714 655540
rect 528002 655528 528008 655540
rect 528060 655528 528066 655580
rect 231578 654780 231584 654832
rect 231636 654820 231642 654832
rect 514754 654820 514760 654832
rect 231636 654792 514760 654820
rect 231636 654780 231642 654792
rect 514754 654780 514760 654792
rect 514812 654780 514818 654832
rect 274542 654508 274548 654560
rect 274600 654548 274606 654560
rect 536006 654548 536012 654560
rect 274600 654520 536012 654548
rect 274600 654508 274606 654520
rect 536006 654508 536012 654520
rect 536064 654508 536070 654560
rect 286962 654440 286968 654492
rect 287020 654480 287026 654492
rect 538766 654480 538772 654492
rect 287020 654452 538772 654480
rect 287020 654440 287026 654452
rect 538766 654440 538772 654452
rect 538824 654440 538830 654492
rect 243722 650632 243728 650684
rect 243780 650672 243786 650684
rect 490374 650672 490380 650684
rect 243780 650644 490380 650672
rect 243780 650632 243786 650644
rect 490374 650632 490380 650644
rect 490432 650632 490438 650684
rect 255958 647844 255964 647896
rect 256016 647884 256022 647896
rect 489178 647884 489184 647896
rect 256016 647856 489184 647884
rect 256016 647844 256022 647856
rect 489178 647844 489184 647856
rect 489236 647844 489242 647896
rect 577590 643084 577596 643136
rect 577648 643124 577654 643136
rect 580718 643124 580724 643136
rect 577648 643096 580724 643124
rect 577648 643084 577654 643096
rect 580718 643084 580724 643096
rect 580776 643084 580782 643136
rect 281442 642336 281448 642388
rect 281500 642376 281506 642388
rect 487890 642376 487896 642388
rect 281500 642348 487896 642376
rect 281500 642336 281506 642348
rect 487890 642336 487896 642348
rect 487948 642336 487954 642388
rect 86862 633360 86868 633412
rect 86920 633400 86926 633412
rect 486970 633400 486976 633412
rect 86920 633372 486976 633400
rect 86920 633360 86926 633372
rect 486970 633360 486976 633372
rect 487028 633360 487034 633412
rect 88242 632884 88248 632936
rect 88300 632924 88306 632936
rect 255958 632924 255964 632936
rect 88300 632896 255964 632924
rect 88300 632884 88306 632896
rect 255958 632884 255964 632896
rect 256016 632884 256022 632936
rect 97994 632816 98000 632868
rect 98052 632856 98058 632868
rect 486878 632856 486884 632868
rect 98052 632828 486884 632856
rect 98052 632816 98058 632828
rect 486878 632816 486884 632828
rect 486936 632816 486942 632868
rect 91094 632748 91100 632800
rect 91152 632788 91158 632800
rect 91922 632788 91928 632800
rect 91152 632760 91928 632788
rect 91152 632748 91158 632760
rect 91922 632748 91928 632760
rect 91980 632788 91986 632800
rect 488442 632788 488448 632800
rect 91980 632760 488448 632788
rect 91980 632748 91986 632760
rect 488442 632748 488448 632760
rect 488500 632748 488506 632800
rect 85850 632720 85856 632732
rect 84166 632692 85856 632720
rect 54294 632272 54300 632324
rect 54352 632312 54358 632324
rect 84166 632312 84194 632692
rect 85850 632680 85856 632692
rect 85908 632720 85914 632732
rect 487062 632720 487068 632732
rect 85908 632692 487068 632720
rect 85908 632680 85914 632692
rect 487062 632680 487068 632692
rect 487120 632680 487126 632732
rect 54352 632284 84194 632312
rect 54352 632272 54358 632284
rect 286226 632272 286232 632324
rect 286284 632312 286290 632324
rect 286962 632312 286968 632324
rect 286284 632284 286968 632312
rect 286284 632272 286290 632284
rect 286962 632272 286968 632284
rect 287020 632312 287026 632324
rect 294138 632312 294144 632324
rect 287020 632284 294144 632312
rect 287020 632272 287026 632284
rect 294138 632272 294144 632284
rect 294196 632272 294202 632324
rect 486878 632272 486884 632324
rect 486936 632312 486942 632324
rect 488074 632312 488080 632324
rect 486936 632284 488080 632312
rect 486936 632272 486942 632284
rect 488074 632272 488080 632284
rect 488132 632272 488138 632324
rect 55950 632204 55956 632256
rect 56008 632244 56014 632256
rect 91094 632244 91100 632256
rect 56008 632216 91100 632244
rect 56008 632204 56014 632216
rect 91094 632204 91100 632216
rect 91152 632204 91158 632256
rect 280154 632204 280160 632256
rect 280212 632244 280218 632256
rect 281442 632244 281448 632256
rect 280212 632216 281448 632244
rect 280212 632204 280218 632216
rect 281442 632204 281448 632216
rect 281500 632244 281506 632256
rect 293034 632244 293040 632256
rect 281500 632216 293040 632244
rect 281500 632204 281506 632216
rect 293034 632204 293040 632216
rect 293092 632204 293098 632256
rect 487062 632204 487068 632256
rect 487120 632244 487126 632256
rect 487982 632244 487988 632256
rect 487120 632216 487988 632244
rect 487120 632204 487126 632216
rect 487982 632204 487988 632216
rect 488040 632204 488046 632256
rect 57606 632136 57612 632188
rect 57664 632176 57670 632188
rect 97994 632176 98000 632188
rect 57664 632148 98000 632176
rect 57664 632136 57670 632148
rect 97994 632136 98000 632148
rect 98052 632136 98058 632188
rect 274542 632136 274548 632188
rect 274600 632176 274606 632188
rect 294322 632176 294328 632188
rect 274600 632148 294328 632176
rect 274600 632136 274606 632148
rect 294322 632136 294328 632148
rect 294380 632136 294386 632188
rect 486970 632136 486976 632188
rect 487028 632176 487034 632188
rect 487890 632176 487896 632188
rect 487028 632148 487896 632176
rect 487028 632136 487034 632148
rect 487890 632136 487896 632148
rect 487948 632136 487954 632188
rect 488442 632136 488448 632188
rect 488500 632176 488506 632188
rect 489178 632176 489184 632188
rect 488500 632148 489184 632176
rect 488500 632136 488506 632148
rect 489178 632136 489184 632148
rect 489236 632136 489242 632188
rect 50982 632068 50988 632120
rect 51040 632108 51046 632120
rect 73706 632108 73712 632120
rect 51040 632080 73712 632108
rect 51040 632068 51046 632080
rect 73706 632068 73712 632080
rect 73764 632108 73770 632120
rect 490558 632108 490564 632120
rect 73764 632080 490564 632108
rect 73764 632068 73770 632080
rect 490558 632068 490564 632080
rect 490616 632068 490622 632120
rect 65886 630640 65892 630692
rect 65944 630680 65950 630692
rect 128814 630680 128820 630692
rect 65944 630652 128820 630680
rect 65944 630640 65950 630652
rect 128814 630640 128820 630652
rect 128872 630640 128878 630692
rect 62758 629620 62764 629672
rect 62816 629660 62822 629672
rect 115934 629660 115940 629672
rect 62816 629632 115940 629660
rect 62816 629620 62822 629632
rect 115934 629620 115940 629632
rect 115992 629620 115998 629672
rect 64414 629552 64420 629604
rect 64472 629592 64478 629604
rect 122006 629592 122012 629604
rect 64472 629564 122012 629592
rect 64472 629552 64478 629564
rect 122006 629552 122012 629564
rect 122064 629552 122070 629604
rect 68922 629484 68928 629536
rect 68980 629524 68986 629536
rect 231302 629524 231308 629536
rect 68980 629496 231308 629524
rect 68980 629484 68986 629496
rect 231302 629484 231308 629496
rect 231360 629484 231366 629536
rect 67450 629416 67456 629468
rect 67508 629456 67514 629468
rect 237374 629456 237380 629468
rect 67508 629428 237380 629456
rect 67508 629416 67514 629428
rect 237374 629416 237380 629428
rect 237432 629416 237438 629468
rect 67542 629348 67548 629400
rect 67600 629388 67606 629400
rect 243446 629388 243452 629400
rect 67600 629360 243452 629388
rect 67600 629348 67606 629360
rect 243446 629348 243452 629360
rect 243504 629348 243510 629400
rect 67450 629280 67456 629332
rect 67508 629320 67514 629332
rect 134150 629320 134156 629332
rect 67508 629292 134156 629320
rect 67508 629280 67514 629292
rect 134150 629280 134156 629292
rect 134208 629280 134214 629332
rect 490558 594056 490564 594108
rect 490616 594096 490622 594108
rect 511258 594096 511264 594108
rect 490616 594068 511264 594096
rect 490616 594056 490622 594068
rect 511258 594056 511264 594068
rect 511316 594056 511322 594108
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 60734 527184 60740 527196
rect 3476 527156 60740 527184
rect 3476 527144 3482 527156
rect 60734 527144 60740 527156
rect 60792 527144 60798 527196
rect 227714 478796 227720 478848
rect 227772 478836 227778 478848
rect 544102 478836 544108 478848
rect 227772 478808 544108 478836
rect 227772 478796 227778 478808
rect 544102 478796 544108 478808
rect 544160 478796 544166 478848
rect 231762 478728 231768 478780
rect 231820 478768 231826 478780
rect 294138 478768 294144 478780
rect 231820 478740 294144 478768
rect 231820 478728 231826 478740
rect 294138 478728 294144 478740
rect 294196 478728 294202 478780
rect 233142 478660 233148 478712
rect 233200 478700 233206 478712
rect 293034 478700 293040 478712
rect 233200 478672 293040 478700
rect 233200 478660 233206 478672
rect 293034 478660 293040 478672
rect 293092 478660 293098 478712
rect 241422 478592 241428 478644
rect 241480 478632 241486 478644
rect 294322 478632 294328 478644
rect 241480 478604 294328 478632
rect 241480 478592 241486 478604
rect 294322 478592 294328 478604
rect 294380 478592 294386 478644
rect 231486 478320 231492 478372
rect 231544 478360 231550 478372
rect 540146 478360 540152 478372
rect 231544 478332 540152 478360
rect 231544 478320 231550 478332
rect 540146 478320 540152 478332
rect 540204 478320 540210 478372
rect 234338 478252 234344 478304
rect 234396 478292 234402 478304
rect 542998 478292 543004 478304
rect 234396 478264 543004 478292
rect 234396 478252 234402 478264
rect 542998 478252 543004 478264
rect 543056 478252 543062 478304
rect 231670 478184 231676 478236
rect 231728 478224 231734 478236
rect 580534 478224 580540 478236
rect 231728 478196 580540 478224
rect 231728 478184 231734 478196
rect 580534 478184 580540 478196
rect 580592 478184 580598 478236
rect 230106 478116 230112 478168
rect 230164 478156 230170 478168
rect 580626 478156 580632 478168
rect 230164 478128 580632 478156
rect 230164 478116 230170 478128
rect 580626 478116 580632 478128
rect 580684 478116 580690 478168
rect 68462 477640 68468 477692
rect 68520 477680 68526 477692
rect 126238 477680 126244 477692
rect 68520 477652 126244 477680
rect 68520 477640 68526 477652
rect 126238 477640 126244 477652
rect 126296 477640 126302 477692
rect 68094 477572 68100 477624
rect 68152 477612 68158 477624
rect 138658 477612 138664 477624
rect 68152 477584 138664 477612
rect 68152 477572 68158 477584
rect 138658 477572 138664 477584
rect 138716 477572 138722 477624
rect 68186 477504 68192 477556
rect 68244 477544 68250 477556
rect 142890 477544 142896 477556
rect 68244 477516 142896 477544
rect 68244 477504 68250 477516
rect 142890 477504 142896 477516
rect 142948 477504 142954 477556
rect 3418 476008 3424 476060
rect 3476 476048 3482 476060
rect 62114 476048 62120 476060
rect 3476 476020 62120 476048
rect 3476 476008 3482 476020
rect 62114 476008 62120 476020
rect 62172 476008 62178 476060
rect 243538 476008 243544 476060
rect 243596 476048 243602 476060
rect 542722 476048 542728 476060
rect 243596 476020 542728 476048
rect 243596 476008 243602 476020
rect 542722 476008 542728 476020
rect 542780 476008 542786 476060
rect 251082 475940 251088 475992
rect 251140 475980 251146 475992
rect 508682 475980 508688 475992
rect 251140 475952 508688 475980
rect 251140 475940 251146 475952
rect 508682 475940 508688 475952
rect 508740 475940 508746 475992
rect 231854 475872 231860 475924
rect 231912 475912 231918 475924
rect 485038 475912 485044 475924
rect 231912 475884 485044 475912
rect 231912 475872 231918 475884
rect 485038 475872 485044 475884
rect 485096 475872 485102 475924
rect 262858 475804 262864 475856
rect 262916 475844 262922 475856
rect 507302 475844 507308 475856
rect 262916 475816 507308 475844
rect 262916 475804 262922 475816
rect 507302 475804 507308 475816
rect 507360 475804 507366 475856
rect 271782 475736 271788 475788
rect 271840 475776 271846 475788
rect 505922 475776 505928 475788
rect 271840 475748 505928 475776
rect 271840 475736 271846 475748
rect 505922 475736 505928 475748
rect 505980 475736 505986 475788
rect 233878 475668 233884 475720
rect 233936 475708 233942 475720
rect 462314 475708 462320 475720
rect 233936 475680 462320 475708
rect 233936 475668 233942 475680
rect 462314 475668 462320 475680
rect 462372 475668 462378 475720
rect 235626 475396 235632 475448
rect 235684 475436 235690 475448
rect 542630 475436 542636 475448
rect 235684 475408 542636 475436
rect 235684 475396 235690 475408
rect 542630 475396 542636 475408
rect 542688 475396 542694 475448
rect 62114 475328 62120 475380
rect 62172 475368 62178 475380
rect 63218 475368 63224 475380
rect 62172 475340 63224 475368
rect 62172 475328 62178 475340
rect 63218 475328 63224 475340
rect 63276 475368 63282 475380
rect 94038 475368 94044 475380
rect 63276 475340 94044 475368
rect 63276 475328 63282 475340
rect 94038 475328 94044 475340
rect 94096 475328 94102 475380
rect 233050 475328 233056 475380
rect 233108 475368 233114 475380
rect 577590 475368 577596 475380
rect 233108 475340 577596 475368
rect 233108 475328 233114 475340
rect 577590 475328 577596 475340
rect 577648 475328 577654 475380
rect 231394 474308 231400 474360
rect 231452 474348 231458 474360
rect 231670 474348 231676 474360
rect 231452 474320 231676 474348
rect 231452 474308 231458 474320
rect 231670 474308 231676 474320
rect 231728 474308 231734 474360
rect 230290 473288 230296 473340
rect 230348 473328 230354 473340
rect 544194 473328 544200 473340
rect 230348 473300 544200 473328
rect 230348 473288 230354 473300
rect 544194 473288 544200 473300
rect 544252 473288 544258 473340
rect 230382 473220 230388 473272
rect 230440 473260 230446 473272
rect 544010 473260 544016 473272
rect 230440 473232 544016 473260
rect 230440 473220 230446 473232
rect 544010 473220 544016 473232
rect 544068 473220 544074 473272
rect 238478 473152 238484 473204
rect 238536 473192 238542 473204
rect 541158 473192 541164 473204
rect 238536 473164 541164 473192
rect 238536 473152 238542 473164
rect 541158 473152 541164 473164
rect 541216 473152 541222 473204
rect 247034 473084 247040 473136
rect 247092 473124 247098 473136
rect 526622 473124 526628 473136
rect 247092 473096 526628 473124
rect 247092 473084 247098 473096
rect 526622 473084 526628 473096
rect 526680 473084 526686 473136
rect 255314 473016 255320 473068
rect 255372 473056 255378 473068
rect 525242 473056 525248 473068
rect 255372 473028 525248 473056
rect 255372 473016 255378 473028
rect 525242 473016 525248 473028
rect 525300 473016 525306 473068
rect 232774 472608 232780 472660
rect 232832 472648 232838 472660
rect 539042 472648 539048 472660
rect 232832 472620 539048 472648
rect 232832 472608 232838 472620
rect 539042 472608 539048 472620
rect 539100 472608 539106 472660
rect 230014 471860 230020 471912
rect 230072 471900 230078 471912
rect 230290 471900 230296 471912
rect 230072 471872 230296 471900
rect 230072 471860 230078 471872
rect 230290 471860 230296 471872
rect 230348 471860 230354 471912
rect 240042 443028 240048 443080
rect 240100 443068 240106 443080
rect 288710 443068 288716 443080
rect 240100 443040 288716 443068
rect 240100 443028 240106 443040
rect 288710 443028 288716 443040
rect 288768 443028 288774 443080
rect 237374 442960 237380 443012
rect 237432 443000 237438 443012
rect 288618 443000 288624 443012
rect 237432 442972 288624 443000
rect 237432 442960 237438 442972
rect 288618 442960 288624 442972
rect 288676 442960 288682 443012
rect 69658 442892 69664 442944
rect 69716 442932 69722 442944
rect 70210 442932 70216 442944
rect 69716 442904 70216 442932
rect 69716 442892 69722 442904
rect 70210 442892 70216 442904
rect 70268 442892 70274 442944
rect 233970 442892 233976 442944
rect 234028 442932 234034 442944
rect 488166 442932 488172 442944
rect 234028 442904 488172 442932
rect 234028 442892 234034 442904
rect 488166 442892 488172 442904
rect 488224 442892 488230 442944
rect 277210 442348 277216 442400
rect 277268 442388 277274 442400
rect 289446 442388 289452 442400
rect 277268 442360 289452 442388
rect 277268 442348 277274 442360
rect 289446 442348 289452 442360
rect 289504 442348 289510 442400
rect 238478 442280 238484 442332
rect 238536 442320 238542 442332
rect 541066 442320 541072 442332
rect 238536 442292 541072 442320
rect 238536 442280 238542 442292
rect 541066 442280 541072 442292
rect 541124 442280 541130 442332
rect 69658 442212 69664 442264
rect 69716 442252 69722 442264
rect 489270 442252 489276 442264
rect 69716 442224 489276 442252
rect 69716 442212 69722 442224
rect 489270 442212 489276 442224
rect 489328 442212 489334 442264
rect 229002 442144 229008 442196
rect 229060 442184 229066 442196
rect 288802 442184 288808 442196
rect 229060 442156 288808 442184
rect 229060 442144 229066 442156
rect 288802 442144 288808 442156
rect 288860 442144 288866 442196
rect 223482 442076 223488 442128
rect 223540 442116 223546 442128
rect 267734 442116 267740 442128
rect 223540 442088 267740 442116
rect 223540 442076 223546 442088
rect 267734 442076 267740 442088
rect 267792 442076 267798 442128
rect 270402 442076 270408 442128
rect 270460 442116 270466 442128
rect 284478 442116 284484 442128
rect 270460 442088 284484 442116
rect 270460 442076 270466 442088
rect 284478 442076 284484 442088
rect 284536 442076 284542 442128
rect 240042 442008 240048 442060
rect 240100 442048 240106 442060
rect 242802 442048 242808 442060
rect 240100 442020 242808 442048
rect 240100 442008 240106 442020
rect 242802 442008 242808 442020
rect 242860 442008 242866 442060
rect 254026 442008 254032 442060
rect 254084 442048 254090 442060
rect 280430 442048 280436 442060
rect 254084 442020 280436 442048
rect 254084 442008 254090 442020
rect 280430 442008 280436 442020
rect 280488 442008 280494 442060
rect 253934 441940 253940 441992
rect 253992 441980 253998 441992
rect 280706 441980 280712 441992
rect 253992 441952 280712 441980
rect 253992 441940 253998 441952
rect 280706 441940 280712 441952
rect 280764 441940 280770 441992
rect 251082 441872 251088 441924
rect 251140 441912 251146 441924
rect 282914 441912 282920 441924
rect 251140 441884 282920 441912
rect 251140 441872 251146 441884
rect 282914 441872 282920 441884
rect 282972 441872 282978 441924
rect 264974 441804 264980 441856
rect 265032 441844 265038 441856
rect 281074 441844 281080 441856
rect 265032 441816 281080 441844
rect 265032 441804 265038 441816
rect 281074 441804 281080 441816
rect 281132 441804 281138 441856
rect 239858 441736 239864 441788
rect 239916 441776 239922 441788
rect 289722 441776 289728 441788
rect 239916 441748 289728 441776
rect 239916 441736 239922 441748
rect 289722 441736 289728 441748
rect 289780 441736 289786 441788
rect 239214 441668 239220 441720
rect 239272 441708 239278 441720
rect 289630 441708 289636 441720
rect 239272 441680 289636 441708
rect 239272 441668 239278 441680
rect 289630 441668 289636 441680
rect 289688 441668 289694 441720
rect 273254 441600 273260 441652
rect 273312 441640 273318 441652
rect 284386 441640 284392 441652
rect 273312 441612 284392 441640
rect 273312 441600 273318 441612
rect 284386 441600 284392 441612
rect 284444 441600 284450 441652
rect 267734 441532 267740 441584
rect 267792 441572 267798 441584
rect 474734 441572 474740 441584
rect 267792 441544 474740 441572
rect 267792 441532 267798 441544
rect 474734 441532 474740 441544
rect 474792 441532 474798 441584
rect 238386 440988 238392 441040
rect 238444 441028 238450 441040
rect 539870 441028 539876 441040
rect 238444 441000 539876 441028
rect 238444 440988 238450 441000
rect 539870 440988 539876 441000
rect 539928 440988 539934 441040
rect 238202 440920 238208 440972
rect 238260 440960 238266 440972
rect 539686 440960 539692 440972
rect 238260 440932 539692 440960
rect 238260 440920 238266 440932
rect 539686 440920 539692 440932
rect 539744 440920 539750 440972
rect 238110 440852 238116 440904
rect 238168 440892 238174 440904
rect 540974 440892 540980 440904
rect 238168 440864 540980 440892
rect 238168 440852 238174 440864
rect 540974 440852 540980 440864
rect 541032 440852 541038 440904
rect 240778 440716 240784 440768
rect 240836 440756 240842 440768
rect 287698 440756 287704 440768
rect 240836 440728 287704 440756
rect 240836 440716 240842 440728
rect 287698 440716 287704 440728
rect 287756 440716 287762 440768
rect 232682 440648 232688 440700
rect 232740 440688 232746 440700
rect 282086 440688 282092 440700
rect 232740 440660 282092 440688
rect 232740 440648 232746 440660
rect 282086 440648 282092 440660
rect 282144 440648 282150 440700
rect 230474 440580 230480 440632
rect 230532 440620 230538 440632
rect 281074 440620 281080 440632
rect 230532 440592 281080 440620
rect 230532 440580 230538 440592
rect 281074 440580 281080 440592
rect 281132 440580 281138 440632
rect 231394 440512 231400 440564
rect 231452 440552 231458 440564
rect 281994 440552 282000 440564
rect 231452 440524 282000 440552
rect 231452 440512 231458 440524
rect 281994 440512 282000 440524
rect 282052 440512 282058 440564
rect 229646 440444 229652 440496
rect 229704 440484 229710 440496
rect 280982 440484 280988 440496
rect 229704 440456 280988 440484
rect 229704 440444 229710 440456
rect 280982 440444 280988 440456
rect 281040 440444 281046 440496
rect 228910 440376 228916 440428
rect 228968 440416 228974 440428
rect 280246 440416 280252 440428
rect 228968 440388 280252 440416
rect 228968 440376 228974 440388
rect 280246 440376 280252 440388
rect 280304 440376 280310 440428
rect 229002 440308 229008 440360
rect 229060 440348 229066 440360
rect 280522 440348 280528 440360
rect 229060 440320 280528 440348
rect 229060 440308 229066 440320
rect 280522 440308 280528 440320
rect 280580 440308 280586 440360
rect 221458 440240 221464 440292
rect 221516 440280 221522 440292
rect 223482 440280 223488 440292
rect 221516 440252 223488 440280
rect 221516 440240 221522 440252
rect 223482 440240 223488 440252
rect 223540 440240 223546 440292
rect 227162 440240 227168 440292
rect 227220 440280 227226 440292
rect 284294 440280 284300 440292
rect 227220 440252 284300 440280
rect 227220 440240 227226 440252
rect 284294 440240 284300 440252
rect 284352 440240 284358 440292
rect 474734 440240 474740 440292
rect 474792 440280 474798 440292
rect 475378 440280 475384 440292
rect 474792 440252 475384 440280
rect 474792 440240 474798 440252
rect 475378 440240 475384 440252
rect 475436 440240 475442 440292
rect 229370 439832 229376 439884
rect 229428 439872 229434 439884
rect 230014 439872 230020 439884
rect 229428 439844 230020 439872
rect 229428 439832 229434 439844
rect 230014 439832 230020 439844
rect 230072 439832 230078 439884
rect 239766 439696 239772 439748
rect 239824 439736 239830 439748
rect 580258 439736 580264 439748
rect 239824 439708 580264 439736
rect 239824 439696 239830 439708
rect 580258 439696 580264 439708
rect 580316 439696 580322 439748
rect 228726 439628 228732 439680
rect 228784 439668 228790 439680
rect 280154 439668 280160 439680
rect 228784 439640 280160 439668
rect 228784 439628 228790 439640
rect 280154 439628 280160 439640
rect 280212 439628 280218 439680
rect 229002 439560 229008 439612
rect 229060 439600 229066 439612
rect 280614 439600 280620 439612
rect 229060 439572 280620 439600
rect 229060 439560 229066 439572
rect 280614 439560 280620 439572
rect 280672 439560 280678 439612
rect 231394 439492 231400 439544
rect 231452 439532 231458 439544
rect 280062 439532 280068 439544
rect 231452 439504 280068 439532
rect 231452 439492 231458 439504
rect 280062 439492 280068 439504
rect 280120 439492 280126 439544
rect 229646 439424 229652 439476
rect 229704 439464 229710 439476
rect 280890 439464 280896 439476
rect 229704 439436 280896 439464
rect 229704 439424 229710 439436
rect 280890 439424 280896 439436
rect 280948 439424 280954 439476
rect 231026 439356 231032 439408
rect 231084 439396 231090 439408
rect 281810 439396 281816 439408
rect 231084 439368 281816 439396
rect 231084 439356 231090 439368
rect 281810 439356 281816 439368
rect 281868 439356 281874 439408
rect 228266 439084 228272 439136
rect 228324 439124 228330 439136
rect 228726 439124 228732 439136
rect 228324 439096 228732 439124
rect 228324 439084 228330 439096
rect 228726 439084 228732 439096
rect 228784 439084 228790 439136
rect 218054 438880 218060 438932
rect 218112 438920 218118 438932
rect 221458 438920 221464 438932
rect 218112 438892 221464 438920
rect 218112 438880 218118 438892
rect 221458 438880 221464 438892
rect 221516 438880 221522 438932
rect 239214 436772 239220 436824
rect 239272 436812 239278 436824
rect 239766 436812 239772 436824
rect 239272 436784 239772 436812
rect 239272 436772 239278 436784
rect 239766 436772 239772 436784
rect 239824 436772 239830 436824
rect 280890 436500 280896 436552
rect 280948 436540 280954 436552
rect 281074 436540 281080 436552
rect 280948 436512 281080 436540
rect 280948 436500 280954 436512
rect 281074 436500 281080 436512
rect 281132 436500 281138 436552
rect 281626 435548 281632 435600
rect 281684 435588 281690 435600
rect 282086 435588 282092 435600
rect 281684 435560 282092 435588
rect 281684 435548 281690 435560
rect 282086 435548 282092 435560
rect 282144 435548 282150 435600
rect 218054 434772 218060 434784
rect 213932 434744 218060 434772
rect 213546 434664 213552 434716
rect 213604 434704 213610 434716
rect 213932 434704 213960 434744
rect 218054 434732 218060 434744
rect 218112 434732 218118 434784
rect 213604 434676 213960 434704
rect 213604 434664 213610 434676
rect 281534 434188 281540 434240
rect 281592 434228 281598 434240
rect 281994 434228 282000 434240
rect 281592 434200 282000 434228
rect 281592 434188 281598 434200
rect 281994 434188 282000 434200
rect 282052 434188 282058 434240
rect 211614 430584 211620 430636
rect 211672 430624 211678 430636
rect 213546 430624 213552 430636
rect 211672 430596 213552 430624
rect 211672 430584 211678 430596
rect 213546 430584 213552 430596
rect 213604 430584 213610 430636
rect 3418 423580 3424 423632
rect 3476 423620 3482 423632
rect 60734 423620 60740 423632
rect 3476 423592 60740 423620
rect 3476 423580 3482 423592
rect 60734 423580 60740 423592
rect 60792 423580 60798 423632
rect 60734 422900 60740 422952
rect 60792 422940 60798 422952
rect 61838 422940 61844 422952
rect 60792 422912 61844 422940
rect 60792 422900 60798 422912
rect 61838 422900 61844 422912
rect 61896 422940 61902 422952
rect 95694 422940 95700 422952
rect 61896 422912 95700 422940
rect 61896 422900 61902 422912
rect 95694 422900 95700 422912
rect 95752 422900 95758 422952
rect 207014 422288 207020 422340
rect 207072 422328 207078 422340
rect 211614 422328 211620 422340
rect 207072 422300 211620 422328
rect 207072 422288 207078 422300
rect 211614 422288 211620 422300
rect 211672 422288 211678 422340
rect 207014 418180 207020 418192
rect 205652 418152 207020 418180
rect 202874 418072 202880 418124
rect 202932 418112 202938 418124
rect 205652 418112 205680 418152
rect 207014 418140 207020 418152
rect 207072 418140 207078 418192
rect 202932 418084 205680 418112
rect 202932 418072 202938 418084
rect 198826 412632 198832 412684
rect 198884 412672 198890 412684
rect 202782 412672 202788 412684
rect 198884 412644 202788 412672
rect 198884 412632 198890 412644
rect 202782 412632 202788 412644
rect 202840 412632 202846 412684
rect 281902 409776 281908 409828
rect 281960 409816 281966 409828
rect 284478 409816 284484 409828
rect 281960 409788 284484 409816
rect 281960 409776 281966 409788
rect 284478 409776 284484 409788
rect 284536 409776 284542 409828
rect 197998 408484 198004 408536
rect 198056 408524 198062 408536
rect 198826 408524 198832 408536
rect 198056 408496 198832 408524
rect 198056 408484 198062 408496
rect 198826 408484 198832 408496
rect 198884 408484 198890 408536
rect 281902 408416 281908 408468
rect 281960 408456 281966 408468
rect 284386 408456 284392 408468
rect 281960 408428 284392 408456
rect 281960 408416 281966 408428
rect 284386 408416 284392 408428
rect 284444 408416 284450 408468
rect 577498 405628 577504 405680
rect 577556 405668 577562 405680
rect 579706 405668 579712 405680
rect 577556 405640 579712 405668
rect 577556 405628 577562 405640
rect 579706 405628 579712 405640
rect 579764 405628 579770 405680
rect 197998 400228 198004 400240
rect 195992 400200 198004 400228
rect 193858 400120 193864 400172
rect 193916 400160 193922 400172
rect 195992 400160 196020 400200
rect 197998 400188 198004 400200
rect 198056 400188 198062 400240
rect 193916 400132 196020 400160
rect 193916 400120 193922 400132
rect 281810 394612 281816 394664
rect 281868 394652 281874 394664
rect 284294 394652 284300 394664
rect 281868 394624 284300 394652
rect 281868 394612 281874 394624
rect 284294 394612 284300 394624
rect 284352 394612 284358 394664
rect 191834 386316 191840 386368
rect 191892 386356 191898 386368
rect 193858 386356 193864 386368
rect 191892 386328 193864 386356
rect 191892 386316 191898 386328
rect 193858 386316 193864 386328
rect 193916 386316 193922 386368
rect 192478 383664 192484 383716
rect 192536 383704 192542 383716
rect 237374 383704 237380 383716
rect 192536 383676 237380 383704
rect 192536 383664 192542 383676
rect 237374 383664 237380 383676
rect 237432 383664 237438 383716
rect 237374 382548 237380 382560
rect 219406 382520 237380 382548
rect 216030 382372 216036 382424
rect 216088 382412 216094 382424
rect 219406 382412 219434 382520
rect 237374 382508 237380 382520
rect 237432 382508 237438 382560
rect 216088 382384 219434 382412
rect 216088 382372 216094 382384
rect 112530 382304 112536 382356
rect 112588 382344 112594 382356
rect 237374 382344 237380 382356
rect 112588 382316 237380 382344
rect 112588 382304 112594 382316
rect 237374 382304 237380 382316
rect 237432 382304 237438 382356
rect 112438 382236 112444 382288
rect 112496 382276 112502 382288
rect 237466 382276 237472 382288
rect 112496 382248 237472 382276
rect 112496 382236 112502 382248
rect 237466 382236 237472 382248
rect 237524 382236 237530 382288
rect 112714 380944 112720 380996
rect 112772 380984 112778 380996
rect 237558 380984 237564 380996
rect 112772 380956 237564 380984
rect 112772 380944 112778 380956
rect 237558 380944 237564 380956
rect 237616 380944 237622 380996
rect 111150 380876 111156 380928
rect 111208 380916 111214 380928
rect 237374 380916 237380 380928
rect 111208 380888 237380 380916
rect 111208 380876 111214 380888
rect 237374 380876 237380 380888
rect 237432 380876 237438 380928
rect 110046 379516 110052 379568
rect 110104 379556 110110 379568
rect 237374 379556 237380 379568
rect 110104 379528 237380 379556
rect 110104 379516 110110 379528
rect 237374 379516 237380 379528
rect 237432 379516 237438 379568
rect 186958 379448 186964 379500
rect 187016 379488 187022 379500
rect 191742 379488 191748 379500
rect 187016 379460 191748 379488
rect 187016 379448 187022 379460
rect 191742 379448 191748 379460
rect 191800 379448 191806 379500
rect 127618 376864 127624 376916
rect 127676 376904 127682 376916
rect 237374 376904 237380 376916
rect 127676 376876 237380 376904
rect 127676 376864 127682 376876
rect 237374 376864 237380 376876
rect 237432 376864 237438 376916
rect 123570 376796 123576 376848
rect 123628 376836 123634 376848
rect 237558 376836 237564 376848
rect 123628 376808 237564 376836
rect 123628 376796 123634 376808
rect 237558 376796 237564 376808
rect 237616 376796 237622 376848
rect 111518 376728 111524 376780
rect 111576 376768 111582 376780
rect 237742 376768 237748 376780
rect 111576 376740 237748 376768
rect 111576 376728 111582 376740
rect 237742 376728 237748 376740
rect 237800 376728 237806 376780
rect 126422 375436 126428 375488
rect 126480 375476 126486 375488
rect 237374 375476 237380 375488
rect 126480 375448 237380 375476
rect 126480 375436 126486 375448
rect 237374 375436 237380 375448
rect 237432 375436 237438 375488
rect 111610 375368 111616 375420
rect 111668 375408 111674 375420
rect 237558 375408 237564 375420
rect 111668 375380 237564 375408
rect 111668 375368 111674 375380
rect 237558 375368 237564 375380
rect 237616 375368 237622 375420
rect 237374 374320 237380 374332
rect 219406 374292 237380 374320
rect 122190 374076 122196 374128
rect 122248 374116 122254 374128
rect 219406 374116 219434 374292
rect 237374 374280 237380 374292
rect 237432 374280 237438 374332
rect 122248 374088 219434 374116
rect 122248 374076 122254 374088
rect 115290 374008 115296 374060
rect 115348 374048 115354 374060
rect 237374 374048 237380 374060
rect 115348 374020 237380 374048
rect 115348 374008 115354 374020
rect 237374 374008 237380 374020
rect 237432 374008 237438 374060
rect 3418 372512 3424 372564
rect 3476 372552 3482 372564
rect 63494 372552 63500 372564
rect 3476 372524 63500 372552
rect 3476 372512 3482 372524
rect 63494 372512 63500 372524
rect 63552 372512 63558 372564
rect 63494 371832 63500 371884
rect 63552 371872 63558 371884
rect 64598 371872 64604 371884
rect 63552 371844 64604 371872
rect 63552 371832 63558 371844
rect 64598 371832 64604 371844
rect 64656 371872 64662 371884
rect 97350 371872 97356 371884
rect 64656 371844 97356 371872
rect 64656 371832 64662 371844
rect 97350 371832 97356 371844
rect 97408 371832 97414 371884
rect 137278 371220 137284 371272
rect 137336 371260 137342 371272
rect 237374 371260 237380 371272
rect 137336 371232 237380 371260
rect 137336 371220 137342 371232
rect 237374 371220 237380 371232
rect 237432 371220 237438 371272
rect 115382 369860 115388 369912
rect 115440 369900 115446 369912
rect 237374 369900 237380 369912
rect 115440 369872 237380 369900
rect 115440 369860 115446 369872
rect 237374 369860 237380 369872
rect 237432 369860 237438 369912
rect 282822 368500 282828 368552
rect 282880 368540 282886 368552
rect 287146 368540 287152 368552
rect 282880 368512 287152 368540
rect 282880 368500 282886 368512
rect 287146 368500 287152 368512
rect 287204 368500 287210 368552
rect 489270 366324 489276 366376
rect 489328 366364 489334 366376
rect 498838 366364 498844 366376
rect 489328 366336 498844 366364
rect 489328 366324 489334 366336
rect 498838 366324 498844 366336
rect 498896 366324 498902 366376
rect 282822 358776 282828 358828
rect 282880 358816 282886 358828
rect 288986 358816 288992 358828
rect 282880 358788 288992 358816
rect 282880 358776 282886 358788
rect 288986 358776 288992 358788
rect 289044 358776 289050 358828
rect 185578 358708 185584 358760
rect 185636 358748 185642 358760
rect 186958 358748 186964 358760
rect 185636 358720 186964 358748
rect 185636 358708 185642 358720
rect 186958 358708 186964 358720
rect 187016 358708 187022 358760
rect 282822 356056 282828 356108
rect 282880 356096 282886 356108
rect 287238 356096 287244 356108
rect 282880 356068 287244 356096
rect 282880 356056 282886 356068
rect 287238 356056 287244 356068
rect 287296 356056 287302 356108
rect 282822 353268 282828 353320
rect 282880 353308 282886 353320
rect 289078 353308 289084 353320
rect 282880 353280 289084 353308
rect 282880 353268 282886 353280
rect 289078 353268 289084 353280
rect 289136 353268 289142 353320
rect 498838 353200 498844 353252
rect 498896 353240 498902 353252
rect 580166 353240 580172 353252
rect 498896 353212 580172 353240
rect 498896 353200 498902 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 60918 352520 60924 352572
rect 60976 352560 60982 352572
rect 69658 352560 69664 352572
rect 60976 352532 69664 352560
rect 60976 352520 60982 352532
rect 69658 352520 69664 352532
rect 69716 352520 69722 352572
rect 282822 347760 282828 347812
rect 282880 347800 282886 347812
rect 291286 347800 291292 347812
rect 282880 347772 291292 347800
rect 282880 347760 282886 347772
rect 291286 347760 291292 347772
rect 291344 347760 291350 347812
rect 182174 347692 182180 347744
rect 182232 347732 182238 347744
rect 185578 347732 185584 347744
rect 182232 347704 185584 347732
rect 182232 347692 182238 347704
rect 185578 347692 185584 347704
rect 185636 347692 185642 347744
rect 59078 344292 59084 344344
rect 59136 344332 59142 344344
rect 182174 344332 182180 344344
rect 59136 344304 182180 344332
rect 59136 344292 59142 344304
rect 182174 344292 182180 344304
rect 182232 344292 182238 344344
rect 475378 344292 475384 344344
rect 475436 344332 475442 344344
rect 497458 344332 497464 344344
rect 475436 344304 497464 344332
rect 475436 344292 475442 344304
rect 497458 344292 497464 344304
rect 497516 344292 497522 344344
rect 216674 343612 216680 343664
rect 216732 343652 216738 343664
rect 235258 343652 235264 343664
rect 216732 343624 235264 343652
rect 216732 343612 216738 343624
rect 235258 343612 235264 343624
rect 235316 343612 235322 343664
rect 282822 343612 282828 343664
rect 282880 343652 282886 343664
rect 287330 343652 287336 343664
rect 282880 343624 287336 343652
rect 282880 343612 282886 343624
rect 287330 343612 287336 343624
rect 287388 343612 287394 343664
rect 63586 342524 63592 342576
rect 63644 342564 63650 342576
rect 86954 342564 86960 342576
rect 63644 342536 86960 342564
rect 63644 342524 63650 342536
rect 86954 342524 86960 342536
rect 87012 342524 87018 342576
rect 66162 342456 66168 342508
rect 66220 342496 66226 342508
rect 92014 342496 92020 342508
rect 66220 342468 92020 342496
rect 66220 342456 66226 342468
rect 92014 342456 92020 342468
rect 92072 342456 92078 342508
rect 43438 342388 43444 342440
rect 43496 342428 43502 342440
rect 105262 342428 105268 342440
rect 43496 342400 105268 342428
rect 43496 342388 43502 342400
rect 105262 342388 105268 342400
rect 105320 342388 105326 342440
rect 15838 342320 15844 342372
rect 15896 342360 15902 342372
rect 106918 342360 106924 342372
rect 15896 342332 106924 342360
rect 15896 342320 15902 342332
rect 106918 342320 106924 342332
rect 106976 342320 106982 342372
rect 11698 342252 11704 342304
rect 11756 342292 11762 342304
rect 108298 342292 108304 342304
rect 11756 342264 108304 342292
rect 11756 342252 11762 342264
rect 108298 342252 108304 342264
rect 108356 342252 108362 342304
rect 99374 341776 99380 341828
rect 99432 341816 99438 341828
rect 100294 341816 100300 341828
rect 99432 341788 100300 341816
rect 99432 341776 99438 341788
rect 100294 341776 100300 341788
rect 100352 341776 100358 341828
rect 65794 341300 65800 341352
rect 65852 341340 65858 341352
rect 228818 341340 228824 341352
rect 65852 341312 228824 341340
rect 65852 341300 65858 341312
rect 228818 341300 228824 341312
rect 228876 341300 228882 341352
rect 39298 341232 39304 341284
rect 39356 341272 39362 341284
rect 104158 341272 104164 341284
rect 39356 341244 104164 341272
rect 39356 341232 39362 341244
rect 104158 341232 104164 341244
rect 104216 341232 104222 341284
rect 215938 341232 215944 341284
rect 215996 341272 216002 341284
rect 237558 341272 237564 341284
rect 215996 341244 237564 341272
rect 215996 341232 216002 341244
rect 237558 341232 237564 341244
rect 237616 341232 237622 341284
rect 25498 341164 25504 341216
rect 25556 341204 25562 341216
rect 99374 341204 99380 341216
rect 25556 341176 99380 341204
rect 25556 341164 25562 341176
rect 99374 341164 99380 341176
rect 99432 341164 99438 341216
rect 213178 341164 213184 341216
rect 213236 341204 213242 341216
rect 237374 341204 237380 341216
rect 213236 341176 237380 341204
rect 213236 341164 213242 341176
rect 237374 341164 237380 341176
rect 237432 341164 237438 341216
rect 70210 341096 70216 341148
rect 70268 341136 70274 341148
rect 225874 341136 225880 341148
rect 70268 341108 225880 341136
rect 70268 341096 70274 341108
rect 225874 341096 225880 341108
rect 225932 341096 225938 341148
rect 70302 341028 70308 341080
rect 70360 341068 70366 341080
rect 228634 341068 228640 341080
rect 70360 341040 228640 341068
rect 70360 341028 70366 341040
rect 228634 341028 228640 341040
rect 228692 341028 228698 341080
rect 67450 340960 67456 341012
rect 67508 341000 67514 341012
rect 228542 341000 228548 341012
rect 67508 340972 228548 341000
rect 67508 340960 67514 340972
rect 228542 340960 228548 340972
rect 228600 340960 228606 341012
rect 228358 340892 228364 340944
rect 228416 340932 228422 340944
rect 237374 340932 237380 340944
rect 228416 340904 237380 340932
rect 228416 340892 228422 340904
rect 237374 340892 237380 340904
rect 237432 340892 237438 340944
rect 43530 339532 43536 339584
rect 43588 339572 43594 339584
rect 102134 339572 102140 339584
rect 43588 339544 102140 339572
rect 43588 339532 43594 339544
rect 102134 339532 102140 339544
rect 102192 339532 102198 339584
rect 29638 339464 29644 339516
rect 29696 339504 29702 339516
rect 98638 339504 98644 339516
rect 29696 339476 98644 339504
rect 29696 339464 29702 339476
rect 98638 339464 98644 339476
rect 98696 339464 98702 339516
rect 3418 320084 3424 320136
rect 3476 320124 3482 320136
rect 29638 320124 29644 320136
rect 3476 320096 29644 320124
rect 3476 320084 3482 320096
rect 29638 320084 29644 320096
rect 29696 320084 29702 320136
rect 235258 300772 235264 300824
rect 235316 300812 235322 300824
rect 237374 300812 237380 300824
rect 235316 300784 237380 300812
rect 235316 300772 235322 300784
rect 237374 300772 237380 300784
rect 237432 300772 237438 300824
rect 497458 299412 497464 299464
rect 497516 299452 497522 299464
rect 580166 299452 580172 299464
rect 497516 299424 580172 299452
rect 497516 299412 497522 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 282822 295332 282828 295384
rect 282880 295372 282886 295384
rect 288526 295372 288532 295384
rect 282880 295344 288532 295372
rect 282880 295332 282886 295344
rect 288526 295332 288532 295344
rect 288584 295332 288590 295384
rect 142890 288328 142896 288380
rect 142948 288368 142954 288380
rect 237374 288368 237380 288380
rect 142948 288340 237380 288368
rect 142948 288328 142954 288340
rect 237374 288328 237380 288340
rect 237432 288328 237438 288380
rect 126238 286968 126244 287020
rect 126296 287008 126302 287020
rect 237374 287008 237380 287020
rect 126296 286980 237380 287008
rect 126296 286968 126302 286980
rect 237374 286968 237380 286980
rect 237432 286968 237438 287020
rect 138658 285608 138664 285660
rect 138716 285648 138722 285660
rect 237374 285648 237380 285660
rect 138716 285620 237380 285648
rect 138716 285608 138722 285620
rect 237374 285608 237380 285620
rect 237432 285608 237438 285660
rect 225874 282820 225880 282872
rect 225932 282860 225938 282872
rect 237374 282860 237380 282872
rect 225932 282832 237380 282860
rect 225932 282820 225938 282832
rect 237374 282820 237380 282832
rect 237432 282820 237438 282872
rect 228818 281460 228824 281512
rect 228876 281500 228882 281512
rect 237558 281500 237564 281512
rect 228876 281472 237564 281500
rect 228876 281460 228882 281472
rect 237558 281460 237564 281472
rect 237616 281460 237622 281512
rect 282822 281460 282828 281512
rect 282880 281500 282886 281512
rect 288802 281500 288808 281512
rect 282880 281472 288808 281500
rect 282880 281460 282886 281472
rect 288802 281460 288808 281472
rect 288860 281460 288866 281512
rect 228634 281392 228640 281444
rect 228692 281432 228698 281444
rect 237374 281432 237380 281444
rect 228692 281404 237380 281432
rect 228692 281392 228698 281404
rect 237374 281392 237380 281404
rect 237432 281392 237438 281444
rect 78950 280100 78956 280152
rect 79008 280140 79014 280152
rect 126422 280140 126428 280152
rect 79008 280112 126428 280140
rect 79008 280100 79014 280112
rect 126422 280100 126428 280112
rect 126480 280100 126486 280152
rect 228542 280100 228548 280152
rect 228600 280140 228606 280152
rect 237374 280140 237380 280152
rect 228600 280112 237380 280140
rect 228600 280100 228606 280112
rect 237374 280100 237380 280112
rect 237432 280100 237438 280152
rect 80054 280032 80060 280084
rect 80112 280072 80118 280084
rect 127618 280072 127624 280084
rect 80112 280044 127624 280072
rect 80112 280032 80118 280044
rect 127618 280032 127624 280044
rect 127676 280032 127682 280084
rect 78582 279964 78588 280016
rect 78640 280004 78646 280016
rect 122190 280004 122196 280016
rect 78640 279976 122196 280004
rect 78640 279964 78646 279976
rect 122190 279964 122196 279976
rect 122248 279964 122254 280016
rect 81434 279896 81440 279948
rect 81492 279936 81498 279948
rect 111610 279936 111616 279948
rect 81492 279908 111616 279936
rect 81492 279896 81498 279908
rect 111610 279896 111616 279908
rect 111668 279896 111674 279948
rect 96522 279828 96528 279880
rect 96580 279868 96586 279880
rect 123570 279868 123576 279880
rect 96580 279840 123576 279868
rect 96580 279828 96586 279840
rect 123570 279828 123576 279840
rect 123628 279828 123634 279880
rect 99374 279760 99380 279812
rect 99432 279800 99438 279812
rect 111518 279800 111524 279812
rect 99432 279772 111524 279800
rect 99432 279760 99438 279772
rect 111518 279760 111524 279772
rect 111576 279760 111582 279812
rect 98638 278672 98644 278724
rect 98696 278712 98702 278724
rect 111150 278712 111156 278724
rect 98696 278684 111156 278712
rect 98696 278672 98702 278684
rect 111150 278672 111156 278684
rect 111208 278672 111214 278724
rect 97902 278604 97908 278656
rect 97960 278644 97966 278656
rect 110046 278644 110052 278656
rect 97960 278616 110052 278644
rect 97960 278604 97966 278616
rect 110046 278604 110052 278616
rect 110104 278604 110110 278656
rect 89714 278536 89720 278588
rect 89772 278576 89778 278588
rect 137278 278576 137284 278588
rect 89772 278548 137284 278576
rect 89772 278536 89778 278548
rect 137278 278536 137284 278548
rect 137336 278536 137342 278588
rect 91094 278468 91100 278520
rect 91152 278508 91158 278520
rect 115382 278508 115388 278520
rect 91152 278480 115388 278508
rect 91152 278468 91158 278480
rect 115382 278468 115388 278480
rect 115440 278468 115446 278520
rect 95142 278400 95148 278452
rect 95200 278440 95206 278452
rect 115290 278440 115296 278452
rect 95200 278412 115296 278440
rect 95200 278400 95206 278412
rect 115290 278400 115296 278412
rect 115348 278400 115354 278452
rect 102134 278332 102140 278384
rect 102192 278372 102198 278384
rect 102192 278344 103514 278372
rect 102192 278332 102198 278344
rect 103486 278304 103514 278344
rect 106182 278332 106188 278384
rect 106240 278372 106246 278384
rect 112438 278372 112444 278384
rect 106240 278344 112444 278372
rect 106240 278332 106246 278344
rect 112438 278332 112444 278344
rect 112496 278332 112502 278384
rect 112530 278332 112536 278384
rect 112588 278332 112594 278384
rect 112548 278304 112576 278332
rect 103486 278276 112576 278304
rect 104802 278196 104808 278248
rect 104860 278236 104866 278248
rect 112714 278236 112720 278248
rect 104860 278208 112720 278236
rect 104860 278196 104866 278208
rect 112714 278196 112720 278208
rect 112772 278196 112778 278248
rect 107378 278128 107384 278180
rect 107436 278168 107442 278180
rect 216030 278168 216036 278180
rect 107436 278140 216036 278168
rect 107436 278128 107442 278140
rect 216030 278128 216036 278140
rect 216088 278128 216094 278180
rect 108298 278060 108304 278112
rect 108356 278100 108362 278112
rect 192478 278100 192484 278112
rect 108356 278072 192484 278100
rect 108356 278060 108362 278072
rect 192478 278060 192484 278072
rect 192536 278060 192542 278112
rect 282822 274592 282828 274644
rect 282880 274632 282886 274644
rect 288710 274632 288716 274644
rect 282880 274604 288716 274632
rect 282880 274592 282886 274604
rect 288710 274592 288716 274604
rect 288768 274592 288774 274644
rect 282822 273164 282828 273216
rect 282880 273204 282886 273216
rect 288618 273204 288624 273216
rect 282880 273176 288624 273204
rect 282880 273164 282886 273176
rect 288618 273164 288624 273176
rect 288676 273164 288682 273216
rect 3418 267656 3424 267708
rect 3476 267696 3482 267708
rect 25498 267696 25504 267708
rect 3476 267668 25504 267696
rect 3476 267656 3482 267668
rect 25498 267656 25504 267668
rect 25556 267656 25562 267708
rect 488074 245556 488080 245608
rect 488132 245596 488138 245608
rect 580166 245596 580172 245608
rect 488132 245568 580172 245596
rect 488132 245556 488138 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 284846 243516 284852 243568
rect 284904 243556 284910 243568
rect 285122 243556 285128 243568
rect 284904 243528 285128 243556
rect 284904 243516 284910 243528
rect 285122 243516 285128 243528
rect 285180 243516 285186 243568
rect 284478 243380 284484 243432
rect 284536 243420 284542 243432
rect 284846 243420 284852 243432
rect 284536 243392 284852 243420
rect 284536 243380 284542 243392
rect 284846 243380 284852 243392
rect 284904 243380 284910 243432
rect 186314 240048 186320 240100
rect 186372 240088 186378 240100
rect 282362 240088 282368 240100
rect 186372 240060 282368 240088
rect 186372 240048 186378 240060
rect 282362 240048 282368 240060
rect 282420 240048 282426 240100
rect 212442 239980 212448 240032
rect 212500 240020 212506 240032
rect 287330 240020 287336 240032
rect 212500 239992 287336 240020
rect 212500 239980 212506 239992
rect 287330 239980 287336 239992
rect 287388 239980 287394 240032
rect 235994 239912 236000 239964
rect 236052 239952 236058 239964
rect 291286 239952 291292 239964
rect 236052 239924 291292 239952
rect 236052 239912 236058 239924
rect 291286 239912 291292 239924
rect 291344 239912 291350 239964
rect 237466 239844 237472 239896
rect 237524 239884 237530 239896
rect 289078 239884 289084 239896
rect 237524 239856 289084 239884
rect 237524 239844 237530 239856
rect 289078 239844 289084 239856
rect 289136 239844 289142 239896
rect 237558 239776 237564 239828
rect 237616 239816 237622 239828
rect 287238 239816 287244 239828
rect 237616 239788 287244 239816
rect 237616 239776 237622 239788
rect 287238 239776 287244 239788
rect 287296 239776 287302 239828
rect 237374 239708 237380 239760
rect 237432 239748 237438 239760
rect 280890 239748 280896 239760
rect 237432 239720 280896 239748
rect 237432 239708 237438 239720
rect 280890 239708 280896 239720
rect 280948 239708 280954 239760
rect 259270 239640 259276 239692
rect 259328 239680 259334 239692
rect 288986 239680 288992 239692
rect 259328 239652 288992 239680
rect 259328 239640 259334 239652
rect 288986 239640 288992 239652
rect 289044 239640 289050 239692
rect 264974 239572 264980 239624
rect 265032 239612 265038 239624
rect 287146 239612 287152 239624
rect 265032 239584 287152 239612
rect 265032 239572 265038 239584
rect 287146 239572 287152 239584
rect 287204 239572 287210 239624
rect 179414 239368 179420 239420
rect 179472 239408 179478 239420
rect 284478 239408 284484 239420
rect 179472 239380 284484 239408
rect 179472 239368 179478 239380
rect 284478 239368 284484 239380
rect 284536 239368 284542 239420
rect 44174 238688 44180 238740
rect 44232 238728 44238 238740
rect 243814 238728 243820 238740
rect 44232 238700 243820 238728
rect 44232 238688 44238 238700
rect 243814 238688 243820 238700
rect 243872 238688 243878 238740
rect 121454 238620 121460 238672
rect 121512 238660 121518 238672
rect 245010 238660 245016 238672
rect 121512 238632 245016 238660
rect 121512 238620 121518 238632
rect 245010 238620 245016 238632
rect 245068 238620 245074 238672
rect 3418 215228 3424 215280
rect 3476 215268 3482 215280
rect 43530 215268 43536 215280
rect 3476 215240 43536 215268
rect 3476 215228 3482 215240
rect 43530 215228 43536 215240
rect 43588 215228 43594 215280
rect 489178 206932 489184 206984
rect 489236 206972 489242 206984
rect 580166 206972 580172 206984
rect 489236 206944 580172 206972
rect 489236 206932 489242 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
rect 487982 166948 487988 167000
rect 488040 166988 488046 167000
rect 580166 166988 580172 167000
rect 488040 166960 580172 166988
rect 488040 166948 488046 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 3418 164160 3424 164212
rect 3476 164200 3482 164212
rect 39298 164200 39304 164212
rect 3476 164172 39304 164200
rect 3476 164160 3482 164172
rect 39298 164160 39304 164172
rect 39356 164160 39362 164212
rect 3418 111732 3424 111784
rect 3476 111772 3482 111784
rect 43438 111772 43444 111784
rect 3476 111744 43444 111772
rect 3476 111732 3482 111744
rect 43438 111732 43444 111744
rect 43496 111732 43502 111784
rect 73062 87252 73068 87304
rect 73120 87292 73126 87304
rect 291838 87292 291844 87304
rect 73120 87264 291844 87292
rect 73120 87252 73126 87264
rect 291838 87252 291844 87264
rect 291896 87252 291902 87304
rect 70118 87184 70124 87236
rect 70176 87224 70182 87236
rect 85022 87224 85028 87236
rect 70176 87196 85028 87224
rect 70176 87184 70182 87196
rect 85022 87184 85028 87196
rect 85080 87184 85086 87236
rect 74442 87116 74448 87168
rect 74500 87156 74506 87168
rect 98730 87156 98736 87168
rect 74500 87128 98736 87156
rect 74500 87116 74506 87128
rect 98730 87116 98736 87128
rect 98788 87116 98794 87168
rect 76466 87048 76472 87100
rect 76524 87088 76530 87100
rect 289078 87088 289084 87100
rect 76524 87060 289084 87088
rect 76524 87048 76530 87060
rect 289078 87048 289084 87060
rect 289136 87048 289142 87100
rect 81158 86980 81164 87032
rect 81216 87020 81222 87032
rect 84838 87020 84844 87032
rect 81216 86992 84844 87020
rect 81216 86980 81222 86992
rect 84838 86980 84844 86992
rect 84896 86980 84902 87032
rect 487890 86912 487896 86964
rect 487948 86952 487954 86964
rect 580166 86952 580172 86964
rect 487948 86924 580172 86952
rect 487948 86912 487954 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 85022 83444 85028 83496
rect 85080 83484 85086 83496
rect 339862 83484 339868 83496
rect 85080 83456 339868 83484
rect 85080 83444 85086 83456
rect 339862 83444 339868 83456
rect 339920 83444 339926 83496
rect 84838 79296 84844 79348
rect 84896 79336 84902 79348
rect 364610 79336 364616 79348
rect 84896 79308 364616 79336
rect 84896 79296 84902 79308
rect 364610 79296 364616 79308
rect 364668 79296 364674 79348
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 15838 71720 15844 71732
rect 3476 71692 15844 71720
rect 3476 71680 3482 71692
rect 15838 71680 15844 71692
rect 15896 71680 15902 71732
rect 98730 51688 98736 51740
rect 98788 51728 98794 51740
rect 350442 51728 350448 51740
rect 98788 51700 350448 51728
rect 98788 51688 98794 51700
rect 350442 51688 350448 51700
rect 350500 51688 350506 51740
rect 511258 46860 511264 46912
rect 511316 46900 511322 46912
rect 580166 46900 580172 46912
rect 511316 46872 580172 46900
rect 511316 46860 511322 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3418 33056 3424 33108
rect 3476 33096 3482 33108
rect 11698 33096 11704 33108
rect 3476 33068 11704 33096
rect 3476 33056 3482 33068
rect 11698 33056 11704 33068
rect 11756 33056 11762 33108
rect 289078 7556 289084 7608
rect 289136 7596 289142 7608
rect 354030 7596 354036 7608
rect 289136 7568 354036 7596
rect 289136 7556 289142 7568
rect 354030 7556 354036 7568
rect 354088 7556 354094 7608
rect 287698 6808 287704 6860
rect 287756 6848 287762 6860
rect 580166 6848 580172 6860
rect 287756 6820 580172 6848
rect 287756 6808 287762 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 291838 4768 291844 4820
rect 291896 4808 291902 4820
rect 346946 4808 346952 4820
rect 291896 4780 346952 4808
rect 291896 4768 291902 4780
rect 346946 4768 346952 4780
rect 347004 4768 347010 4820
rect 243538 4088 243544 4140
rect 243596 4128 243602 4140
rect 288526 4128 288532 4140
rect 243596 4100 288532 4128
rect 243596 4088 243602 4100
rect 288526 4088 288532 4100
rect 288584 4088 288590 4140
rect 271782 4020 271788 4072
rect 271840 4060 271846 4072
rect 283834 4060 283840 4072
rect 271840 4032 283840 4060
rect 271840 4020 271846 4032
rect 283834 4020 283840 4032
rect 283892 4020 283898 4072
rect 446398 3408 446404 3460
rect 446456 3448 446462 3460
rect 583386 3448 583392 3460
rect 446456 3420 583392 3448
rect 446456 3408 446462 3420
rect 583386 3408 583392 3420
rect 583444 3408 583450 3460
rect 442902 2796 442908 2848
rect 442960 2836 442966 2848
rect 580994 2836 581000 2848
rect 442960 2808 581000 2836
rect 442960 2796 442966 2808
rect 580994 2796 581000 2808
rect 581052 2796 581058 2848
<< via1 >>
rect 485044 700272 485096 700324
rect 527180 700272 527232 700324
rect 3424 683136 3476 683188
rect 87604 683136 87656 683188
rect 487804 657500 487856 657552
rect 534908 657500 534960 657552
rect 487896 657432 487948 657484
rect 537668 657432 537720 657484
rect 486884 657364 486936 657416
rect 496268 657364 496320 657416
rect 503168 657364 503220 657416
rect 580448 657364 580500 657416
rect 487160 657296 487212 657348
rect 497648 657296 497700 657348
rect 505100 657296 505152 657348
rect 530768 657296 530820 657348
rect 490380 657228 490432 657280
rect 529388 657228 529440 657280
rect 490472 657160 490524 657212
rect 533528 657160 533580 657212
rect 489184 657092 489236 657144
rect 532148 657092 532200 657144
rect 488448 657024 488500 657076
rect 494888 657024 494940 657076
rect 487068 656956 487120 657008
rect 493508 656956 493560 657008
rect 486976 656888 487028 656940
rect 492128 656888 492180 656940
rect 494704 656888 494756 656940
rect 504548 656888 504600 656940
rect 514760 656888 514812 656940
rect 526628 656888 526680 656940
rect 224960 656140 225012 656192
rect 503168 656140 503220 656192
rect 504548 655732 504600 655784
rect 580632 655732 580684 655784
rect 500408 655664 500460 655716
rect 577504 655664 577556 655716
rect 489276 655596 489328 655648
rect 499028 655596 499080 655648
rect 501788 655596 501840 655648
rect 580356 655596 580408 655648
rect 237656 655528 237708 655580
rect 528008 655528 528060 655580
rect 231584 654780 231636 654832
rect 514760 654780 514812 654832
rect 274548 654508 274600 654560
rect 536012 654508 536064 654560
rect 286968 654440 287020 654492
rect 538772 654440 538824 654492
rect 243728 650632 243780 650684
rect 490380 650632 490432 650684
rect 255964 647844 256016 647896
rect 489184 647844 489236 647896
rect 577596 643084 577648 643136
rect 580724 643084 580776 643136
rect 281448 642336 281500 642388
rect 487896 642336 487948 642388
rect 86868 633360 86920 633412
rect 486976 633360 487028 633412
rect 88248 632884 88300 632936
rect 255964 632884 256016 632936
rect 98000 632816 98052 632868
rect 486884 632816 486936 632868
rect 91100 632748 91152 632800
rect 91928 632748 91980 632800
rect 488448 632748 488500 632800
rect 54300 632272 54352 632324
rect 85856 632680 85908 632732
rect 487068 632680 487120 632732
rect 286232 632272 286284 632324
rect 286968 632272 287020 632324
rect 294144 632272 294196 632324
rect 486884 632272 486936 632324
rect 488080 632272 488132 632324
rect 55956 632204 56008 632256
rect 91100 632204 91152 632256
rect 280160 632204 280212 632256
rect 281448 632204 281500 632256
rect 293040 632204 293092 632256
rect 487068 632204 487120 632256
rect 487988 632204 488040 632256
rect 57612 632136 57664 632188
rect 98000 632136 98052 632188
rect 274548 632136 274600 632188
rect 294328 632136 294380 632188
rect 486976 632136 487028 632188
rect 487896 632136 487948 632188
rect 488448 632136 488500 632188
rect 489184 632136 489236 632188
rect 50988 632068 51040 632120
rect 73712 632068 73764 632120
rect 490564 632068 490616 632120
rect 65892 630640 65944 630692
rect 128820 630640 128872 630692
rect 62764 629620 62816 629672
rect 115940 629620 115992 629672
rect 64420 629552 64472 629604
rect 122012 629552 122064 629604
rect 68928 629484 68980 629536
rect 231308 629484 231360 629536
rect 67456 629416 67508 629468
rect 237380 629416 237432 629468
rect 67548 629348 67600 629400
rect 243452 629348 243504 629400
rect 67456 629280 67508 629332
rect 134156 629280 134208 629332
rect 490564 594056 490616 594108
rect 511264 594056 511316 594108
rect 3424 527144 3476 527196
rect 60740 527144 60792 527196
rect 227720 478796 227772 478848
rect 544108 478796 544160 478848
rect 231768 478728 231820 478780
rect 294144 478728 294196 478780
rect 233148 478660 233200 478712
rect 293040 478660 293092 478712
rect 241428 478592 241480 478644
rect 294328 478592 294380 478644
rect 231492 478320 231544 478372
rect 540152 478320 540204 478372
rect 234344 478252 234396 478304
rect 543004 478252 543056 478304
rect 231676 478184 231728 478236
rect 580540 478184 580592 478236
rect 230112 478116 230164 478168
rect 580632 478116 580684 478168
rect 68468 477640 68520 477692
rect 126244 477640 126296 477692
rect 68100 477572 68152 477624
rect 138664 477572 138716 477624
rect 68192 477504 68244 477556
rect 142896 477504 142948 477556
rect 3424 476008 3476 476060
rect 62120 476008 62172 476060
rect 243544 476008 243596 476060
rect 542728 476008 542780 476060
rect 251088 475940 251140 475992
rect 508688 475940 508740 475992
rect 231860 475872 231912 475924
rect 485044 475872 485096 475924
rect 262864 475804 262916 475856
rect 507308 475804 507360 475856
rect 271788 475736 271840 475788
rect 505928 475736 505980 475788
rect 233884 475668 233936 475720
rect 462320 475668 462372 475720
rect 235632 475396 235684 475448
rect 542636 475396 542688 475448
rect 62120 475328 62172 475380
rect 63224 475328 63276 475380
rect 94044 475328 94096 475380
rect 233056 475328 233108 475380
rect 577596 475328 577648 475380
rect 231400 474308 231452 474360
rect 231676 474308 231728 474360
rect 230296 473288 230348 473340
rect 544200 473288 544252 473340
rect 230388 473220 230440 473272
rect 544016 473220 544068 473272
rect 238484 473152 238536 473204
rect 541164 473152 541216 473204
rect 247040 473084 247092 473136
rect 526628 473084 526680 473136
rect 255320 473016 255372 473068
rect 525248 473016 525300 473068
rect 232780 472608 232832 472660
rect 539048 472608 539100 472660
rect 230020 471860 230072 471912
rect 230296 471860 230348 471912
rect 240048 443028 240100 443080
rect 288716 443028 288768 443080
rect 237380 442960 237432 443012
rect 288624 442960 288676 443012
rect 69664 442892 69716 442944
rect 70216 442892 70268 442944
rect 233976 442892 234028 442944
rect 488172 442892 488224 442944
rect 277216 442348 277268 442400
rect 289452 442348 289504 442400
rect 238484 442280 238536 442332
rect 541072 442280 541124 442332
rect 69664 442212 69716 442264
rect 489276 442212 489328 442264
rect 229008 442144 229060 442196
rect 288808 442144 288860 442196
rect 223488 442076 223540 442128
rect 267740 442076 267792 442128
rect 270408 442076 270460 442128
rect 284484 442076 284536 442128
rect 240048 442008 240100 442060
rect 242808 442008 242860 442060
rect 254032 442008 254084 442060
rect 280436 442008 280488 442060
rect 253940 441940 253992 441992
rect 280712 441940 280764 441992
rect 251088 441872 251140 441924
rect 282920 441872 282972 441924
rect 264980 441804 265032 441856
rect 281080 441804 281132 441856
rect 239864 441736 239916 441788
rect 289728 441736 289780 441788
rect 239220 441668 239272 441720
rect 289636 441668 289688 441720
rect 273260 441600 273312 441652
rect 284392 441600 284444 441652
rect 267740 441532 267792 441584
rect 474740 441532 474792 441584
rect 238392 440988 238444 441040
rect 539876 440988 539928 441040
rect 238208 440920 238260 440972
rect 539692 440920 539744 440972
rect 238116 440852 238168 440904
rect 540980 440852 541032 440904
rect 240784 440716 240836 440768
rect 287704 440716 287756 440768
rect 232688 440648 232740 440700
rect 282092 440648 282144 440700
rect 230480 440580 230532 440632
rect 281080 440580 281132 440632
rect 231400 440512 231452 440564
rect 282000 440512 282052 440564
rect 229652 440444 229704 440496
rect 280988 440444 281040 440496
rect 228916 440376 228968 440428
rect 280252 440376 280304 440428
rect 229008 440308 229060 440360
rect 280528 440308 280580 440360
rect 221464 440240 221516 440292
rect 223488 440240 223540 440292
rect 227168 440240 227220 440292
rect 284300 440240 284352 440292
rect 474740 440240 474792 440292
rect 475384 440240 475436 440292
rect 229376 439832 229428 439884
rect 230020 439832 230072 439884
rect 239772 439696 239824 439748
rect 580264 439696 580316 439748
rect 228732 439628 228784 439680
rect 280160 439628 280212 439680
rect 229008 439560 229060 439612
rect 280620 439560 280672 439612
rect 231400 439492 231452 439544
rect 280068 439492 280120 439544
rect 229652 439424 229704 439476
rect 280896 439424 280948 439476
rect 231032 439356 231084 439408
rect 281816 439356 281868 439408
rect 228272 439084 228324 439136
rect 228732 439084 228784 439136
rect 218060 438880 218112 438932
rect 221464 438880 221516 438932
rect 239220 436772 239272 436824
rect 239772 436772 239824 436824
rect 280896 436500 280948 436552
rect 281080 436500 281132 436552
rect 281632 435548 281684 435600
rect 282092 435548 282144 435600
rect 213552 434664 213604 434716
rect 218060 434732 218112 434784
rect 281540 434188 281592 434240
rect 282000 434188 282052 434240
rect 211620 430584 211672 430636
rect 213552 430584 213604 430636
rect 3424 423580 3476 423632
rect 60740 423580 60792 423632
rect 60740 422900 60792 422952
rect 61844 422900 61896 422952
rect 95700 422900 95752 422952
rect 207020 422288 207072 422340
rect 211620 422288 211672 422340
rect 202880 418072 202932 418124
rect 207020 418140 207072 418192
rect 198832 412632 198884 412684
rect 202788 412632 202840 412684
rect 281908 409776 281960 409828
rect 284484 409776 284536 409828
rect 198004 408484 198056 408536
rect 198832 408484 198884 408536
rect 281908 408416 281960 408468
rect 284392 408416 284444 408468
rect 577504 405628 577556 405680
rect 579712 405628 579764 405680
rect 193864 400120 193916 400172
rect 198004 400188 198056 400240
rect 281816 394612 281868 394664
rect 284300 394612 284352 394664
rect 191840 386316 191892 386368
rect 193864 386316 193916 386368
rect 192484 383664 192536 383716
rect 237380 383664 237432 383716
rect 216036 382372 216088 382424
rect 237380 382508 237432 382560
rect 112536 382304 112588 382356
rect 237380 382304 237432 382356
rect 112444 382236 112496 382288
rect 237472 382236 237524 382288
rect 112720 380944 112772 380996
rect 237564 380944 237616 380996
rect 111156 380876 111208 380928
rect 237380 380876 237432 380928
rect 110052 379516 110104 379568
rect 237380 379516 237432 379568
rect 186964 379448 187016 379500
rect 191748 379448 191800 379500
rect 127624 376864 127676 376916
rect 237380 376864 237432 376916
rect 123576 376796 123628 376848
rect 237564 376796 237616 376848
rect 111524 376728 111576 376780
rect 237748 376728 237800 376780
rect 126428 375436 126480 375488
rect 237380 375436 237432 375488
rect 111616 375368 111668 375420
rect 237564 375368 237616 375420
rect 122196 374076 122248 374128
rect 237380 374280 237432 374332
rect 115296 374008 115348 374060
rect 237380 374008 237432 374060
rect 3424 372512 3476 372564
rect 63500 372512 63552 372564
rect 63500 371832 63552 371884
rect 64604 371832 64656 371884
rect 97356 371832 97408 371884
rect 137284 371220 137336 371272
rect 237380 371220 237432 371272
rect 115388 369860 115440 369912
rect 237380 369860 237432 369912
rect 282828 368500 282880 368552
rect 287152 368500 287204 368552
rect 489276 366324 489328 366376
rect 498844 366324 498896 366376
rect 282828 358776 282880 358828
rect 288992 358776 289044 358828
rect 185584 358708 185636 358760
rect 186964 358708 187016 358760
rect 282828 356056 282880 356108
rect 287244 356056 287296 356108
rect 282828 353268 282880 353320
rect 289084 353268 289136 353320
rect 498844 353200 498896 353252
rect 580172 353200 580224 353252
rect 60924 352520 60976 352572
rect 69664 352520 69716 352572
rect 282828 347760 282880 347812
rect 291292 347760 291344 347812
rect 182180 347692 182232 347744
rect 185584 347692 185636 347744
rect 59084 344292 59136 344344
rect 182180 344292 182232 344344
rect 475384 344292 475436 344344
rect 497464 344292 497516 344344
rect 216680 343612 216732 343664
rect 235264 343612 235316 343664
rect 282828 343612 282880 343664
rect 287336 343612 287388 343664
rect 63592 342524 63644 342576
rect 86960 342524 87012 342576
rect 66168 342456 66220 342508
rect 92020 342456 92072 342508
rect 43444 342388 43496 342440
rect 105268 342388 105320 342440
rect 15844 342320 15896 342372
rect 106924 342320 106976 342372
rect 11704 342252 11756 342304
rect 108304 342252 108356 342304
rect 99380 341776 99432 341828
rect 100300 341776 100352 341828
rect 65800 341300 65852 341352
rect 228824 341300 228876 341352
rect 39304 341232 39356 341284
rect 104164 341232 104216 341284
rect 215944 341232 215996 341284
rect 237564 341232 237616 341284
rect 25504 341164 25556 341216
rect 99380 341164 99432 341216
rect 213184 341164 213236 341216
rect 237380 341164 237432 341216
rect 70216 341096 70268 341148
rect 225880 341096 225932 341148
rect 70308 341028 70360 341080
rect 228640 341028 228692 341080
rect 67456 340960 67508 341012
rect 228548 340960 228600 341012
rect 228364 340892 228416 340944
rect 237380 340892 237432 340944
rect 43536 339532 43588 339584
rect 102140 339532 102192 339584
rect 29644 339464 29696 339516
rect 98644 339464 98696 339516
rect 3424 320084 3476 320136
rect 29644 320084 29696 320136
rect 235264 300772 235316 300824
rect 237380 300772 237432 300824
rect 497464 299412 497516 299464
rect 580172 299412 580224 299464
rect 282828 295332 282880 295384
rect 288532 295332 288584 295384
rect 142896 288328 142948 288380
rect 237380 288328 237432 288380
rect 126244 286968 126296 287020
rect 237380 286968 237432 287020
rect 138664 285608 138716 285660
rect 237380 285608 237432 285660
rect 225880 282820 225932 282872
rect 237380 282820 237432 282872
rect 228824 281460 228876 281512
rect 237564 281460 237616 281512
rect 282828 281460 282880 281512
rect 288808 281460 288860 281512
rect 228640 281392 228692 281444
rect 237380 281392 237432 281444
rect 78956 280100 79008 280152
rect 126428 280100 126480 280152
rect 228548 280100 228600 280152
rect 237380 280100 237432 280152
rect 80060 280032 80112 280084
rect 127624 280032 127676 280084
rect 78588 279964 78640 280016
rect 122196 279964 122248 280016
rect 81440 279896 81492 279948
rect 111616 279896 111668 279948
rect 96528 279828 96580 279880
rect 123576 279828 123628 279880
rect 99380 279760 99432 279812
rect 111524 279760 111576 279812
rect 98644 278672 98696 278724
rect 111156 278672 111208 278724
rect 97908 278604 97960 278656
rect 110052 278604 110104 278656
rect 89720 278536 89772 278588
rect 137284 278536 137336 278588
rect 91100 278468 91152 278520
rect 115388 278468 115440 278520
rect 95148 278400 95200 278452
rect 115296 278400 115348 278452
rect 102140 278332 102192 278384
rect 106188 278332 106240 278384
rect 112444 278332 112496 278384
rect 112536 278332 112588 278384
rect 104808 278196 104860 278248
rect 112720 278196 112772 278248
rect 107384 278128 107436 278180
rect 216036 278128 216088 278180
rect 108304 278060 108356 278112
rect 192484 278060 192536 278112
rect 282828 274592 282880 274644
rect 288716 274592 288768 274644
rect 282828 273164 282880 273216
rect 288624 273164 288676 273216
rect 3424 267656 3476 267708
rect 25504 267656 25556 267708
rect 488080 245556 488132 245608
rect 580172 245556 580224 245608
rect 284852 243516 284904 243568
rect 285128 243516 285180 243568
rect 284484 243380 284536 243432
rect 284852 243380 284904 243432
rect 186320 240048 186372 240100
rect 282368 240048 282420 240100
rect 212448 239980 212500 240032
rect 287336 239980 287388 240032
rect 236000 239912 236052 239964
rect 291292 239912 291344 239964
rect 237472 239844 237524 239896
rect 289084 239844 289136 239896
rect 237564 239776 237616 239828
rect 287244 239776 287296 239828
rect 237380 239708 237432 239760
rect 280896 239708 280948 239760
rect 259276 239640 259328 239692
rect 288992 239640 289044 239692
rect 264980 239572 265032 239624
rect 287152 239572 287204 239624
rect 179420 239368 179472 239420
rect 284484 239368 284536 239420
rect 44180 238688 44232 238740
rect 243820 238688 243872 238740
rect 121460 238620 121512 238672
rect 245016 238620 245068 238672
rect 3424 215228 3476 215280
rect 43536 215228 43588 215280
rect 489184 206932 489236 206984
rect 580172 206932 580224 206984
rect 487988 166948 488040 167000
rect 580172 166948 580224 167000
rect 3424 164160 3476 164212
rect 39304 164160 39356 164212
rect 3424 111732 3476 111784
rect 43444 111732 43496 111784
rect 73068 87252 73120 87304
rect 291844 87252 291896 87304
rect 70124 87184 70176 87236
rect 85028 87184 85080 87236
rect 74448 87116 74500 87168
rect 98736 87116 98788 87168
rect 76472 87048 76524 87100
rect 289084 87048 289136 87100
rect 81164 86980 81216 87032
rect 84844 86980 84896 87032
rect 487896 86912 487948 86964
rect 580172 86912 580224 86964
rect 85028 83444 85080 83496
rect 339868 83444 339920 83496
rect 84844 79296 84896 79348
rect 364616 79296 364668 79348
rect 3424 71680 3476 71732
rect 15844 71680 15896 71732
rect 98736 51688 98788 51740
rect 350448 51688 350500 51740
rect 511264 46860 511316 46912
rect 580172 46860 580224 46912
rect 3424 33056 3476 33108
rect 11704 33056 11756 33108
rect 289084 7556 289136 7608
rect 354036 7556 354088 7608
rect 287704 6808 287756 6860
rect 580172 6808 580224 6860
rect 291844 4768 291896 4820
rect 346952 4768 347004 4820
rect 243544 4088 243596 4140
rect 288532 4088 288584 4140
rect 271788 4020 271840 4072
rect 283840 4020 283892 4072
rect 446404 3408 446456 3460
rect 583392 3408 583444 3460
rect 442908 2796 442960 2848
rect 581000 2796 581052 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 4066 553480 4122 553489
rect 4066 553415 4122 553424
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3974 502344 4030 502353
rect 3974 502279 4030 502288
rect 3424 476060 3476 476066
rect 3424 476002 3476 476008
rect 3436 475697 3464 476002
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3988 474065 4016 502279
rect 3974 474056 4030 474065
rect 3974 473991 4030 474000
rect 4080 453393 4108 553415
rect 4066 453384 4122 453393
rect 4066 453319 4122 453328
rect 3424 423632 3476 423638
rect 3422 423600 3424 423609
rect 3476 423600 3478 423609
rect 3422 423535 3478 423544
rect 3424 372564 3476 372570
rect 3424 372506 3476 372512
rect 3436 371385 3464 372506
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 8128 364993 8156 703520
rect 24320 700505 24348 703520
rect 24306 700496 24362 700505
rect 24306 700431 24362 700440
rect 40512 700369 40540 703520
rect 60002 700496 60058 700505
rect 60002 700431 60058 700440
rect 40498 700360 40554 700369
rect 40498 700295 40554 700304
rect 54300 632324 54352 632330
rect 54300 632266 54352 632272
rect 52642 632224 52698 632233
rect 52642 632159 52698 632168
rect 50988 632120 51040 632126
rect 50988 632062 51040 632068
rect 48134 442504 48190 442513
rect 48134 442439 48190 442448
rect 8114 364984 8170 364993
rect 8114 364919 8170 364928
rect 5262 349208 5318 349217
rect 5262 349143 5318 349152
rect 3424 320136 3476 320142
rect 3424 320078 3476 320084
rect 3436 319297 3464 320078
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3424 267708 3476 267714
rect 3424 267650 3476 267656
rect 3436 267209 3464 267650
rect 3422 267200 3478 267209
rect 3422 267135 3478 267144
rect 3424 215280 3476 215286
rect 3424 215222 3476 215228
rect 3436 214985 3464 215222
rect 3422 214976 3478 214985
rect 3422 214911 3478 214920
rect 3424 164212 3476 164218
rect 3424 164154 3476 164160
rect 3436 162897 3464 164154
rect 3422 162888 3478 162897
rect 3422 162823 3478 162832
rect 3424 111784 3476 111790
rect 3424 111726 3476 111732
rect 3436 110673 3464 111726
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 4066 94480 4122 94489
rect 4066 94415 4122 94424
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 570 51776 626 51785
rect 570 51711 626 51720
rect 584 480 612 51711
rect 3424 33108 3476 33114
rect 3424 33050 3476 33056
rect 3436 32473 3464 33050
rect 3422 32464 3478 32473
rect 3422 32399 3478 32408
rect 2870 18864 2926 18873
rect 2870 18799 2926 18808
rect 1674 4040 1730 4049
rect 1674 3975 1730 3984
rect 1688 480 1716 3975
rect 2884 480 2912 18799
rect 4080 480 4108 94415
rect 5276 480 5304 349143
rect 6458 348120 6514 348129
rect 6458 348055 6514 348064
rect 6472 480 6500 348055
rect 43444 342440 43496 342446
rect 43444 342382 43496 342388
rect 15844 342372 15896 342378
rect 15844 342314 15896 342320
rect 11704 342304 11756 342310
rect 11704 342246 11756 342252
rect 8758 95840 8814 95849
rect 8758 95775 8814 95784
rect 7562 40896 7618 40905
rect 7562 40831 7618 40840
rect 7576 4049 7604 40831
rect 7654 4992 7710 5001
rect 7654 4927 7710 4936
rect 7562 4040 7618 4049
rect 7562 3975 7618 3984
rect 7668 480 7696 4927
rect 8772 480 8800 95775
rect 11716 33114 11744 342246
rect 14738 235376 14794 235385
rect 14738 235311 14794 235320
rect 11704 33108 11756 33114
rect 11704 33050 11756 33056
rect 12346 6216 12402 6225
rect 12346 6151 12402 6160
rect 9954 3360 10010 3369
rect 9954 3295 10010 3304
rect 9968 480 9996 3295
rect 12360 480 12388 6151
rect 13542 3632 13598 3641
rect 13542 3567 13598 3576
rect 13556 480 13584 3567
rect 14752 480 14780 235311
rect 15856 71738 15884 342314
rect 39304 341284 39356 341290
rect 39304 341226 39356 341232
rect 25504 341216 25556 341222
rect 25504 341158 25556 341164
rect 18234 269784 18290 269793
rect 18234 269719 18290 269728
rect 17038 237552 17094 237561
rect 17038 237487 17094 237496
rect 15844 71732 15896 71738
rect 15844 71674 15896 71680
rect 17052 480 17080 237487
rect 18248 480 18276 269719
rect 23018 268424 23074 268433
rect 23018 268359 23074 268368
rect 21822 237416 21878 237425
rect 21822 237351 21878 237360
rect 19430 2952 19486 2961
rect 19430 2887 19486 2896
rect 19444 480 19472 2887
rect 21836 480 21864 237351
rect 23032 480 23060 268359
rect 25516 267714 25544 341158
rect 29644 339516 29696 339522
rect 29644 339458 29696 339464
rect 29656 320142 29684 339458
rect 29644 320136 29696 320142
rect 29644 320078 29696 320084
rect 25504 267708 25556 267714
rect 25504 267650 25556 267656
rect 31298 264208 31354 264217
rect 31298 264143 31354 264152
rect 30102 238096 30158 238105
rect 30102 238031 30158 238040
rect 26514 237960 26570 237969
rect 26514 237895 26570 237904
rect 24214 225584 24270 225593
rect 24214 225519 24270 225528
rect 24228 480 24256 225519
rect 25502 218648 25558 218657
rect 25502 218583 25558 218592
rect 25516 3369 25544 218583
rect 25502 3360 25558 3369
rect 25502 3295 25558 3304
rect 26528 480 26556 237895
rect 27710 102776 27766 102785
rect 27710 102711 27766 102720
rect 27724 480 27752 102711
rect 28906 3496 28962 3505
rect 28906 3431 28962 3440
rect 28920 480 28948 3431
rect 30116 480 30144 238031
rect 31312 480 31340 264143
rect 34794 244896 34850 244905
rect 34794 244831 34850 244840
rect 33598 238232 33654 238241
rect 33598 238167 33654 238176
rect 32402 203552 32458 203561
rect 32402 203487 32458 203496
rect 32416 3505 32444 203487
rect 32402 3496 32458 3505
rect 32402 3431 32458 3440
rect 32402 2816 32458 2825
rect 32402 2751 32458 2760
rect 32416 480 32444 2751
rect 33612 480 33640 238167
rect 34808 480 34836 244831
rect 35990 238776 36046 238785
rect 35990 238711 36046 238720
rect 36004 480 36032 238711
rect 37186 238368 37242 238377
rect 37186 238303 37242 238312
rect 37200 480 37228 238303
rect 39316 164218 39344 341226
rect 40682 238504 40738 238513
rect 40682 238439 40738 238448
rect 39578 233880 39634 233889
rect 39578 233815 39634 233824
rect 39304 164212 39356 164218
rect 39304 164154 39356 164160
rect 38382 104136 38438 104145
rect 38382 104071 38438 104080
rect 38396 480 38424 104071
rect 39592 480 39620 233815
rect 40696 480 40724 238439
rect 43074 228304 43130 228313
rect 43074 228239 43130 228248
rect 41878 105496 41934 105505
rect 41878 105431 41934 105440
rect 41892 480 41920 105431
rect 43088 480 43116 228239
rect 43456 111790 43484 342382
rect 43536 339584 43588 339590
rect 43536 339526 43588 339532
rect 43548 215286 43576 339526
rect 48148 325009 48176 442439
rect 50618 367704 50674 367713
rect 50618 367639 50674 367648
rect 48226 340096 48282 340105
rect 48226 340031 48282 340040
rect 48134 325000 48190 325009
rect 48134 324935 48190 324944
rect 48240 295089 48268 340031
rect 48226 295080 48282 295089
rect 48226 295015 48282 295024
rect 44180 238740 44232 238746
rect 44180 238682 44232 238688
rect 44192 237561 44220 238682
rect 44270 238640 44326 238649
rect 44270 238575 44326 238584
rect 44178 237552 44234 237561
rect 44178 237487 44234 237496
rect 43536 215280 43588 215286
rect 43536 215222 43588 215228
rect 43444 111784 43496 111790
rect 43444 111726 43496 111732
rect 44284 480 44312 238575
rect 46662 174584 46718 174593
rect 46662 174519 46718 174528
rect 45466 106856 45522 106865
rect 45466 106791 45522 106800
rect 45480 480 45508 106791
rect 46676 480 46704 174519
rect 48042 81696 48098 81705
rect 48042 81631 48098 81640
rect 47582 64016 47638 64025
rect 47582 63951 47638 63960
rect 47490 57216 47546 57225
rect 47490 57151 47546 57160
rect 47504 18601 47532 57151
rect 47596 19961 47624 63951
rect 47950 62656 48006 62665
rect 47950 62591 48006 62600
rect 47858 61296 47914 61305
rect 47858 61231 47914 61240
rect 47766 59936 47822 59945
rect 47766 59871 47822 59880
rect 47674 58576 47730 58585
rect 47674 58511 47730 58520
rect 47688 28257 47716 58511
rect 47674 28248 47730 28257
rect 47674 28183 47730 28192
rect 47780 26897 47808 59871
rect 47766 26888 47822 26897
rect 47766 26823 47822 26832
rect 47872 24177 47900 61231
rect 47858 24168 47914 24177
rect 47858 24103 47914 24112
rect 47964 22681 47992 62591
rect 48056 42265 48084 81631
rect 48134 80336 48190 80345
rect 48134 80271 48190 80280
rect 48148 49065 48176 80271
rect 48240 51513 48268 295015
rect 50632 280786 50660 367639
rect 51000 340218 51028 632062
rect 52656 340218 52684 632159
rect 54312 340218 54340 632266
rect 55956 632256 56008 632262
rect 55956 632198 56008 632204
rect 55968 340218 55996 632198
rect 57612 632188 57664 632194
rect 57612 632130 57664 632136
rect 57624 340218 57652 632130
rect 60016 444145 60044 700431
rect 69938 633176 69994 633185
rect 69938 633111 69994 633120
rect 69846 632904 69902 632913
rect 69846 632839 69902 632848
rect 64786 632632 64842 632641
rect 64786 632567 64842 632576
rect 60646 632088 60702 632097
rect 60646 632023 60702 632032
rect 60554 580000 60610 580009
rect 60554 579935 60610 579944
rect 60568 579601 60596 579935
rect 60554 579592 60610 579601
rect 60554 579527 60610 579536
rect 60002 444136 60058 444145
rect 60002 444071 60058 444080
rect 59084 344344 59136 344350
rect 59084 344286 59136 344292
rect 50954 340190 51028 340218
rect 52610 340190 52684 340218
rect 54266 340190 54340 340218
rect 55922 340190 55996 340218
rect 57578 340190 57652 340218
rect 50954 339932 50982 340190
rect 52610 339932 52638 340190
rect 54266 339932 54294 340190
rect 55922 339932 55950 340190
rect 57578 339932 57606 340190
rect 59096 339674 59124 344286
rect 60568 342961 60596 579527
rect 60660 343097 60688 632023
rect 62026 631544 62082 631553
rect 62026 631479 62082 631488
rect 61934 629776 61990 629785
rect 61934 629711 61990 629720
rect 61842 629640 61898 629649
rect 61842 629575 61898 629584
rect 60738 527232 60794 527241
rect 60738 527167 60740 527176
rect 60792 527167 60794 527176
rect 61750 527232 61806 527241
rect 61750 527167 61806 527176
rect 60740 527138 60792 527144
rect 60740 423632 60792 423638
rect 60740 423574 60792 423580
rect 60752 422958 60780 423574
rect 60740 422952 60792 422958
rect 60740 422894 60792 422900
rect 60924 352572 60976 352578
rect 60924 352514 60976 352520
rect 60646 343088 60702 343097
rect 60646 343023 60702 343032
rect 60554 342952 60610 342961
rect 60554 342887 60610 342896
rect 60936 340218 60964 352514
rect 61764 343641 61792 527167
rect 61856 422958 61884 629575
rect 61844 422952 61896 422958
rect 61844 422894 61896 422900
rect 61750 343632 61806 343641
rect 61750 343567 61806 343576
rect 61948 343233 61976 629711
rect 62040 344185 62068 631479
rect 63406 631272 63462 631281
rect 63406 631207 63462 631216
rect 63222 630320 63278 630329
rect 63222 630255 63278 630264
rect 63130 630184 63186 630193
rect 63130 630119 63186 630128
rect 62764 629672 62816 629678
rect 62764 629614 62816 629620
rect 62776 625154 62804 629614
rect 62592 625126 62804 625154
rect 62120 476060 62172 476066
rect 62120 476002 62172 476008
rect 62132 475386 62160 476002
rect 62120 475380 62172 475386
rect 62120 475322 62172 475328
rect 62026 344176 62082 344185
rect 62026 344111 62082 344120
rect 61934 343224 61990 343233
rect 61934 343159 61990 343168
rect 62592 340218 62620 625126
rect 63144 342689 63172 630119
rect 63236 475386 63264 630255
rect 63224 475380 63276 475386
rect 63224 475322 63276 475328
rect 63420 343482 63448 631207
rect 64694 629912 64750 629921
rect 64694 629847 64750 629856
rect 64420 629604 64472 629610
rect 64420 629546 64472 629552
rect 64432 625154 64460 629546
rect 64602 629504 64658 629513
rect 64602 629439 64658 629448
rect 64248 625126 64460 625154
rect 63500 372564 63552 372570
rect 63500 372506 63552 372512
rect 63512 371890 63540 372506
rect 63500 371884 63552 371890
rect 63500 371826 63552 371832
rect 63420 343454 63632 343482
rect 63130 342680 63186 342689
rect 63130 342615 63186 342624
rect 63604 342582 63632 343454
rect 63592 342576 63644 342582
rect 63592 342518 63644 342524
rect 64248 340218 64276 625126
rect 64616 371890 64644 629439
rect 64604 371884 64656 371890
rect 64604 371826 64656 371832
rect 64708 343505 64736 629847
rect 64694 343496 64750 343505
rect 64694 343431 64750 343440
rect 64800 342825 64828 632567
rect 66074 632496 66130 632505
rect 66074 632431 66130 632440
rect 65892 630692 65944 630698
rect 65892 630634 65944 630640
rect 65798 492688 65854 492697
rect 65798 492623 65854 492632
rect 64786 342816 64842 342825
rect 64786 342751 64842 342760
rect 65812 341358 65840 492623
rect 65800 341352 65852 341358
rect 65800 341294 65852 341300
rect 65904 340218 65932 630634
rect 65982 629368 66038 629377
rect 65982 629303 66038 629312
rect 65996 478145 66024 629303
rect 65982 478136 66038 478145
rect 65982 478071 66038 478080
rect 66088 477873 66116 632431
rect 66166 631408 66222 631417
rect 66166 631343 66222 631352
rect 66180 629354 66208 631343
rect 69202 630864 69258 630873
rect 69202 630799 69258 630808
rect 68926 630320 68982 630329
rect 68926 630255 68982 630264
rect 67362 630048 67418 630057
rect 67362 629983 67418 629992
rect 66902 629368 66958 629377
rect 66180 629326 66300 629354
rect 66272 629082 66300 629326
rect 66902 629303 66958 629312
rect 66180 629054 66300 629082
rect 66074 477864 66130 477873
rect 66074 477799 66130 477808
rect 66180 345014 66208 629054
rect 66916 527241 66944 629303
rect 66902 527232 66958 527241
rect 66902 527167 66958 527176
rect 67376 478689 67404 629983
rect 67454 629640 67510 629649
rect 67454 629575 67510 629584
rect 68282 629640 68338 629649
rect 68282 629575 68338 629584
rect 67468 629474 67496 629575
rect 67546 629504 67602 629513
rect 67456 629468 67508 629474
rect 67546 629439 67602 629448
rect 67456 629410 67508 629416
rect 67560 629406 67588 629439
rect 67548 629400 67600 629406
rect 67548 629342 67600 629348
rect 67456 629332 67508 629338
rect 67456 629274 67508 629280
rect 67468 625154 67496 629274
rect 67468 625126 67588 625154
rect 67454 540968 67510 540977
rect 67454 540903 67510 540912
rect 67362 478680 67418 478689
rect 67362 478615 67418 478624
rect 66088 344986 66208 345014
rect 66088 343369 66116 344986
rect 67468 344593 67496 540903
rect 67454 344584 67510 344593
rect 67454 344519 67510 344528
rect 66166 343632 66222 343641
rect 66166 343567 66222 343576
rect 66074 343360 66130 343369
rect 66074 343295 66130 343304
rect 66180 342514 66208 343567
rect 66168 342508 66220 342514
rect 66168 342450 66220 342456
rect 67454 342136 67510 342145
rect 67454 342071 67510 342080
rect 67468 341018 67496 342071
rect 67456 341012 67508 341018
rect 67456 340954 67508 340960
rect 67560 340218 67588 625126
rect 68296 579601 68324 629575
rect 68940 629542 68968 630255
rect 68928 629536 68980 629542
rect 68928 629478 68980 629484
rect 68742 604480 68798 604489
rect 68742 604415 68798 604424
rect 68650 601080 68706 601089
rect 68650 601015 68706 601024
rect 68282 579592 68338 579601
rect 68282 579527 68338 579536
rect 68098 531312 68154 531321
rect 68098 531247 68154 531256
rect 67914 523016 67970 523025
rect 67914 522951 67970 522960
rect 67928 478802 67956 522951
rect 68112 478938 68140 531247
rect 68466 525872 68522 525881
rect 68466 525807 68522 525816
rect 68190 517576 68246 517585
rect 68190 517511 68246 517520
rect 68204 479505 68232 517511
rect 68282 507920 68338 507929
rect 68282 507855 68338 507864
rect 68190 479496 68246 479505
rect 68190 479431 68246 479440
rect 68112 478910 68232 478938
rect 67928 478774 68140 478802
rect 68112 477630 68140 478774
rect 68100 477624 68152 477630
rect 68100 477566 68152 477572
rect 68204 477562 68232 478910
rect 68192 477556 68244 477562
rect 68192 477498 68244 477504
rect 68296 468489 68324 507855
rect 68480 477698 68508 525807
rect 68558 500848 68614 500857
rect 68558 500783 68614 500792
rect 68468 477692 68520 477698
rect 68468 477634 68520 477640
rect 68282 468480 68338 468489
rect 68282 468415 68338 468424
rect 68572 446457 68600 500783
rect 68664 476785 68692 601015
rect 68650 476776 68706 476785
rect 68650 476711 68706 476720
rect 68756 475425 68784 604415
rect 68834 514040 68890 514049
rect 68834 513975 68890 513984
rect 68742 475416 68798 475425
rect 68742 475351 68798 475360
rect 68558 446448 68614 446457
rect 68558 446383 68614 446392
rect 68848 351121 68876 513975
rect 68926 483032 68982 483041
rect 68926 482967 68982 482976
rect 68834 351112 68890 351121
rect 68834 351047 68890 351056
rect 68940 340785 68968 482967
rect 68926 340776 68982 340785
rect 68926 340711 68982 340720
rect 60890 340190 60964 340218
rect 62546 340190 62620 340218
rect 64202 340190 64276 340218
rect 65858 340190 65932 340218
rect 67514 340190 67588 340218
rect 60890 339932 60918 340190
rect 62546 339932 62574 340190
rect 64202 339932 64230 340190
rect 65858 339932 65886 340190
rect 67514 339932 67542 340190
rect 68940 340105 68968 340711
rect 69216 340218 69244 630799
rect 69570 571296 69626 571305
rect 69570 571231 69626 571240
rect 69584 340241 69612 571231
rect 69754 487384 69810 487393
rect 69754 487319 69810 487328
rect 69768 478553 69796 487319
rect 69754 478544 69810 478553
rect 69754 478479 69810 478488
rect 69860 478417 69888 632839
rect 69846 478408 69902 478417
rect 69846 478343 69902 478352
rect 69952 478281 69980 633111
rect 70030 632768 70086 632777
rect 70030 632703 70086 632712
rect 69938 478272 69994 478281
rect 69938 478207 69994 478216
rect 70044 477601 70072 632703
rect 72988 631553 73016 703520
rect 89180 700369 89208 703520
rect 86222 700360 86278 700369
rect 86222 700295 86278 700304
rect 89166 700360 89222 700369
rect 89166 700295 89222 700304
rect 85856 632732 85908 632738
rect 85856 632674 85908 632680
rect 79782 632224 79838 632233
rect 79782 632159 79838 632168
rect 73712 632120 73764 632126
rect 73712 632062 73764 632068
rect 72974 631544 73030 631553
rect 72974 631479 73030 631488
rect 70214 631000 70270 631009
rect 70214 630935 70270 630944
rect 70122 496360 70178 496369
rect 70122 496295 70178 496304
rect 70030 477592 70086 477601
rect 70030 477527 70086 477536
rect 69664 442944 69716 442950
rect 69664 442886 69716 442892
rect 69676 442270 69704 442886
rect 69664 442264 69716 442270
rect 69664 442206 69716 442212
rect 69676 352578 69704 442206
rect 69664 352572 69716 352578
rect 69664 352514 69716 352520
rect 69170 340190 69244 340218
rect 69570 340232 69626 340241
rect 68926 340096 68982 340105
rect 68926 340031 68982 340040
rect 69170 339932 69198 340190
rect 69570 340167 69626 340176
rect 70136 340105 70164 496295
rect 70228 442950 70256 630935
rect 70582 630728 70638 630737
rect 70582 630663 70638 630672
rect 70216 442944 70268 442950
rect 70216 442886 70268 442892
rect 70306 342136 70362 342145
rect 70306 342071 70362 342080
rect 70214 342000 70270 342009
rect 70214 341935 70270 341944
rect 70228 341154 70256 341935
rect 70216 341148 70268 341154
rect 70216 341090 70268 341096
rect 70320 341086 70348 342071
rect 70490 341864 70546 341873
rect 70490 341799 70546 341808
rect 70504 341465 70532 341799
rect 70490 341456 70546 341465
rect 70490 341391 70546 341400
rect 70308 341080 70360 341086
rect 70308 341022 70360 341028
rect 70122 340096 70178 340105
rect 70122 340031 70178 340040
rect 70596 339946 70624 630663
rect 73724 629884 73752 632062
rect 79796 629884 79824 632159
rect 85868 629884 85896 632674
rect 86236 632369 86264 700295
rect 87604 683188 87656 683194
rect 87604 683130 87656 683136
rect 86868 633412 86920 633418
rect 86868 633354 86920 633360
rect 86222 632360 86278 632369
rect 86222 632295 86278 632304
rect 86236 631417 86264 632295
rect 86880 632233 86908 633354
rect 87616 632233 87644 683130
rect 104070 634128 104126 634137
rect 104070 634063 104126 634072
rect 88246 633176 88302 633185
rect 88246 633111 88302 633120
rect 88260 632942 88288 633111
rect 88248 632936 88300 632942
rect 88248 632878 88300 632884
rect 98000 632868 98052 632874
rect 98000 632810 98052 632816
rect 91100 632800 91152 632806
rect 91100 632742 91152 632748
rect 91928 632800 91980 632806
rect 91928 632742 91980 632748
rect 91112 632262 91140 632742
rect 91100 632256 91152 632262
rect 86866 632224 86922 632233
rect 86866 632159 86922 632168
rect 87602 632224 87658 632233
rect 91100 632198 91152 632204
rect 87602 632159 87658 632168
rect 86222 631408 86278 631417
rect 86222 631343 86278 631352
rect 87616 631281 87644 632159
rect 87602 631272 87658 631281
rect 87602 631207 87658 631216
rect 91940 629884 91968 632742
rect 98012 632194 98040 632810
rect 98000 632188 98052 632194
rect 98000 632130 98052 632136
rect 98012 629884 98040 632130
rect 104084 629884 104112 634063
rect 105464 633321 105492 703520
rect 137848 700505 137876 703520
rect 154132 700641 154160 703520
rect 170324 700777 170352 703520
rect 202800 700777 202828 703520
rect 218992 700913 219020 703520
rect 218978 700904 219034 700913
rect 218978 700839 219034 700848
rect 170310 700768 170366 700777
rect 170310 700703 170366 700712
rect 189722 700768 189778 700777
rect 189722 700703 189778 700712
rect 202786 700768 202842 700777
rect 202786 700703 202842 700712
rect 154118 700632 154174 700641
rect 154118 700567 154174 700576
rect 137834 700496 137890 700505
rect 137834 700431 137890 700440
rect 134430 657928 134486 657937
rect 134430 657863 134486 657872
rect 129002 655616 129058 655625
rect 129002 655551 129058 655560
rect 122286 653576 122342 653585
rect 122286 653511 122342 653520
rect 116214 653440 116270 653449
rect 116214 653375 116270 653384
rect 105450 633312 105506 633321
rect 105450 633247 105506 633256
rect 110142 631000 110198 631009
rect 110142 630935 110198 630944
rect 110156 629884 110184 630935
rect 116228 629898 116256 653375
rect 115952 629884 116256 629898
rect 115952 629870 116242 629884
rect 115952 629678 115980 629870
rect 115940 629672 115992 629678
rect 122300 629626 122328 653511
rect 129016 634814 129044 655551
rect 128832 634786 129044 634814
rect 128832 630698 128860 634786
rect 128820 630692 128872 630698
rect 128820 630634 128872 630640
rect 128832 629898 128860 630634
rect 134444 629898 134472 657863
rect 183006 657520 183062 657529
rect 183006 657455 183062 657464
rect 140042 656568 140098 656577
rect 140042 656503 140098 656512
rect 140056 654134 140084 656503
rect 152462 655888 152518 655897
rect 152462 655823 152518 655832
rect 146942 655752 146998 655761
rect 146942 655687 146998 655696
rect 140056 654106 140176 654134
rect 140148 630873 140176 654106
rect 140134 630864 140190 630873
rect 140134 630799 140190 630808
rect 140502 630864 140558 630873
rect 140502 630799 140558 630808
rect 128386 629870 128860 629898
rect 134168 629884 134472 629898
rect 140516 629884 140544 630799
rect 146956 630737 146984 655687
rect 152476 634814 152504 655823
rect 159362 654800 159418 654809
rect 159362 654735 159418 654744
rect 152476 634786 152688 634814
rect 152660 632777 152688 634786
rect 152646 632768 152702 632777
rect 152646 632703 152702 632712
rect 146942 630728 146998 630737
rect 146942 630663 146998 630672
rect 146956 629898 146984 630663
rect 134168 629870 134458 629884
rect 146602 629870 146984 629898
rect 152660 629884 152688 632703
rect 159376 632641 159404 654735
rect 170862 652080 170918 652089
rect 170862 652015 170918 652024
rect 164790 634264 164846 634273
rect 164790 634199 164846 634208
rect 158718 632632 158774 632641
rect 158718 632567 158774 632576
rect 159362 632632 159418 632641
rect 159362 632567 159418 632576
rect 158732 629884 158760 632567
rect 164804 632505 164832 634199
rect 164790 632496 164846 632505
rect 164790 632431 164846 632440
rect 164804 629884 164832 632431
rect 170876 630193 170904 652015
rect 176934 635488 176990 635497
rect 176934 635423 176990 635432
rect 170862 630184 170918 630193
rect 170862 630119 170918 630128
rect 170876 629884 170904 630119
rect 176658 630048 176714 630057
rect 176658 629983 176714 629992
rect 176672 629898 176700 629983
rect 176948 629898 176976 635423
rect 183020 629921 183048 657455
rect 189736 657121 189764 700703
rect 235184 657529 235212 703520
rect 267660 701049 267688 703520
rect 267646 701040 267702 701049
rect 267646 700975 267702 700984
rect 283852 700233 283880 703520
rect 292854 701040 292910 701049
rect 292854 700975 292910 700984
rect 292762 700768 292818 700777
rect 292762 700703 292818 700712
rect 292578 700632 292634 700641
rect 292578 700567 292634 700576
rect 283838 700224 283894 700233
rect 283838 700159 283894 700168
rect 235170 657520 235226 657529
rect 235170 657455 235226 657464
rect 189078 657112 189134 657121
rect 189078 657047 189134 657056
rect 189722 657112 189778 657121
rect 189722 657047 189778 657056
rect 176672 629884 176976 629898
rect 183006 629912 183062 629921
rect 176672 629870 176962 629884
rect 115940 629614 115992 629620
rect 122024 629612 122328 629626
rect 122024 629610 122314 629612
rect 122012 629604 122314 629610
rect 122064 629598 122314 629604
rect 122012 629546 122064 629552
rect 134168 629338 134196 629870
rect 183006 629847 183062 629856
rect 189092 629785 189120 657047
rect 225510 656432 225566 656441
rect 225510 656367 225566 656376
rect 213182 656296 213238 656305
rect 213182 656231 213238 656240
rect 200762 656160 200818 656169
rect 200762 656095 200818 656104
rect 195242 656024 195298 656033
rect 195242 655959 195298 655968
rect 195256 633321 195284 655959
rect 200776 654134 200804 656095
rect 207662 654528 207718 654537
rect 207662 654463 207718 654472
rect 200776 654106 200896 654134
rect 195242 633312 195298 633321
rect 195242 633247 195298 633256
rect 195256 629898 195284 633247
rect 200868 632369 200896 654106
rect 200854 632360 200910 632369
rect 200854 632295 200910 632304
rect 201222 632360 201278 632369
rect 201222 632295 201278 632304
rect 195178 629870 195284 629898
rect 201236 629884 201264 632295
rect 207676 632233 207704 654463
rect 207662 632224 207718 632233
rect 207662 632159 207718 632168
rect 207676 629898 207704 632159
rect 213196 632097 213224 656231
rect 224960 656192 225012 656198
rect 224960 656134 225012 656140
rect 224972 655625 225000 656134
rect 224958 655616 225014 655625
rect 224958 655551 225014 655560
rect 219438 654664 219494 654673
rect 219438 654599 219494 654608
rect 213182 632088 213238 632097
rect 213182 632023 213238 632032
rect 207322 629870 207704 629898
rect 213196 629898 213224 632023
rect 213196 629870 213394 629898
rect 189078 629776 189134 629785
rect 189078 629711 189134 629720
rect 219452 629649 219480 654599
rect 219438 629640 219494 629649
rect 219438 629575 219494 629584
rect 225524 629513 225552 656367
rect 237656 655580 237708 655586
rect 237656 655522 237708 655528
rect 231584 654832 231636 654838
rect 231584 654774 231636 654780
rect 231596 629898 231624 654774
rect 231320 629884 231624 629898
rect 231320 629870 231610 629884
rect 231320 629542 231348 629870
rect 231308 629536 231360 629542
rect 225510 629504 225566 629513
rect 237668 629490 237696 655522
rect 274548 654560 274600 654566
rect 274548 654502 274600 654508
rect 262126 653712 262182 653721
rect 262126 653647 262182 653656
rect 243728 650684 243780 650690
rect 243728 650626 243780 650632
rect 243740 629898 243768 650626
rect 249798 649224 249854 649233
rect 249798 649159 249854 649168
rect 231308 629478 231360 629484
rect 237392 629476 237696 629490
rect 243464 629884 243768 629898
rect 243464 629870 243754 629884
rect 237392 629474 237682 629476
rect 225510 629439 225566 629448
rect 237380 629468 237682 629474
rect 237432 629462 237682 629468
rect 237380 629410 237432 629416
rect 243464 629406 243492 629870
rect 249812 629649 249840 649159
rect 255964 647896 256016 647902
rect 255964 647838 256016 647844
rect 255976 632942 256004 647838
rect 255964 632936 256016 632942
rect 255964 632878 256016 632884
rect 255976 629898 256004 632878
rect 262140 632097 262168 653647
rect 268014 632224 268070 632233
rect 274560 632194 274588 654502
rect 286968 654492 287020 654498
rect 286968 654434 287020 654440
rect 281448 642388 281500 642394
rect 281448 642330 281500 642336
rect 281460 632262 281488 642330
rect 286980 632330 287008 654434
rect 289818 636848 289874 636857
rect 289818 636783 289874 636792
rect 289832 633321 289860 636783
rect 289818 633312 289874 633321
rect 289818 633247 289874 633256
rect 286232 632324 286284 632330
rect 286232 632266 286284 632272
rect 286968 632324 287020 632330
rect 286968 632266 287020 632272
rect 280160 632256 280212 632262
rect 280160 632198 280212 632204
rect 281448 632256 281500 632262
rect 281448 632198 281500 632204
rect 268014 632159 268070 632168
rect 274548 632188 274600 632194
rect 262126 632088 262182 632097
rect 262126 632023 262182 632032
rect 262140 629898 262168 632023
rect 255898 629870 256004 629898
rect 261970 629870 262168 629898
rect 268028 629884 268056 632159
rect 274548 632130 274600 632136
rect 274560 629898 274588 632130
rect 274114 629870 274588 629898
rect 280172 629884 280200 632198
rect 286244 629884 286272 632266
rect 249798 629640 249854 629649
rect 249798 629575 249854 629584
rect 243452 629400 243504 629406
rect 243452 629342 243504 629348
rect 134156 629332 134208 629338
rect 134156 629274 134208 629280
rect 291290 605976 291346 605985
rect 291290 605911 291346 605920
rect 289910 564496 289966 564505
rect 289910 564431 289966 564440
rect 289818 552392 289874 552401
rect 289818 552327 289874 552336
rect 289358 507920 289414 507929
rect 289358 507855 289414 507864
rect 289372 489914 289400 507855
rect 289542 499760 289598 499769
rect 289542 499695 289598 499704
rect 289450 491328 289506 491337
rect 289450 491263 289506 491272
rect 289188 489886 289400 489914
rect 288990 480312 289046 480321
rect 288990 480247 289046 480256
rect 278226 480176 278282 480185
rect 72514 477592 72570 477601
rect 72514 477527 72570 477536
rect 70674 341456 70730 341465
rect 70674 341391 70730 341400
rect 70688 341057 70716 341391
rect 70674 341048 70730 341057
rect 70674 340983 70730 340992
rect 72528 340218 72556 477527
rect 73724 389473 73752 480148
rect 79138 478680 79194 478689
rect 79138 478615 79194 478624
rect 75826 477864 75882 477873
rect 75826 477799 75882 477808
rect 73710 389464 73766 389473
rect 73710 389399 73766 389408
rect 73710 342816 73766 342825
rect 73710 342751 73766 342760
rect 72482 340190 72556 340218
rect 70596 339918 70840 339946
rect 72482 339932 72510 340190
rect 73724 339946 73752 342751
rect 75840 340218 75868 477799
rect 77298 342680 77354 342689
rect 77298 342615 77354 342624
rect 75794 340190 75868 340218
rect 73724 339918 74152 339946
rect 75794 339932 75822 340190
rect 77312 339946 77340 342615
rect 79152 340218 79180 478615
rect 79796 390017 79824 480148
rect 84106 478408 84162 478417
rect 84106 478343 84162 478352
rect 79782 390008 79838 390017
rect 79782 389943 79838 389952
rect 80334 343496 80390 343505
rect 80334 343431 80390 343440
rect 79106 340190 79180 340218
rect 77312 339918 77464 339946
rect 79106 339932 79134 340190
rect 80348 339946 80376 343431
rect 81990 343224 82046 343233
rect 81990 343159 82046 343168
rect 82004 339946 82032 343159
rect 84120 340218 84148 478343
rect 85868 390561 85896 480148
rect 91940 391105 91968 480148
rect 94044 475380 94096 475386
rect 94044 475322 94096 475328
rect 91926 391096 91982 391105
rect 91926 391031 91982 391040
rect 85854 390552 85910 390561
rect 85854 390487 85910 390496
rect 85578 343360 85634 343369
rect 85578 343295 85634 343304
rect 84074 340190 84148 340218
rect 80348 339918 80776 339946
rect 82004 339918 82432 339946
rect 84074 339932 84102 340190
rect 85592 339946 85620 343295
rect 88614 343088 88670 343097
rect 88614 343023 88670 343032
rect 86960 342576 87012 342582
rect 86960 342518 87012 342524
rect 86972 339946 87000 342518
rect 88628 339946 88656 343023
rect 90270 342952 90326 342961
rect 90270 342887 90326 342896
rect 90284 339946 90312 342887
rect 92020 342508 92072 342514
rect 92020 342450 92072 342456
rect 92032 339946 92060 342450
rect 94056 340218 94084 475322
rect 95700 422952 95752 422958
rect 95700 422894 95752 422900
rect 95712 340218 95740 422894
rect 98012 391649 98040 480148
rect 99378 478272 99434 478281
rect 99378 478207 99434 478216
rect 102322 478272 102378 478281
rect 102322 478207 102378 478216
rect 99010 478136 99066 478145
rect 99010 478071 99066 478080
rect 97998 391640 98054 391649
rect 97998 391575 98054 391584
rect 97356 371884 97408 371890
rect 97356 371826 97408 371832
rect 97368 340218 97396 371826
rect 99024 340218 99052 478071
rect 99392 341834 99420 478207
rect 99380 341828 99432 341834
rect 99380 341770 99432 341776
rect 100300 341828 100352 341834
rect 100300 341770 100352 341776
rect 99392 341222 99420 341770
rect 99380 341216 99432 341222
rect 99380 341158 99432 341164
rect 94010 340190 94084 340218
rect 95666 340190 95740 340218
rect 97322 340190 97396 340218
rect 98978 340190 99052 340218
rect 85592 339918 85744 339946
rect 86972 339918 87400 339946
rect 88628 339918 89056 339946
rect 90284 339918 90712 339946
rect 92032 339918 92368 339946
rect 94010 339932 94038 340190
rect 95666 339932 95694 340190
rect 97322 339932 97350 340190
rect 98978 339946 99006 340190
rect 98656 339932 99006 339946
rect 100312 339946 100340 341770
rect 102336 340218 102364 478207
rect 104084 392193 104112 480148
rect 104162 478408 104218 478417
rect 104162 478343 104218 478352
rect 104070 392184 104126 392193
rect 104070 392119 104126 392128
rect 104176 341290 104204 478343
rect 105542 478000 105598 478009
rect 105542 477935 105598 477944
rect 105556 345014 105584 477935
rect 108302 477864 108358 477873
rect 108302 477799 108358 477808
rect 106922 477728 106978 477737
rect 106922 477663 106978 477672
rect 105280 344986 105584 345014
rect 105280 342446 105308 344986
rect 105268 342440 105320 342446
rect 105268 342382 105320 342388
rect 104164 341284 104216 341290
rect 104164 341226 104216 341232
rect 102290 340190 102364 340218
rect 98656 339918 98992 339932
rect 100312 339918 100648 339946
rect 59096 339646 59248 339674
rect 98656 339522 98684 339918
rect 102290 339674 102318 340190
rect 104176 339946 104204 341226
rect 103960 339918 104204 339946
rect 105280 339946 105308 342382
rect 106936 342378 106964 477663
rect 106924 342372 106976 342378
rect 106924 342314 106976 342320
rect 106936 339946 106964 342314
rect 108316 342310 108344 477799
rect 110156 454753 110184 480148
rect 110142 454744 110198 454753
rect 110142 454679 110198 454688
rect 112994 440736 113050 440745
rect 112994 440671 113050 440680
rect 111062 388376 111118 388385
rect 111062 388311 111118 388320
rect 110052 379568 110104 379574
rect 110052 379510 110104 379516
rect 108304 342304 108356 342310
rect 108304 342246 108356 342252
rect 108316 339946 108344 342246
rect 105280 339918 105616 339946
rect 106936 339918 107272 339946
rect 108316 339918 108928 339946
rect 102152 339660 102318 339674
rect 102152 339646 102304 339660
rect 102152 339590 102180 339646
rect 102140 339584 102192 339590
rect 102140 339526 102192 339532
rect 98644 339516 98696 339522
rect 98644 339458 98696 339464
rect 50632 280758 50968 280786
rect 78956 280152 79008 280158
rect 69156 280120 69212 280129
rect 52624 280078 52960 280106
rect 54280 280078 54616 280106
rect 55936 280078 56272 280106
rect 57592 280078 57744 280106
rect 52932 277409 52960 280078
rect 54588 278769 54616 280078
rect 54574 278760 54630 278769
rect 54574 278695 54630 278704
rect 56244 278633 56272 280078
rect 56230 278624 56286 278633
rect 56230 278559 56286 278568
rect 52918 277400 52974 277409
rect 52918 277335 52974 277344
rect 57716 277137 57744 280078
rect 59234 279834 59262 280092
rect 60904 280078 61240 280106
rect 62560 280078 62896 280106
rect 64216 280078 64552 280106
rect 65872 280078 66208 280106
rect 59234 279806 59308 279834
rect 57702 277128 57758 277137
rect 57702 277063 57758 277072
rect 59280 277001 59308 279806
rect 59266 276992 59322 277001
rect 59266 276927 59322 276936
rect 61212 276865 61240 280078
rect 61198 276856 61254 276865
rect 61198 276791 61254 276800
rect 62868 276729 62896 280078
rect 64524 277953 64552 280078
rect 64510 277944 64566 277953
rect 64510 277879 64566 277888
rect 66180 277273 66208 280078
rect 67514 279834 67542 280092
rect 74124 280120 74180 280129
rect 70840 280078 71176 280106
rect 72496 280078 72832 280106
rect 69156 280055 69212 280064
rect 67514 279806 67588 279834
rect 67560 279177 67588 279806
rect 71148 279721 71176 280078
rect 71134 279712 71190 279721
rect 71134 279647 71190 279656
rect 67546 279168 67602 279177
rect 67546 279103 67602 279112
rect 72804 279041 72832 280078
rect 74124 280055 74180 280064
rect 75794 279834 75822 280092
rect 77464 280078 77800 280106
rect 96526 280120 96582 280129
rect 78956 280094 79008 280100
rect 75794 279806 75868 279834
rect 75840 279313 75868 279806
rect 75826 279304 75882 279313
rect 75826 279239 75882 279248
rect 72790 279032 72846 279041
rect 72790 278967 72846 278976
rect 77772 278905 77800 280078
rect 78588 280016 78640 280022
rect 78968 279993 78996 280094
rect 79120 280078 79456 280106
rect 78588 279958 78640 279964
rect 78954 279984 79010 279993
rect 78600 279177 78628 279958
rect 78954 279919 79010 279928
rect 79428 279585 79456 280078
rect 80060 280084 80112 280090
rect 80060 280026 80112 280032
rect 79414 279576 79470 279585
rect 79414 279511 79470 279520
rect 78586 279168 78642 279177
rect 78586 279103 78642 279112
rect 80072 279041 80100 280026
rect 80762 279857 80790 280092
rect 82432 280078 82768 280106
rect 81440 279948 81492 279954
rect 81440 279890 81492 279896
rect 80748 279848 80804 279857
rect 80748 279783 80804 279792
rect 81452 279721 81480 279890
rect 81438 279712 81494 279721
rect 82740 279698 82768 280078
rect 84074 279834 84102 280092
rect 85744 280078 86080 280106
rect 87400 280078 87736 280106
rect 89056 280078 89392 280106
rect 90712 280078 91048 280106
rect 84074 279806 84148 279834
rect 83002 279712 83058 279721
rect 82740 279670 83002 279698
rect 81438 279647 81494 279656
rect 83002 279647 83058 279656
rect 83094 279440 83150 279449
rect 83370 279440 83426 279449
rect 83150 279398 83370 279426
rect 83094 279375 83150 279384
rect 83370 279375 83426 279384
rect 80058 279032 80114 279041
rect 80058 278967 80114 278976
rect 77758 278896 77814 278905
rect 77758 278831 77814 278840
rect 84120 278089 84148 279806
rect 84106 278080 84162 278089
rect 84106 278015 84162 278024
rect 86052 277817 86080 280078
rect 86038 277808 86094 277817
rect 86038 277743 86094 277752
rect 87708 277681 87736 280078
rect 89364 278497 89392 280078
rect 89718 278624 89774 278633
rect 89718 278559 89720 278568
rect 89772 278559 89774 278568
rect 89720 278530 89772 278536
rect 89350 278488 89406 278497
rect 89350 278423 89406 278432
rect 91020 278361 91048 280078
rect 92354 279834 92382 280092
rect 94024 280078 94360 280106
rect 95680 280078 96016 280106
rect 92354 279806 92428 279834
rect 92400 278769 92428 279806
rect 91098 278760 91154 278769
rect 91098 278695 91154 278704
rect 92386 278760 92442 278769
rect 92386 278695 92442 278704
rect 91112 278526 91140 278695
rect 91100 278520 91152 278526
rect 91100 278462 91152 278468
rect 91006 278352 91062 278361
rect 91006 278287 91062 278296
rect 94332 278225 94360 280078
rect 95988 279177 96016 280078
rect 100620 280120 100676 280129
rect 97336 280078 97672 280106
rect 98992 280078 99328 280106
rect 96526 280055 96582 280064
rect 96540 279886 96568 280055
rect 96528 279880 96580 279886
rect 96528 279822 96580 279828
rect 95974 279168 96030 279177
rect 95974 279103 96030 279112
rect 95148 278452 95200 278458
rect 95148 278394 95200 278400
rect 94318 278216 94374 278225
rect 94318 278151 94374 278160
rect 95160 277953 95188 278394
rect 97644 277953 97672 280078
rect 98644 278724 98696 278730
rect 98644 278666 98696 278672
rect 97908 278656 97960 278662
rect 97908 278598 97960 278604
rect 97920 278089 97948 278598
rect 97906 278080 97962 278089
rect 97906 278015 97962 278024
rect 95146 277944 95202 277953
rect 95146 277879 95202 277888
rect 97630 277944 97686 277953
rect 97630 277879 97686 277888
rect 98656 277817 98684 278666
rect 99300 278089 99328 280078
rect 102304 280078 102640 280106
rect 103960 280078 104296 280106
rect 105616 280078 105952 280106
rect 107272 280078 107608 280106
rect 100620 280055 100676 280064
rect 99380 279812 99432 279818
rect 99380 279754 99432 279760
rect 99392 279585 99420 279754
rect 99378 279576 99434 279585
rect 99378 279511 99434 279520
rect 102138 278488 102194 278497
rect 102138 278423 102194 278432
rect 102152 278390 102180 278423
rect 102140 278384 102192 278390
rect 102140 278326 102192 278332
rect 99286 278080 99342 278089
rect 99286 278015 99342 278024
rect 98642 277808 98698 277817
rect 98642 277743 98698 277752
rect 87694 277672 87750 277681
rect 87694 277607 87750 277616
rect 102612 277545 102640 280078
rect 104268 278497 104296 280078
rect 104254 278488 104310 278497
rect 104254 278423 104310 278432
rect 104808 278248 104860 278254
rect 104808 278190 104860 278196
rect 104820 277681 104848 278190
rect 105924 277817 105952 280078
rect 107580 278769 107608 280078
rect 108914 279834 108942 280092
rect 108914 279806 108988 279834
rect 107382 278760 107438 278769
rect 107382 278695 107438 278704
rect 107566 278760 107622 278769
rect 107566 278695 107622 278704
rect 106188 278384 106240 278390
rect 106186 278352 106188 278361
rect 106240 278352 106242 278361
rect 106186 278287 106242 278296
rect 107396 278186 107424 278695
rect 108960 278633 108988 279806
rect 110064 278662 110092 379510
rect 111076 278769 111104 388311
rect 111246 386744 111302 386753
rect 111246 386679 111302 386688
rect 111156 380928 111208 380934
rect 111156 380870 111208 380876
rect 111062 278760 111118 278769
rect 111168 278730 111196 380870
rect 111062 278695 111118 278704
rect 111156 278724 111208 278730
rect 111156 278666 111208 278672
rect 110052 278656 110104 278662
rect 108946 278624 109002 278633
rect 110052 278598 110104 278604
rect 108946 278559 109002 278568
rect 108302 278216 108358 278225
rect 107384 278180 107436 278186
rect 108302 278151 108358 278160
rect 107384 278122 107436 278128
rect 108316 278118 108344 278151
rect 108304 278112 108356 278118
rect 108304 278054 108356 278060
rect 105910 277808 105966 277817
rect 105910 277743 105966 277752
rect 104806 277672 104862 277681
rect 104806 277607 104862 277616
rect 111260 277545 111288 386679
rect 111430 385656 111486 385665
rect 111430 385591 111486 385600
rect 111338 379128 111394 379137
rect 111338 379063 111394 379072
rect 111352 279857 111380 379063
rect 111338 279848 111394 279857
rect 111338 279783 111394 279792
rect 111444 278089 111472 385591
rect 112626 384568 112682 384577
rect 112626 384503 112682 384512
rect 112536 382356 112588 382362
rect 112536 382298 112588 382304
rect 112444 382288 112496 382294
rect 112444 382230 112496 382236
rect 111524 376780 111576 376786
rect 111524 376722 111576 376728
rect 111536 279818 111564 376722
rect 111616 375420 111668 375426
rect 111616 375362 111668 375368
rect 111628 279954 111656 375362
rect 111616 279948 111668 279954
rect 111616 279890 111668 279896
rect 111524 279812 111576 279818
rect 111524 279754 111576 279760
rect 112456 278390 112484 382230
rect 112548 278390 112576 382298
rect 112640 279177 112668 384503
rect 112720 380996 112772 381002
rect 112720 380938 112772 380944
rect 112626 279168 112682 279177
rect 112626 279103 112682 279112
rect 112444 278384 112496 278390
rect 112444 278326 112496 278332
rect 112536 278384 112588 278390
rect 112536 278326 112588 278332
rect 112732 278254 112760 380938
rect 113008 339425 113036 440671
rect 113086 439104 113142 439113
rect 113086 439039 113142 439048
rect 112994 339416 113050 339425
rect 112994 339351 113050 339360
rect 113100 322969 113128 439039
rect 116228 431225 116256 480148
rect 116214 431216 116270 431225
rect 116214 431151 116270 431160
rect 122300 393825 122328 480148
rect 123482 479496 123538 479505
rect 123482 479431 123538 479440
rect 122286 393816 122342 393825
rect 122286 393751 122342 393760
rect 116582 387832 116638 387841
rect 116582 387767 116638 387776
rect 115202 386200 115258 386209
rect 115202 386135 115258 386144
rect 114006 380216 114062 380225
rect 114006 380151 114062 380160
rect 113822 379672 113878 379681
rect 113822 379607 113878 379616
rect 113086 322960 113142 322969
rect 113086 322895 113142 322904
rect 113836 279993 113864 379607
rect 113822 279984 113878 279993
rect 113822 279919 113878 279928
rect 114020 279721 114048 380151
rect 115216 280129 115244 386135
rect 115296 374060 115348 374066
rect 115296 374002 115348 374008
rect 115202 280120 115258 280129
rect 115202 280055 115258 280064
rect 114006 279712 114062 279721
rect 114006 279647 114062 279656
rect 115308 278458 115336 374002
rect 115388 369912 115440 369918
rect 115388 369854 115440 369860
rect 115400 278526 115428 369854
rect 116398 318064 116454 318073
rect 116398 317999 116454 318008
rect 115388 278520 115440 278526
rect 115388 278462 115440 278468
rect 115296 278452 115348 278458
rect 115296 278394 115348 278400
rect 112720 278248 112772 278254
rect 112720 278190 112772 278196
rect 111430 278080 111486 278089
rect 111430 278015 111486 278024
rect 102598 277536 102654 277545
rect 102598 277471 102654 277480
rect 111246 277536 111302 277545
rect 111246 277471 111302 277480
rect 66166 277264 66222 277273
rect 66166 277199 66222 277208
rect 62854 276720 62910 276729
rect 62854 276655 62910 276664
rect 98642 272640 98698 272649
rect 98642 272575 98698 272584
rect 87970 224224 88026 224233
rect 87970 224159 88026 224168
rect 85670 204912 85726 204921
rect 85670 204847 85726 204856
rect 52918 87816 52974 87825
rect 52918 87751 52974 87760
rect 50986 85912 51042 85921
rect 50908 85870 50986 85898
rect 50908 84810 50936 85870
rect 50986 85847 51042 85856
rect 52932 84946 52960 87751
rect 63866 87680 63922 87689
rect 63866 87615 63922 87624
rect 59266 87544 59322 87553
rect 59266 87479 59322 87488
rect 57610 87272 57666 87281
rect 57610 87207 57666 87216
rect 54666 87136 54722 87145
rect 54588 87094 54666 87122
rect 54588 84946 54616 87094
rect 54666 87071 54722 87080
rect 56506 86184 56562 86193
rect 56152 86142 56506 86170
rect 56152 84946 56180 86142
rect 56506 86119 56562 86128
rect 57624 84946 57652 87207
rect 59280 84946 59308 87479
rect 62026 87408 62082 87417
rect 62026 87343 62082 87352
rect 60646 85776 60702 85785
rect 60646 85711 60702 85720
rect 60660 84946 60688 85711
rect 62040 85082 62068 87343
rect 52624 84918 52960 84946
rect 54188 84918 54616 84946
rect 55752 84918 56180 84946
rect 57316 84918 57652 84946
rect 58880 84918 59308 84946
rect 60444 84918 60688 84946
rect 61994 85054 62068 85082
rect 61994 84932 62022 85054
rect 63880 84946 63908 87615
rect 84934 87544 84990 87553
rect 84934 87479 84990 87488
rect 73068 87304 73120 87310
rect 73068 87246 73120 87252
rect 70124 87236 70176 87242
rect 70124 87178 70176 87184
rect 65614 87000 65670 87009
rect 65536 86958 65614 86986
rect 65536 84946 65564 86958
rect 65614 86935 65670 86944
rect 68650 86048 68706 86057
rect 68650 85983 68706 85992
rect 66994 85640 67050 85649
rect 66994 85575 67050 85584
rect 67008 84946 67036 85575
rect 68664 84946 68692 85983
rect 70136 84946 70164 87178
rect 73080 84946 73108 87246
rect 74448 87168 74500 87174
rect 74448 87110 74500 87116
rect 74460 85082 74488 87110
rect 76472 87100 76524 87106
rect 76472 87042 76524 87048
rect 63572 84918 63908 84946
rect 65136 84918 65564 84946
rect 66700 84918 67036 84946
rect 68264 84918 68692 84946
rect 69828 84918 70164 84946
rect 72956 84918 73108 84946
rect 74368 85054 74488 85082
rect 74368 84810 74396 85054
rect 76484 84946 76512 87042
rect 81164 87032 81216 87038
rect 81164 86974 81216 86980
rect 84844 87032 84896 87038
rect 84844 86974 84896 86980
rect 81176 84946 81204 86974
rect 76084 84918 76512 84946
rect 80776 84918 81204 84946
rect 82312 84960 82368 84969
rect 82312 84895 82368 84904
rect 77620 84824 77676 84833
rect 50908 84782 51060 84810
rect 74368 84782 74520 84810
rect 77620 84759 77676 84768
rect 71364 84688 71420 84697
rect 71364 84623 71420 84632
rect 79184 84552 79240 84561
rect 83904 84510 84332 84538
rect 79184 84487 79240 84496
rect 84304 83473 84332 84510
rect 84290 83464 84346 83473
rect 84290 83399 84346 83408
rect 84856 79354 84884 86974
rect 84948 80753 84976 87479
rect 85028 87236 85080 87242
rect 85028 87178 85080 87184
rect 85040 83502 85068 87178
rect 85028 83496 85080 83502
rect 85028 83438 85080 83444
rect 84934 80744 84990 80753
rect 84934 80679 84990 80688
rect 84844 79348 84896 79354
rect 84844 79290 84896 79296
rect 49330 78976 49386 78985
rect 49330 78911 49386 78920
rect 49238 69456 49294 69465
rect 49238 69391 49294 69400
rect 49054 68096 49110 68105
rect 49054 68031 49110 68040
rect 48226 51504 48282 51513
rect 48226 51439 48282 51448
rect 48134 49056 48190 49065
rect 48134 48991 48190 49000
rect 49068 48929 49096 68031
rect 49146 54496 49202 54505
rect 49146 54431 49202 54440
rect 49054 48920 49110 48929
rect 49054 48855 49110 48864
rect 48042 42256 48098 42265
rect 48042 42191 48098 42200
rect 49160 30977 49188 54431
rect 49252 39273 49280 69391
rect 49344 44849 49372 78911
rect 49606 77616 49662 77625
rect 49606 77551 49662 77560
rect 49514 74896 49570 74905
rect 49514 74831 49570 74840
rect 49422 72176 49478 72185
rect 49422 72111 49478 72120
rect 49330 44840 49386 44849
rect 49330 44775 49386 44784
rect 49238 39264 49294 39273
rect 49238 39199 49294 39208
rect 49436 37913 49464 72111
rect 49422 37904 49478 37913
rect 49422 37839 49478 37848
rect 49528 35193 49556 74831
rect 49514 35184 49570 35193
rect 49514 35119 49570 35128
rect 49620 32473 49648 77551
rect 50250 75984 50306 75993
rect 50250 75919 50306 75928
rect 50158 70408 50214 70417
rect 50158 70343 50214 70352
rect 50066 52592 50122 52601
rect 50066 52527 50122 52536
rect 50080 43625 50108 52527
rect 50066 43616 50122 43625
rect 50066 43551 50122 43560
rect 49606 32464 49662 32473
rect 49606 32399 49662 32408
rect 49146 30968 49202 30977
rect 49146 30903 49202 30912
rect 47950 22672 48006 22681
rect 47950 22607 48006 22616
rect 47582 19952 47638 19961
rect 47582 19887 47638 19896
rect 47490 18592 47546 18601
rect 47490 18527 47546 18536
rect 50172 17241 50200 70343
rect 50264 33833 50292 75919
rect 50434 73264 50490 73273
rect 50434 73199 50490 73208
rect 50342 66328 50398 66337
rect 50342 66263 50398 66272
rect 50250 33824 50306 33833
rect 50250 33759 50306 33768
rect 50356 25537 50384 66263
rect 50448 36553 50476 73199
rect 50618 65104 50674 65113
rect 50618 65039 50674 65048
rect 50526 55584 50582 55593
rect 50526 55519 50582 55528
rect 50434 36544 50490 36553
rect 50434 36479 50490 36488
rect 50540 29617 50568 55519
rect 50632 46345 50660 65039
rect 84658 53272 84714 53281
rect 84658 53207 84714 53216
rect 83278 50552 83334 50561
rect 83278 50487 83334 50496
rect 50876 50102 51028 50130
rect 52256 50102 52408 50130
rect 53636 50102 53788 50130
rect 51000 47841 51028 50102
rect 50986 47832 51042 47841
rect 50986 47767 51042 47776
rect 52380 47705 52408 50102
rect 52366 47696 52422 47705
rect 52366 47631 52422 47640
rect 53760 47569 53788 50102
rect 55002 49858 55030 50116
rect 56396 50102 56548 50130
rect 57776 50102 57928 50130
rect 55002 49830 55076 49858
rect 53746 47560 53802 47569
rect 53746 47495 53802 47504
rect 50618 46336 50674 46345
rect 50618 46271 50674 46280
rect 51354 38040 51410 38049
rect 51354 37975 51410 37984
rect 50526 29608 50582 29617
rect 50526 29543 50582 29552
rect 50342 25528 50398 25537
rect 50342 25463 50398 25472
rect 50158 17232 50214 17241
rect 50158 17167 50214 17176
rect 48962 7848 49018 7857
rect 48962 7783 49018 7792
rect 47858 6352 47914 6361
rect 47858 6287 47914 6296
rect 47872 480 47900 6287
rect 48976 480 49004 7783
rect 50158 3496 50214 3505
rect 50158 3431 50214 3440
rect 50172 480 50200 3431
rect 51368 480 51396 37975
rect 51722 36680 51778 36689
rect 51722 36615 51778 36624
rect 51736 3505 51764 36615
rect 52550 27160 52606 27169
rect 52550 27095 52606 27104
rect 51722 3496 51778 3505
rect 51722 3431 51778 3440
rect 52564 480 52592 27095
rect 53746 27024 53802 27033
rect 53746 26959 53802 26968
rect 53760 480 53788 26959
rect 54942 6488 54998 6497
rect 54942 6423 54998 6432
rect 54956 480 54984 6423
rect 55048 4865 55076 49830
rect 56520 46209 56548 50102
rect 57900 47818 57928 50102
rect 59142 49858 59170 50116
rect 60522 49858 60550 50116
rect 61902 49858 61930 50116
rect 63282 49858 63310 50116
rect 64662 49858 64690 50116
rect 66042 49858 66070 50116
rect 67422 49858 67450 50116
rect 68802 49858 68830 50116
rect 70182 49858 70210 50116
rect 71562 49858 71590 50116
rect 72942 49858 72970 50116
rect 74336 50102 74488 50130
rect 75716 50102 75868 50130
rect 59142 49830 59216 49858
rect 60522 49830 60596 49858
rect 61902 49830 61976 49858
rect 63282 49830 63356 49858
rect 64662 49830 64736 49858
rect 66042 49830 66116 49858
rect 67422 49830 67496 49858
rect 68802 49830 68876 49858
rect 70182 49830 70256 49858
rect 71562 49830 71636 49858
rect 72942 49830 73016 49858
rect 57900 47790 58664 47818
rect 56506 46200 56562 46209
rect 56506 46135 56562 46144
rect 56046 29880 56102 29889
rect 56046 29815 56102 29824
rect 55034 4856 55090 4865
rect 55034 4791 55090 4800
rect 56060 480 56088 29815
rect 58636 8945 58664 47790
rect 59188 10305 59216 49830
rect 59634 28520 59690 28529
rect 59634 28455 59690 28464
rect 59174 10296 59230 10305
rect 59174 10231 59230 10240
rect 58622 8936 58678 8945
rect 58622 8871 58678 8880
rect 58438 6624 58494 6633
rect 58438 6559 58494 6568
rect 57242 3496 57298 3505
rect 57242 3431 57298 3440
rect 57256 480 57284 3431
rect 58452 480 58480 6559
rect 59648 480 59676 28455
rect 60568 11665 60596 49830
rect 61948 13025 61976 49830
rect 63222 31104 63278 31113
rect 63222 31039 63278 31048
rect 61934 13016 61990 13025
rect 61934 12951 61990 12960
rect 60554 11656 60610 11665
rect 60554 11591 60610 11600
rect 62026 6760 62082 6769
rect 62026 6695 62082 6704
rect 60830 3360 60886 3369
rect 60830 3295 60886 3304
rect 60844 480 60872 3295
rect 62040 480 62068 6695
rect 63236 480 63264 31039
rect 63328 14521 63356 49830
rect 64708 43489 64736 49830
rect 64694 43480 64750 43489
rect 64694 43415 64750 43424
rect 65522 24304 65578 24313
rect 65522 24239 65578 24248
rect 64326 18728 64382 18737
rect 64326 18663 64382 18672
rect 63314 14512 63370 14521
rect 63314 14447 63370 14456
rect 64340 480 64368 18663
rect 65536 480 65564 24239
rect 66088 15881 66116 49830
rect 67468 42129 67496 49830
rect 67454 42120 67510 42129
rect 67454 42055 67510 42064
rect 68848 40633 68876 49830
rect 68834 40624 68890 40633
rect 68834 40559 68890 40568
rect 66718 32736 66774 32745
rect 66718 32671 66774 32680
rect 66074 15872 66130 15881
rect 66074 15807 66130 15816
rect 66732 480 66760 32671
rect 70228 21457 70256 49830
rect 70306 34096 70362 34105
rect 70306 34031 70362 34040
rect 70214 21448 70270 21457
rect 70214 21383 70270 21392
rect 69110 20088 69166 20097
rect 69110 20023 69166 20032
rect 67914 3768 67970 3777
rect 67914 3703 67970 3712
rect 67928 480 67956 3703
rect 69124 480 69152 20023
rect 70320 480 70348 34031
rect 71502 32600 71558 32609
rect 71502 32535 71558 32544
rect 71516 480 71544 32535
rect 71608 10441 71636 49830
rect 72988 21321 73016 49830
rect 74460 47025 74488 50102
rect 75840 47818 75868 50102
rect 77082 49858 77110 50116
rect 78476 50102 78628 50130
rect 77082 49830 77156 49858
rect 75840 47790 76604 47818
rect 74446 47016 74502 47025
rect 74446 46951 74502 46960
rect 75182 47016 75238 47025
rect 75182 46951 75238 46960
rect 73802 35320 73858 35329
rect 73802 35255 73858 35264
rect 72974 21312 73030 21321
rect 72974 21247 73030 21256
rect 71594 10432 71650 10441
rect 71594 10367 71650 10376
rect 72606 6896 72662 6905
rect 72606 6831 72662 6840
rect 72620 480 72648 6831
rect 73816 480 73844 35255
rect 74998 28384 75054 28393
rect 74998 28319 75054 28328
rect 75012 480 75040 28319
rect 75196 11801 75224 46951
rect 76576 13161 76604 47790
rect 77128 14657 77156 49830
rect 78600 47818 78628 50102
rect 79842 49858 79870 50116
rect 81222 49858 81250 50116
rect 82616 50102 82768 50130
rect 79842 49830 79916 49858
rect 81222 49830 81296 49858
rect 78600 47790 79364 47818
rect 77390 36816 77446 36825
rect 77390 36751 77446 36760
rect 77114 14648 77170 14657
rect 77114 14583 77170 14592
rect 76562 13152 76618 13161
rect 76562 13087 76618 13096
rect 75182 11792 75238 11801
rect 75182 11727 75238 11736
rect 76194 6080 76250 6089
rect 76194 6015 76250 6024
rect 76208 480 76236 6015
rect 77404 480 77432 36751
rect 79336 16017 79364 47790
rect 79690 25664 79746 25673
rect 79690 25599 79746 25608
rect 79322 16008 79378 16017
rect 79322 15943 79378 15952
rect 78586 7712 78642 7721
rect 78586 7647 78642 7656
rect 78600 480 78628 7647
rect 79704 480 79732 25599
rect 79888 17377 79916 49830
rect 81268 40769 81296 49830
rect 82740 47977 82768 50102
rect 82726 47968 82782 47977
rect 82726 47903 82782 47912
rect 81254 40760 81310 40769
rect 81254 40695 81310 40704
rect 80886 33960 80942 33969
rect 80886 33895 80942 33904
rect 79874 17368 79930 17377
rect 79874 17303 79930 17312
rect 80900 480 80928 33895
rect 82082 29744 82138 29753
rect 82082 29679 82138 29688
rect 82096 480 82124 29679
rect 83292 480 83320 50487
rect 83982 49858 84010 50116
rect 83982 49830 84056 49858
rect 83462 47968 83518 47977
rect 83462 47903 83518 47912
rect 83476 22817 83504 47903
rect 84028 39409 84056 49830
rect 84014 39400 84070 39409
rect 84014 39335 84070 39344
rect 83462 22808 83518 22817
rect 83462 22743 83518 22752
rect 84672 6914 84700 53207
rect 84488 6886 84700 6914
rect 84488 480 84516 6886
rect 85684 480 85712 204847
rect 86866 91760 86922 91769
rect 86866 91695 86922 91704
rect 86222 87816 86278 87825
rect 86222 87751 86278 87760
rect 86236 51785 86264 87751
rect 86406 87272 86462 87281
rect 86406 87207 86462 87216
rect 86420 53145 86448 87207
rect 86406 53136 86462 53145
rect 86406 53071 86462 53080
rect 86222 51776 86278 51785
rect 86222 51711 86278 51720
rect 86880 480 86908 91695
rect 87602 90400 87658 90409
rect 87602 90335 87658 90344
rect 87616 52601 87644 90335
rect 87878 87680 87934 87689
rect 87878 87615 87934 87624
rect 87694 87136 87750 87145
rect 87694 87071 87750 87080
rect 86958 52592 87014 52601
rect 86958 52527 87014 52536
rect 87602 52592 87658 52601
rect 87602 52527 87658 52536
rect 86972 40905 87000 52527
rect 87708 50289 87736 87071
rect 87892 54641 87920 87615
rect 87878 54632 87934 54641
rect 87878 54567 87934 54576
rect 87694 50280 87750 50289
rect 87694 50215 87750 50224
rect 86958 40896 87014 40905
rect 86958 40831 87014 40840
rect 87984 480 88012 224159
rect 96250 221504 96306 221513
rect 96250 221439 96306 221448
rect 92754 220144 92810 220153
rect 92754 220079 92810 220088
rect 91742 214568 91798 214577
rect 91742 214503 91798 214512
rect 90362 213208 90418 213217
rect 90362 213143 90418 213152
rect 89166 89040 89222 89049
rect 89166 88975 89222 88984
rect 89180 480 89208 88975
rect 90376 480 90404 213143
rect 91558 97200 91614 97209
rect 91558 97135 91614 97144
rect 90638 87408 90694 87417
rect 90638 87343 90694 87352
rect 90454 87000 90510 87009
rect 90454 86935 90510 86944
rect 90468 9081 90496 86935
rect 90652 69601 90680 87343
rect 90638 69592 90694 69601
rect 90638 69527 90694 69536
rect 90454 9072 90510 9081
rect 90454 9007 90510 9016
rect 91572 480 91600 97135
rect 91756 3505 91784 214503
rect 91742 3496 91798 3505
rect 91742 3431 91798 3440
rect 92768 480 92796 220079
rect 93950 211848 94006 211857
rect 93950 211783 94006 211792
rect 93964 480 93992 211783
rect 95146 98696 95202 98705
rect 95146 98631 95202 98640
rect 95160 480 95188 98631
rect 96264 480 96292 221439
rect 97446 210352 97502 210361
rect 97446 210287 97502 210296
rect 97460 480 97488 210287
rect 98656 480 98684 272575
rect 105726 243536 105782 243545
rect 105726 243471 105782 243480
rect 101402 239592 101458 239601
rect 101402 239527 101458 239536
rect 99838 229800 99894 229809
rect 99838 229735 99894 229744
rect 98736 87168 98788 87174
rect 98736 87110 98788 87116
rect 98748 51746 98776 87110
rect 98736 51740 98788 51746
rect 98736 51682 98788 51688
rect 99852 480 99880 229735
rect 101034 177304 101090 177313
rect 101034 177239 101090 177248
rect 101048 480 101076 177239
rect 101416 3777 101444 239527
rect 103334 226944 103390 226953
rect 103334 226879 103390 226888
rect 102230 100056 102286 100065
rect 102230 99991 102286 100000
rect 101402 3768 101458 3777
rect 101402 3703 101458 3712
rect 102244 480 102272 99991
rect 103348 480 103376 226879
rect 104530 208992 104586 209001
rect 104530 208927 104586 208936
rect 104544 480 104572 208927
rect 105740 480 105768 243471
rect 114006 236736 114062 236745
rect 114006 236671 114062 236680
rect 106922 234016 106978 234025
rect 106922 233951 106978 233960
rect 106936 480 106964 233951
rect 110510 222864 110566 222873
rect 110510 222799 110566 222808
rect 108118 178664 108174 178673
rect 108118 178599 108174 178608
rect 108132 480 108160 178599
rect 109314 5128 109370 5137
rect 109314 5063 109370 5072
rect 109328 480 109356 5063
rect 110524 480 110552 222799
rect 112810 101416 112866 101425
rect 112810 101351 112866 101360
rect 111614 93120 111670 93129
rect 111614 93055 111670 93064
rect 111628 480 111656 93055
rect 112824 480 112852 101351
rect 114020 480 114048 236671
rect 115202 207632 115258 207641
rect 115202 207567 115258 207576
rect 115216 480 115244 207567
rect 116412 480 116440 317999
rect 116596 277817 116624 387767
rect 119434 387288 119490 387297
rect 119434 387223 119490 387232
rect 117962 385112 118018 385121
rect 117962 385047 118018 385056
rect 117976 277953 118004 385047
rect 119342 331256 119398 331265
rect 119342 331191 119398 331200
rect 117962 277944 118018 277953
rect 117962 277879 118018 277888
rect 116582 277808 116638 277817
rect 116582 277743 116638 277752
rect 118790 3904 118846 3913
rect 118790 3839 118846 3848
rect 117594 3496 117650 3505
rect 117594 3431 117650 3440
rect 117608 480 117636 3431
rect 118804 480 118832 3839
rect 119356 3641 119384 331191
rect 119448 278497 119476 387223
rect 120722 378584 120778 378593
rect 120722 378519 120778 378528
rect 120736 279313 120764 378519
rect 122196 374128 122248 374134
rect 122196 374070 122248 374076
rect 122102 373688 122158 373697
rect 122102 373623 122158 373632
rect 120722 279304 120778 279313
rect 120722 279239 120778 279248
rect 119434 278488 119490 278497
rect 119434 278423 119490 278432
rect 122116 276729 122144 373623
rect 122208 280022 122236 374070
rect 123496 285025 123524 479431
rect 126244 477692 126296 477698
rect 126244 477634 126296 477640
rect 123576 376848 123628 376854
rect 123576 376790 123628 376796
rect 123482 285016 123538 285025
rect 123482 284951 123538 284960
rect 122196 280016 122248 280022
rect 122196 279958 122248 279964
rect 123588 279886 123616 376790
rect 123666 373144 123722 373153
rect 123666 373079 123722 373088
rect 123576 279880 123628 279886
rect 123576 279822 123628 279828
rect 123680 276865 123708 373079
rect 126256 287026 126284 477634
rect 128372 394369 128400 480148
rect 134444 394913 134472 480148
rect 138664 477624 138716 477630
rect 138664 477566 138716 477572
rect 134430 394904 134486 394913
rect 134430 394839 134486 394848
rect 128358 394360 128414 394369
rect 128358 394295 128414 394304
rect 126334 388920 126390 388929
rect 126334 388855 126390 388864
rect 126244 287020 126296 287026
rect 126244 286962 126296 286968
rect 126348 278633 126376 388855
rect 127624 376916 127676 376922
rect 127624 376858 127676 376864
rect 126428 375488 126480 375494
rect 126428 375430 126480 375436
rect 126440 280158 126468 375430
rect 126428 280152 126480 280158
rect 126428 280094 126480 280100
rect 127636 280090 127664 376858
rect 127714 372600 127770 372609
rect 127714 372535 127770 372544
rect 127624 280084 127676 280090
rect 127624 280026 127676 280032
rect 126334 278624 126390 278633
rect 126334 278559 126390 278568
rect 127728 277001 127756 372535
rect 130382 372056 130438 372065
rect 130382 371991 130438 372000
rect 130396 277137 130424 371991
rect 137284 371272 137336 371278
rect 137284 371214 137336 371220
rect 134522 370424 134578 370433
rect 134522 370359 134578 370368
rect 134536 277409 134564 370359
rect 137296 278594 137324 371214
rect 138676 285666 138704 477566
rect 140516 395457 140544 480148
rect 142896 477556 142948 477562
rect 142896 477498 142948 477504
rect 140502 395448 140558 395457
rect 140502 395383 140558 395392
rect 140042 374776 140098 374785
rect 140042 374711 140098 374720
rect 138664 285660 138716 285666
rect 138664 285602 138716 285608
rect 137284 278588 137336 278594
rect 137284 278530 137336 278536
rect 134522 277400 134578 277409
rect 134522 277335 134578 277344
rect 140056 277273 140084 374711
rect 142802 339416 142858 339425
rect 142802 339351 142858 339360
rect 140042 277264 140098 277273
rect 140042 277199 140098 277208
rect 130382 277128 130438 277137
rect 130382 277063 130438 277072
rect 127714 276992 127770 277001
rect 127714 276927 127770 276936
rect 123666 276856 123722 276865
rect 123666 276791 123722 276800
rect 122102 276720 122158 276729
rect 122102 276655 122158 276664
rect 123482 265568 123538 265577
rect 123482 265503 123538 265512
rect 121460 238672 121512 238678
rect 121460 238614 121512 238620
rect 121472 237425 121500 238614
rect 122286 237824 122342 237833
rect 122286 237759 122342 237768
rect 121458 237416 121514 237425
rect 121458 237351 121514 237360
rect 121090 232520 121146 232529
rect 121090 232455 121146 232464
rect 119894 3768 119950 3777
rect 119894 3703 119950 3712
rect 119342 3632 119398 3641
rect 119342 3567 119398 3576
rect 119908 480 119936 3703
rect 121104 480 121132 232455
rect 122300 480 122328 237759
rect 123496 480 123524 265503
rect 141238 235512 141294 235521
rect 141238 235447 141294 235456
rect 126978 232656 127034 232665
rect 126978 232591 127034 232600
rect 126242 206272 126298 206281
rect 126242 206207 126298 206216
rect 126256 3913 126284 206207
rect 126242 3904 126298 3913
rect 126242 3839 126298 3848
rect 124678 3632 124734 3641
rect 124678 3567 124734 3576
rect 124692 480 124720 3567
rect 126992 480 127020 232591
rect 130566 225720 130622 225729
rect 130566 225655 130622 225664
rect 130580 480 130608 225655
rect 134154 220280 134210 220289
rect 134154 220215 134210 220224
rect 134168 480 134196 220215
rect 137650 200696 137706 200705
rect 137650 200631 137706 200640
rect 137664 480 137692 200631
rect 141252 480 141280 235447
rect 142816 34105 142844 339351
rect 142908 288386 142936 477498
rect 146588 396001 146616 480148
rect 151174 474056 151230 474065
rect 151174 473991 151230 474000
rect 146574 395992 146630 396001
rect 146574 395927 146630 395936
rect 146942 345400 146998 345409
rect 146942 345335 146998 345344
rect 142896 288380 142948 288386
rect 142896 288322 142948 288328
rect 144734 197976 144790 197985
rect 144734 197911 144790 197920
rect 142802 34096 142858 34105
rect 142802 34031 142858 34040
rect 144748 480 144776 197911
rect 146956 5137 146984 345335
rect 151082 336696 151138 336705
rect 151082 336631 151138 336640
rect 148322 239320 148378 239329
rect 148322 239255 148378 239264
rect 146942 5128 146998 5137
rect 146942 5063 146998 5072
rect 148336 480 148364 239255
rect 151096 27169 151124 336631
rect 151188 301889 151216 473991
rect 152660 396545 152688 480148
rect 155222 468480 155278 468489
rect 155222 468415 155278 468424
rect 152646 396536 152702 396545
rect 152646 396471 152702 396480
rect 151174 301880 151230 301889
rect 151174 301815 151230 301824
rect 155236 275777 155264 468415
rect 158732 397089 158760 480148
rect 164804 464409 164832 480148
rect 164790 464400 164846 464409
rect 164790 464335 164846 464344
rect 170876 398177 170904 480148
rect 176948 398721 176976 480148
rect 183020 399265 183048 480148
rect 189092 474065 189120 480148
rect 189078 474056 189134 474065
rect 189078 473991 189134 474000
rect 195164 400353 195192 480148
rect 199474 446448 199530 446457
rect 199474 446383 199530 446392
rect 198832 412684 198884 412690
rect 198832 412626 198884 412632
rect 198844 408542 198872 412626
rect 198004 408536 198056 408542
rect 198004 408478 198056 408484
rect 198832 408536 198884 408542
rect 198832 408478 198884 408484
rect 195150 400344 195206 400353
rect 195150 400279 195206 400288
rect 198016 400246 198044 408478
rect 198004 400240 198056 400246
rect 198004 400182 198056 400188
rect 193864 400172 193916 400178
rect 193864 400114 193916 400120
rect 183006 399256 183062 399265
rect 183006 399191 183062 399200
rect 176934 398712 176990 398721
rect 176934 398647 176990 398656
rect 170862 398168 170918 398177
rect 170862 398103 170918 398112
rect 158718 397080 158774 397089
rect 158718 397015 158774 397024
rect 193876 386374 193904 400114
rect 191840 386368 191892 386374
rect 191840 386310 191892 386316
rect 193864 386368 193916 386374
rect 193864 386310 193916 386316
rect 191852 379522 191880 386310
rect 192484 383716 192536 383722
rect 192484 383658 192536 383664
rect 191760 379506 191880 379522
rect 186964 379500 187016 379506
rect 186964 379442 187016 379448
rect 191748 379500 191880 379506
rect 191800 379494 191880 379500
rect 191748 379442 191800 379448
rect 186976 358766 187004 379442
rect 185584 358760 185636 358766
rect 185584 358702 185636 358708
rect 186964 358760 187016 358766
rect 186964 358702 187016 358708
rect 159362 349752 159418 349761
rect 159362 349687 159418 349696
rect 155222 275768 155278 275777
rect 155222 275703 155278 275712
rect 158902 239048 158958 239057
rect 158902 238983 158958 238992
rect 155406 231160 155462 231169
rect 155406 231095 155462 231104
rect 151818 196616 151874 196625
rect 151818 196551 151874 196560
rect 151082 27160 151138 27169
rect 151082 27095 151138 27104
rect 151832 480 151860 196551
rect 155420 480 155448 231095
rect 158916 480 158944 238983
rect 159376 18873 159404 349687
rect 185596 347750 185624 358702
rect 182180 347744 182232 347750
rect 182180 347686 182232 347692
rect 185584 347744 185636 347750
rect 185584 347686 185636 347692
rect 163502 347032 163558 347041
rect 163502 346967 163558 346976
rect 162490 236872 162546 236881
rect 162490 236807 162546 236816
rect 159362 18864 159418 18873
rect 159362 18799 159418 18808
rect 162504 480 162532 236807
rect 163516 3777 163544 346967
rect 182192 344350 182220 347686
rect 182180 344344 182232 344350
rect 182180 344286 182232 344292
rect 174542 343224 174598 343233
rect 174542 343159 174598 343168
rect 173162 239184 173218 239193
rect 173162 239119 173218 239128
rect 166078 228440 166134 228449
rect 166078 228375 166134 228384
rect 163502 3768 163558 3777
rect 163502 3703 163558 3712
rect 166092 480 166120 228375
rect 169574 3768 169630 3777
rect 169574 3703 169630 3712
rect 169588 480 169616 3703
rect 173176 480 173204 239119
rect 174556 98705 174584 343159
rect 175922 338872 175978 338881
rect 175922 338807 175978 338816
rect 174542 98696 174598 98705
rect 174542 98631 174598 98640
rect 175936 32745 175964 338807
rect 178682 337784 178738 337793
rect 178682 337719 178738 337728
rect 176658 239456 176714 239465
rect 176658 239391 176714 239400
rect 175922 32736 175978 32745
rect 175922 32671 175978 32680
rect 176672 480 176700 239391
rect 178696 28529 178724 337719
rect 188342 337240 188398 337249
rect 188342 337175 188398 337184
rect 184202 335608 184258 335617
rect 184202 335543 184258 335552
rect 179420 239420 179472 239426
rect 179420 239362 179472 239368
rect 179432 238785 179460 239362
rect 180246 238912 180302 238921
rect 180246 238847 180302 238856
rect 179418 238776 179474 238785
rect 179418 238711 179474 238720
rect 178682 28520 178738 28529
rect 178682 28455 178738 28464
rect 180260 480 180288 238847
rect 183742 235648 183798 235657
rect 183742 235583 183798 235592
rect 183756 480 183784 235583
rect 184216 106865 184244 335543
rect 186962 333976 187018 333985
rect 186962 333911 187018 333920
rect 186976 244905 187004 333911
rect 186962 244896 187018 244905
rect 186962 244831 187018 244840
rect 186320 240100 186372 240106
rect 186320 240042 186372 240048
rect 186332 239601 186360 240042
rect 186318 239592 186374 239601
rect 186318 239527 186374 239536
rect 187330 238776 187386 238785
rect 187330 238711 187386 238720
rect 184202 106856 184258 106865
rect 184202 106791 184258 106800
rect 187344 480 187372 238711
rect 188356 29889 188384 337175
rect 191102 335064 191158 335073
rect 191102 334999 191158 335008
rect 190826 229936 190882 229945
rect 190826 229871 190882 229880
rect 188342 29880 188398 29889
rect 188342 29815 188398 29824
rect 190840 480 190868 229871
rect 191116 105505 191144 334999
rect 192496 278118 192524 383658
rect 199382 345944 199438 345953
rect 199382 345879 199438 345888
rect 195242 340504 195298 340513
rect 195242 340439 195298 340448
rect 192484 278112 192536 278118
rect 192484 278054 192536 278060
rect 194414 231296 194470 231305
rect 194414 231231 194470 231240
rect 191102 105496 191158 105505
rect 191102 105431 191158 105440
rect 194428 480 194456 231231
rect 195256 36825 195284 340439
rect 198002 334520 198058 334529
rect 198002 334455 198058 334464
rect 197910 234152 197966 234161
rect 197910 234087 197966 234096
rect 195242 36816 195298 36825
rect 195242 36751 195298 36760
rect 197924 480 197952 234087
rect 198016 104145 198044 334455
rect 198002 104136 198058 104145
rect 198002 104071 198058 104080
rect 199396 101425 199424 345879
rect 199488 275233 199516 446383
rect 201236 400897 201264 480148
rect 207020 422340 207072 422346
rect 207020 422282 207072 422288
rect 207032 418198 207060 422282
rect 207020 418192 207072 418198
rect 207020 418134 207072 418140
rect 202880 418124 202932 418130
rect 202880 418066 202932 418072
rect 202892 415426 202920 418066
rect 202800 415398 202920 415426
rect 202800 412690 202828 415398
rect 202788 412684 202840 412690
rect 202788 412626 202840 412632
rect 207308 401441 207336 480148
rect 211802 431216 211858 431225
rect 211802 431151 211858 431160
rect 211620 430636 211672 430642
rect 211620 430578 211672 430584
rect 211632 422346 211660 430578
rect 211620 422340 211672 422346
rect 211620 422282 211672 422288
rect 207294 401432 207350 401441
rect 207294 401367 207350 401376
rect 201222 400888 201278 400897
rect 201222 400823 201278 400832
rect 211816 393281 211844 431151
rect 213380 401985 213408 480148
rect 214654 475416 214710 475425
rect 214654 475351 214710 475360
rect 213552 434716 213604 434722
rect 213552 434658 213604 434664
rect 213564 430642 213592 434658
rect 213552 430636 213604 430642
rect 213552 430578 213604 430584
rect 213366 401976 213422 401985
rect 213366 401911 213422 401920
rect 211802 393272 211858 393281
rect 211802 393207 211858 393216
rect 210422 348664 210478 348673
rect 210422 348599 210478 348608
rect 202142 344856 202198 344865
rect 202142 344791 202198 344800
rect 199474 275224 199530 275233
rect 199474 275159 199530 275168
rect 202156 243545 202184 344791
rect 203522 338328 203578 338337
rect 203522 338263 203578 338272
rect 202142 243536 202198 243545
rect 202142 243471 202198 243480
rect 201498 237008 201554 237017
rect 201498 236943 201554 236952
rect 199382 101416 199438 101425
rect 199382 101351 199438 101360
rect 201512 480 201540 236943
rect 203536 31113 203564 338263
rect 206282 336152 206338 336161
rect 206282 336087 206338 336096
rect 205086 223000 205142 223009
rect 205086 222935 205142 222944
rect 203522 31104 203578 31113
rect 203522 31039 203578 31048
rect 205100 480 205128 222935
rect 206296 7857 206324 336087
rect 209042 332888 209098 332897
rect 209042 332823 209098 332832
rect 208582 232792 208638 232801
rect 208582 232727 208638 232736
rect 206282 7848 206338 7857
rect 206282 7783 206338 7792
rect 208596 480 208624 232727
rect 209056 102785 209084 332823
rect 209042 102776 209098 102785
rect 209042 102711 209098 102720
rect 210436 94489 210464 348599
rect 211802 342680 211858 342689
rect 211802 342615 211858 342624
rect 211816 97209 211844 342615
rect 213184 341216 213236 341222
rect 213184 341158 213236 341164
rect 212448 240032 212500 240038
rect 212448 239974 212500 239980
rect 212460 239329 212488 239974
rect 212446 239320 212502 239329
rect 212722 239320 212778 239329
rect 212446 239255 212502 239264
rect 212552 239278 212722 239306
rect 212552 239170 212580 239278
rect 212722 239255 212778 239264
rect 212184 239142 212580 239170
rect 211802 97200 211858 97209
rect 211802 97135 211858 97144
rect 210422 94480 210478 94489
rect 210422 94415 210478 94424
rect 212184 480 212212 239142
rect 213196 53281 213224 341158
rect 214562 330168 214618 330177
rect 214562 330103 214618 330112
rect 214576 90409 214604 330103
rect 214668 288289 214696 475351
rect 215942 474056 215998 474065
rect 215942 473991 215998 474000
rect 215956 399809 215984 473991
rect 218702 443048 218758 443057
rect 218702 442983 218758 442992
rect 218060 438932 218112 438938
rect 218060 438874 218112 438880
rect 218072 434790 218100 438874
rect 218060 434784 218112 434790
rect 218060 434726 218112 434732
rect 215942 399800 215998 399809
rect 215942 399735 215998 399744
rect 216036 382424 216088 382430
rect 216036 382366 216088 382372
rect 215944 341284 215996 341290
rect 215944 341226 215996 341232
rect 214654 288280 214710 288289
rect 214654 288215 214710 288224
rect 215666 224360 215722 224369
rect 215666 224295 215722 224304
rect 214562 90400 214618 90409
rect 214562 90335 214618 90344
rect 213182 53272 213238 53281
rect 213182 53207 213238 53216
rect 215680 480 215708 224295
rect 215956 224233 215984 341226
rect 216048 278186 216076 382366
rect 216126 347576 216182 347585
rect 216126 347511 216182 347520
rect 216036 278180 216088 278186
rect 216036 278122 216088 278128
rect 216140 265577 216168 347511
rect 217322 344312 217378 344321
rect 217322 344247 217378 344256
rect 216678 344176 216734 344185
rect 216678 344111 216734 344120
rect 216692 343670 216720 344111
rect 216680 343664 216732 343670
rect 216680 343606 216732 343612
rect 216126 265568 216182 265577
rect 216126 265503 216182 265512
rect 215942 224224 215998 224233
rect 215942 224159 215998 224168
rect 217336 100065 217364 344247
rect 218716 305969 218744 442983
rect 219452 402529 219480 480148
rect 224774 477592 224830 477601
rect 224774 477527 224830 477536
rect 224222 476776 224278 476785
rect 224222 476711 224278 476720
rect 222106 469840 222162 469849
rect 222106 469775 222162 469784
rect 222014 440872 222070 440881
rect 222014 440807 222070 440816
rect 221464 440292 221516 440298
rect 221464 440234 221516 440240
rect 221476 438938 221504 440234
rect 221464 438932 221516 438938
rect 221464 438874 221516 438880
rect 219438 402520 219494 402529
rect 219438 402455 219494 402464
rect 220082 339960 220138 339969
rect 220082 339895 220138 339904
rect 218702 305960 218758 305969
rect 218702 305895 218758 305904
rect 219254 203688 219310 203697
rect 219254 203623 219310 203632
rect 217322 100056 217378 100065
rect 217322 99991 217378 100000
rect 219268 480 219296 203623
rect 220096 35329 220124 339895
rect 222028 299441 222056 440807
rect 222120 328001 222148 469775
rect 223488 442128 223540 442134
rect 223488 442070 223540 442076
rect 223500 440298 223528 442070
rect 223488 440292 223540 440298
rect 223488 440234 223540 440240
rect 222842 343768 222898 343777
rect 222842 343703 222898 343712
rect 222106 327992 222162 328001
rect 222106 327927 222162 327936
rect 222014 299432 222070 299441
rect 222014 299367 222070 299376
rect 222856 272649 222884 343703
rect 224236 287745 224264 476711
rect 224788 410009 224816 477527
rect 224866 470112 224922 470121
rect 224866 470047 224922 470056
rect 224774 410000 224830 410009
rect 224774 409935 224830 409944
rect 224314 332344 224370 332353
rect 224314 332279 224370 332288
rect 224222 287736 224278 287745
rect 224222 287671 224278 287680
rect 222842 272640 222898 272649
rect 222842 272575 222898 272584
rect 224328 268433 224356 332279
rect 224880 327457 224908 470047
rect 225524 403073 225552 480148
rect 227720 478848 227772 478854
rect 227720 478790 227772 478796
rect 231214 478816 231270 478825
rect 227732 477601 227760 478790
rect 231214 478751 231270 478760
rect 228454 478680 228510 478689
rect 228454 478615 228510 478624
rect 227718 477592 227774 477601
rect 227718 477527 227774 477536
rect 227626 475688 227682 475697
rect 227626 475623 227682 475632
rect 227534 475008 227590 475017
rect 227534 474943 227590 474952
rect 227442 473104 227498 473113
rect 227442 473039 227498 473048
rect 227350 472968 227406 472977
rect 227350 472903 227406 472912
rect 227258 472288 227314 472297
rect 227258 472223 227314 472232
rect 226062 470384 226118 470393
rect 226062 470319 226118 470328
rect 225970 469976 226026 469985
rect 225970 469911 226026 469920
rect 225510 403064 225566 403073
rect 225510 402999 225566 403008
rect 225602 344992 225658 345001
rect 225602 344927 225658 344936
rect 225418 344448 225474 344457
rect 225418 344383 225474 344392
rect 224866 327448 224922 327457
rect 224866 327383 224922 327392
rect 225432 283393 225460 344383
rect 225418 283384 225474 283393
rect 225418 283319 225474 283328
rect 225616 271969 225644 344927
rect 225786 344040 225842 344049
rect 225786 343975 225842 343984
rect 225694 333432 225750 333441
rect 225694 333367 225750 333376
rect 225602 271960 225658 271969
rect 225602 271895 225658 271904
rect 224314 268424 224370 268433
rect 224314 268359 224370 268368
rect 225708 264217 225736 333367
rect 225800 283937 225828 343975
rect 225880 341148 225932 341154
rect 225880 341090 225932 341096
rect 225786 283928 225842 283937
rect 225786 283863 225842 283872
rect 225892 282878 225920 341090
rect 225984 328545 226012 469911
rect 225970 328536 226026 328545
rect 225970 328471 226026 328480
rect 226076 325281 226104 470319
rect 226246 470248 226302 470257
rect 226246 470183 226302 470192
rect 226154 442232 226210 442241
rect 226154 442167 226210 442176
rect 226062 325272 226118 325281
rect 226062 325207 226118 325216
rect 226168 295361 226196 442167
rect 226260 319297 226288 470183
rect 226982 454744 227038 454753
rect 226982 454679 227038 454688
rect 226890 444136 226946 444145
rect 226890 444071 226946 444080
rect 226904 443873 226932 444071
rect 226890 443864 226946 443873
rect 226890 443799 226946 443808
rect 226996 392737 227024 454679
rect 227166 440328 227222 440337
rect 227166 440263 227168 440272
rect 227220 440263 227222 440272
rect 227168 440234 227220 440240
rect 226982 392728 227038 392737
rect 226982 392663 227038 392672
rect 227272 363905 227300 472223
rect 227258 363896 227314 363905
rect 227258 363831 227314 363840
rect 227364 357921 227392 472903
rect 227350 357912 227406 357921
rect 227350 357847 227406 357856
rect 227456 355201 227484 473039
rect 227548 356833 227576 474943
rect 227534 356824 227590 356833
rect 227534 356759 227590 356768
rect 227442 355192 227498 355201
rect 227442 355127 227498 355136
rect 227074 351112 227130 351121
rect 227074 351047 227130 351056
rect 226982 330712 227038 330721
rect 226982 330647 227038 330656
rect 226246 319288 226302 319297
rect 226246 319223 226302 319232
rect 226154 295352 226210 295361
rect 226154 295287 226210 295296
rect 225880 282872 225932 282878
rect 225880 282814 225932 282820
rect 225694 264208 225750 264217
rect 225694 264143 225750 264152
rect 222750 230072 222806 230081
rect 222750 230007 222806 230016
rect 220082 35320 220138 35329
rect 220082 35255 220138 35264
rect 222764 480 222792 230007
rect 226338 221640 226394 221649
rect 226338 221575 226394 221584
rect 226352 480 226380 221575
rect 226996 95849 227024 330647
rect 227088 276321 227116 351047
rect 227166 346488 227222 346497
rect 227166 346423 227222 346432
rect 227180 318073 227208 346423
rect 227166 318064 227222 318073
rect 227166 317999 227222 318008
rect 227640 299169 227668 475623
rect 228178 475280 228234 475289
rect 228178 475215 228234 475224
rect 227626 299160 227682 299169
rect 227626 299095 227682 299104
rect 228192 297537 228220 475215
rect 228362 470520 228418 470529
rect 228362 470455 228418 470464
rect 228270 442776 228326 442785
rect 228270 442711 228326 442720
rect 228284 439142 228312 442711
rect 228272 439136 228324 439142
rect 228272 439078 228324 439084
rect 228376 406065 228404 470455
rect 228362 406056 228418 406065
rect 228362 405991 228418 406000
rect 228468 405793 228496 478615
rect 230112 478168 230164 478174
rect 230112 478110 230164 478116
rect 228822 475144 228878 475153
rect 228822 475079 228878 475088
rect 228638 472696 228694 472705
rect 228638 472631 228694 472640
rect 228546 472152 228602 472161
rect 228546 472087 228602 472096
rect 228454 405784 228510 405793
rect 228454 405719 228510 405728
rect 228560 364449 228588 472087
rect 228546 364440 228602 364449
rect 228546 364375 228602 364384
rect 228652 363361 228680 472631
rect 228732 439680 228784 439686
rect 228732 439622 228784 439628
rect 228744 439249 228772 439622
rect 228730 439240 228786 439249
rect 228730 439175 228786 439184
rect 228732 439136 228784 439142
rect 228732 439078 228784 439084
rect 228638 363352 228694 363361
rect 228638 363287 228694 363296
rect 228454 344584 228510 344593
rect 228454 344519 228510 344528
rect 228364 340944 228416 340950
rect 228364 340886 228416 340892
rect 228178 297528 228234 297537
rect 228178 297463 228234 297472
rect 227074 276312 227130 276321
rect 227074 276247 227130 276256
rect 226982 95840 227038 95849
rect 226982 95775 227038 95784
rect 228376 33969 228404 340886
rect 228468 281761 228496 344519
rect 228640 341080 228692 341086
rect 228640 341022 228692 341028
rect 228548 341012 228600 341018
rect 228548 340954 228600 340960
rect 228454 281752 228510 281761
rect 228454 281687 228510 281696
rect 228560 280158 228588 340954
rect 228652 281450 228680 341022
rect 228744 331401 228772 439078
rect 228836 357377 228864 475079
rect 230124 472954 230152 478110
rect 230386 475416 230442 475425
rect 230386 475351 230442 475360
rect 230202 474872 230258 474881
rect 230202 474807 230258 474816
rect 230032 472926 230152 472954
rect 229742 472560 229798 472569
rect 229742 472495 229798 472504
rect 229008 442196 229060 442202
rect 229008 442138 229060 442144
rect 229020 442105 229048 442138
rect 229006 442096 229062 442105
rect 229006 442031 229062 442040
rect 229650 442096 229706 442105
rect 229650 442031 229706 442040
rect 229664 441697 229692 442031
rect 229650 441688 229706 441697
rect 229650 441623 229706 441632
rect 229006 440872 229062 440881
rect 229006 440807 229062 440816
rect 228916 440428 228968 440434
rect 228916 440370 228968 440376
rect 228928 440337 228956 440370
rect 229020 440366 229048 440807
rect 229650 440736 229706 440745
rect 229650 440671 229706 440680
rect 229664 440502 229692 440671
rect 229652 440496 229704 440502
rect 229652 440438 229704 440444
rect 229008 440360 229060 440366
rect 228914 440328 228970 440337
rect 229008 440302 229060 440308
rect 228914 440263 228970 440272
rect 228914 440192 228970 440201
rect 228914 440127 228970 440136
rect 228822 357368 228878 357377
rect 228822 357303 228878 357312
rect 228824 341352 228876 341358
rect 228824 341294 228876 341300
rect 228730 331392 228786 331401
rect 228730 331327 228786 331336
rect 228836 281518 228864 341294
rect 228928 304065 228956 440127
rect 229650 440056 229706 440065
rect 229650 439991 229706 440000
rect 229376 439884 229428 439890
rect 229376 439826 229428 439832
rect 229388 439657 229416 439826
rect 229664 439657 229692 439991
rect 229374 439648 229430 439657
rect 229008 439612 229060 439618
rect 229374 439583 229430 439592
rect 229650 439648 229706 439657
rect 229650 439583 229706 439592
rect 229008 439554 229060 439560
rect 229020 439385 229048 439554
rect 229652 439476 229704 439482
rect 229652 439418 229704 439424
rect 229006 439376 229062 439385
rect 229006 439311 229062 439320
rect 229664 439113 229692 439418
rect 229650 439104 229706 439113
rect 229650 439039 229706 439048
rect 229756 340785 229784 472495
rect 230032 471918 230060 472926
rect 230110 472832 230166 472841
rect 230110 472767 230166 472776
rect 230020 471912 230072 471918
rect 230020 471854 230072 471860
rect 230018 439920 230074 439929
rect 230018 439855 230020 439864
rect 230072 439855 230074 439864
rect 230020 439826 230072 439832
rect 230124 361729 230152 472767
rect 230110 361720 230166 361729
rect 230110 361655 230166 361664
rect 230216 356289 230244 474807
rect 230400 473362 230428 475351
rect 230296 473340 230348 473346
rect 230400 473334 230520 473362
rect 230296 473282 230348 473288
rect 230308 472025 230336 473282
rect 230388 473272 230440 473278
rect 230388 473214 230440 473220
rect 230400 472433 230428 473214
rect 230386 472424 230442 472433
rect 230386 472359 230442 472368
rect 230492 472274 230520 473334
rect 230400 472246 230520 472274
rect 230294 472016 230350 472025
rect 230294 471951 230350 471960
rect 230296 471912 230348 471918
rect 230296 471854 230348 471860
rect 230202 356280 230258 356289
rect 230202 356215 230258 356224
rect 229742 340776 229798 340785
rect 229742 340711 229798 340720
rect 229756 329769 229784 340711
rect 230308 334121 230336 471854
rect 230294 334112 230350 334121
rect 230294 334047 230350 334056
rect 229834 331800 229890 331809
rect 229834 331735 229890 331744
rect 229742 329760 229798 329769
rect 229742 329695 229798 329704
rect 228914 304056 228970 304065
rect 228914 303991 228970 304000
rect 228824 281512 228876 281518
rect 228824 281454 228876 281460
rect 228640 281444 228692 281450
rect 228640 281386 228692 281392
rect 228548 280152 228600 280158
rect 228548 280094 228600 280100
rect 229848 269793 229876 331735
rect 230400 296993 230428 472246
rect 231122 464400 231178 464409
rect 231122 464335 231178 464344
rect 230480 440632 230532 440638
rect 230478 440600 230480 440609
rect 230532 440600 230534 440609
rect 230478 440535 230534 440544
rect 231032 439408 231084 439414
rect 231032 439350 231084 439356
rect 231044 439113 231072 439350
rect 231030 439104 231086 439113
rect 231030 439039 231086 439048
rect 231136 397633 231164 464335
rect 231228 404705 231256 478751
rect 231492 478372 231544 478378
rect 231492 478314 231544 478320
rect 231504 475674 231532 478314
rect 231412 475646 231532 475674
rect 231412 474366 231440 475646
rect 231490 475552 231546 475561
rect 231490 475487 231546 475496
rect 231400 474360 231452 474366
rect 231400 474302 231452 474308
rect 231306 474192 231362 474201
rect 231306 474127 231362 474136
rect 231214 404696 231270 404705
rect 231214 404631 231270 404640
rect 231122 397624 231178 397633
rect 231122 397559 231178 397568
rect 231320 366625 231348 474127
rect 231400 440564 231452 440570
rect 231400 440506 231452 440512
rect 231412 440337 231440 440506
rect 231398 440328 231454 440337
rect 231398 440263 231454 440272
rect 231400 439544 231452 439550
rect 231400 439486 231452 439492
rect 231306 366616 231362 366625
rect 231306 366551 231362 366560
rect 231214 364984 231270 364993
rect 231214 364919 231270 364928
rect 230938 342000 230994 342009
rect 230938 341935 230994 341944
rect 230386 296984 230442 296993
rect 230386 296919 230442 296928
rect 230952 279041 230980 341935
rect 231122 341320 231178 341329
rect 231122 341255 231178 341264
rect 230938 279032 230994 279041
rect 230938 278967 230994 278976
rect 231136 278497 231164 341255
rect 231228 301345 231256 364919
rect 231306 341864 231362 341873
rect 231306 341799 231362 341808
rect 231214 301336 231270 301345
rect 231214 301271 231270 301280
rect 231122 278488 231178 278497
rect 231122 278423 231178 278432
rect 231320 277953 231348 341799
rect 231412 324465 231440 439486
rect 231504 350305 231532 475487
rect 231596 403617 231624 480148
rect 234526 479632 234582 479641
rect 234526 479567 234582 479576
rect 231768 478780 231820 478786
rect 231768 478722 231820 478728
rect 231676 478236 231728 478242
rect 231676 478178 231728 478184
rect 231688 474450 231716 478178
rect 231780 477873 231808 478722
rect 233148 478712 233200 478718
rect 233148 478654 233200 478660
rect 231766 477864 231822 477873
rect 231766 477799 231822 477808
rect 233160 477737 233188 478654
rect 234344 478304 234396 478310
rect 234344 478246 234396 478252
rect 233146 477728 233202 477737
rect 233146 477663 233202 477672
rect 231860 475924 231912 475930
rect 231860 475866 231912 475872
rect 231872 475425 231900 475866
rect 233884 475720 233936 475726
rect 233884 475662 233936 475668
rect 231858 475416 231914 475425
rect 231858 475351 231914 475360
rect 232870 475416 232926 475425
rect 232870 475351 232926 475360
rect 233056 475380 233108 475386
rect 231688 474422 231808 474450
rect 231676 474360 231728 474366
rect 231676 474302 231728 474308
rect 231582 403608 231638 403617
rect 231582 403543 231638 403552
rect 231582 369880 231638 369889
rect 231582 369815 231638 369824
rect 231596 367713 231624 369815
rect 231582 367704 231638 367713
rect 231582 367639 231638 367648
rect 231490 350296 231546 350305
rect 231490 350231 231546 350240
rect 231490 341184 231546 341193
rect 231490 341119 231546 341128
rect 231398 324456 231454 324465
rect 231398 324391 231454 324400
rect 231504 279585 231532 341119
rect 231688 329089 231716 474302
rect 231674 329080 231730 329089
rect 231674 329015 231730 329024
rect 231780 320929 231808 474422
rect 232780 472660 232832 472666
rect 232780 472602 232832 472608
rect 232688 440700 232740 440706
rect 232688 440642 232740 440648
rect 232700 440337 232728 440642
rect 232686 440328 232742 440337
rect 232686 440263 232742 440272
rect 232792 369345 232820 472602
rect 232778 369336 232834 369345
rect 232778 369271 232834 369280
rect 232884 355745 232912 475351
rect 233056 475322 233108 475328
rect 232962 469704 233018 469713
rect 232962 469639 233018 469648
rect 232870 355736 232926 355745
rect 232870 355671 232926 355680
rect 232976 326913 233004 469639
rect 232962 326904 233018 326913
rect 232962 326839 233018 326848
rect 231766 320920 231822 320929
rect 231766 320855 231822 320864
rect 233068 313313 233096 475322
rect 233896 475289 233924 475662
rect 233882 475280 233938 475289
rect 233882 475215 233938 475224
rect 234250 475280 234306 475289
rect 234250 475215 234306 475224
rect 233146 465760 233202 465769
rect 233146 465695 233202 465704
rect 233054 313304 233110 313313
rect 233054 313239 233110 313248
rect 233160 296449 233188 465695
rect 234158 451888 234214 451897
rect 234158 451823 234214 451832
rect 233790 449168 233846 449177
rect 233790 449103 233846 449112
rect 233804 447134 233832 449103
rect 233804 447106 234108 447134
rect 233882 446448 233938 446457
rect 233804 446406 233882 446434
rect 233804 437474 233832 446406
rect 233882 446383 233938 446392
rect 233974 444952 234030 444961
rect 233896 444910 233974 444938
rect 233896 441266 233924 444910
rect 233974 444887 234030 444896
rect 233976 442944 234028 442950
rect 233976 442886 234028 442892
rect 233988 441697 234016 442886
rect 233974 441688 234030 441697
rect 233974 441623 234030 441632
rect 233896 441238 234016 441266
rect 233804 437446 233924 437474
rect 233896 313857 233924 437446
rect 233882 313848 233938 313857
rect 233882 313783 233938 313792
rect 233988 312769 234016 441238
rect 234080 314945 234108 447106
rect 234066 314936 234122 314945
rect 234066 314871 234122 314880
rect 233974 312760 234030 312769
rect 233974 312695 234030 312704
rect 234172 312225 234200 451823
rect 234264 322561 234292 475215
rect 234250 322552 234306 322561
rect 234250 322487 234306 322496
rect 234356 321473 234384 478246
rect 234434 471200 234490 471209
rect 234434 471135 234490 471144
rect 234342 321464 234398 321473
rect 234342 321399 234398 321408
rect 234448 313313 234476 471135
rect 234540 320385 234568 479567
rect 235632 475448 235684 475454
rect 235632 475390 235684 475396
rect 235446 458960 235502 458969
rect 235446 458895 235502 458904
rect 235078 453248 235134 453257
rect 235078 453183 235134 453192
rect 234986 448216 235042 448225
rect 234986 448151 235042 448160
rect 234894 440192 234950 440201
rect 234894 440127 234950 440136
rect 234908 439385 234936 440127
rect 234894 439376 234950 439385
rect 234894 439311 234950 439320
rect 235000 351937 235028 448151
rect 235092 368257 235120 453183
rect 235170 450664 235226 450673
rect 235170 450599 235226 450608
rect 235078 368248 235134 368257
rect 235078 368183 235134 368192
rect 235184 365537 235212 450599
rect 235354 445360 235410 445369
rect 235354 445295 235410 445304
rect 235262 443592 235318 443601
rect 235262 443527 235318 443536
rect 235170 365528 235226 365537
rect 235170 365463 235226 365472
rect 235276 353569 235304 443527
rect 235368 354657 235396 445295
rect 235460 364993 235488 458895
rect 235538 446856 235594 446865
rect 235538 446791 235594 446800
rect 235446 364984 235502 364993
rect 235446 364919 235502 364928
rect 235354 354648 235410 354657
rect 235354 354583 235410 354592
rect 235262 353560 235318 353569
rect 235262 353495 235318 353504
rect 235552 353025 235580 446791
rect 235644 444145 235672 475390
rect 237102 471336 237158 471345
rect 237102 471271 237158 471280
rect 235814 467256 235870 467265
rect 235814 467191 235870 467200
rect 235722 467120 235778 467129
rect 235722 467055 235778 467064
rect 235630 444136 235686 444145
rect 235630 444071 235686 444080
rect 235736 367713 235764 467055
rect 235722 367704 235778 367713
rect 235722 367639 235778 367648
rect 235828 367169 235856 467191
rect 235906 465896 235962 465905
rect 235906 465831 235962 465840
rect 235814 367160 235870 367169
rect 235814 367095 235870 367104
rect 235538 353016 235594 353025
rect 235538 352951 235594 352960
rect 234986 351928 235042 351937
rect 234986 351863 235042 351872
rect 235920 351393 235948 465831
rect 236918 464400 236974 464409
rect 236918 464335 236974 464344
rect 236826 460184 236882 460193
rect 236826 460119 236882 460128
rect 236734 448080 236790 448089
rect 236734 448015 236790 448024
rect 236642 447808 236698 447817
rect 236642 447743 236698 447752
rect 236458 445224 236514 445233
rect 236458 445159 236514 445168
rect 236472 362817 236500 445159
rect 236550 443728 236606 443737
rect 236550 443663 236606 443672
rect 236458 362808 236514 362817
rect 236458 362743 236514 362752
rect 236564 360641 236592 443663
rect 236550 360632 236606 360641
rect 236550 360567 236606 360576
rect 236656 360097 236684 447743
rect 236642 360088 236698 360097
rect 236642 360023 236698 360032
rect 236748 354113 236776 448015
rect 236840 359553 236868 460119
rect 236826 359544 236882 359553
rect 236826 359479 236882 359488
rect 236932 358465 236960 464335
rect 237010 462904 237066 462913
rect 237010 462839 237066 462848
rect 236918 358456 236974 358465
rect 236918 358391 236974 358400
rect 236734 354104 236790 354113
rect 236734 354039 236790 354048
rect 235906 351384 235962 351393
rect 235906 351319 235962 351328
rect 237024 350849 237052 462839
rect 237116 359009 237144 471271
rect 237194 468616 237250 468625
rect 237194 468551 237250 468560
rect 237102 359000 237158 359009
rect 237102 358935 237158 358944
rect 237208 352481 237236 468551
rect 237286 450800 237342 450809
rect 237286 450735 237342 450744
rect 237194 352472 237250 352481
rect 237194 352407 237250 352416
rect 237010 350840 237066 350849
rect 237010 350775 237066 350784
rect 235264 343664 235316 343670
rect 235264 343606 235316 343612
rect 234526 320376 234582 320385
rect 234526 320311 234582 320320
rect 234434 313304 234490 313313
rect 234434 313239 234490 313248
rect 234158 312216 234214 312225
rect 234158 312151 234214 312160
rect 235276 300830 235304 343606
rect 235814 341048 235870 341057
rect 235814 340983 235870 340992
rect 235828 324737 235856 340983
rect 235906 340912 235962 340921
rect 235906 340847 235962 340856
rect 235814 324728 235870 324737
rect 235814 324663 235870 324672
rect 235920 314401 235948 340847
rect 235906 314392 235962 314401
rect 235906 314327 235962 314336
rect 235906 307728 235962 307737
rect 235906 307663 235962 307672
rect 235264 300824 235316 300830
rect 235264 300766 235316 300772
rect 233146 296440 233202 296449
rect 233146 296375 233202 296384
rect 231490 279576 231546 279585
rect 231490 279511 231546 279520
rect 231306 277944 231362 277953
rect 231306 277879 231362 277888
rect 235920 277409 235948 307663
rect 237300 298625 237328 450735
rect 237378 443864 237434 443873
rect 237378 443799 237434 443808
rect 237562 443864 237618 443873
rect 237562 443799 237618 443808
rect 237392 443018 237420 443799
rect 237576 443601 237604 443799
rect 237562 443592 237618 443601
rect 237562 443527 237618 443536
rect 237380 443012 237432 443018
rect 237380 442954 237432 442960
rect 237668 404161 237696 480148
rect 243740 478825 243768 480148
rect 244830 479768 244886 479777
rect 244830 479703 244886 479712
rect 243726 478816 243782 478825
rect 243726 478751 243782 478760
rect 241428 478644 241480 478650
rect 241428 478586 241480 478592
rect 241440 478009 241468 478586
rect 241794 478544 241850 478553
rect 241794 478479 241850 478488
rect 241426 478000 241482 478009
rect 241426 477935 241482 477944
rect 238484 473204 238536 473210
rect 238484 473146 238536 473152
rect 238496 472025 238524 473146
rect 238482 472016 238538 472025
rect 238482 471951 238538 471960
rect 239494 454744 239550 454753
rect 239494 454679 239550 454688
rect 239402 446992 239458 447001
rect 239402 446927 239458 446936
rect 238574 446720 238630 446729
rect 238574 446655 238630 446664
rect 238298 443592 238354 443601
rect 238298 443527 238354 443536
rect 238022 443456 238078 443465
rect 238022 443391 238078 443400
rect 237654 404152 237710 404161
rect 237654 404087 237710 404096
rect 237378 384024 237434 384033
rect 237378 383959 237434 383968
rect 237392 383722 237420 383959
rect 237380 383716 237432 383722
rect 237380 383658 237432 383664
rect 237378 383480 237434 383489
rect 237378 383415 237434 383424
rect 237392 382566 237420 383415
rect 237470 382936 237526 382945
rect 237470 382871 237526 382880
rect 237380 382560 237432 382566
rect 237380 382502 237432 382508
rect 237378 382392 237434 382401
rect 237378 382327 237380 382336
rect 237432 382327 237434 382336
rect 237380 382298 237432 382304
rect 237484 382294 237512 382871
rect 237472 382288 237524 382294
rect 237472 382230 237524 382236
rect 237562 381848 237618 381857
rect 237562 381783 237618 381792
rect 237378 381304 237434 381313
rect 237378 381239 237434 381248
rect 237392 380934 237420 381239
rect 237576 381002 237604 381783
rect 237564 380996 237616 381002
rect 237564 380938 237616 380944
rect 237380 380928 237432 380934
rect 237380 380870 237432 380876
rect 237378 380760 237434 380769
rect 237378 380695 237434 380704
rect 237392 379574 237420 380695
rect 237380 379568 237432 379574
rect 237380 379510 237432 379516
rect 237746 378040 237802 378049
rect 237746 377975 237802 377984
rect 237562 377496 237618 377505
rect 237562 377431 237618 377440
rect 237378 376952 237434 376961
rect 237378 376887 237380 376896
rect 237432 376887 237434 376896
rect 237380 376858 237432 376864
rect 237576 376854 237604 377431
rect 237564 376848 237616 376854
rect 237564 376790 237616 376796
rect 237760 376786 237788 377975
rect 237748 376780 237800 376786
rect 237748 376722 237800 376728
rect 237562 376408 237618 376417
rect 237562 376343 237618 376352
rect 237378 375864 237434 375873
rect 237378 375799 237434 375808
rect 237392 375494 237420 375799
rect 237380 375488 237432 375494
rect 237380 375430 237432 375436
rect 237576 375426 237604 376343
rect 237564 375420 237616 375426
rect 237564 375362 237616 375368
rect 237378 375320 237434 375329
rect 237378 375255 237434 375264
rect 237392 374338 237420 375255
rect 237380 374332 237432 374338
rect 237380 374274 237432 374280
rect 237378 374232 237434 374241
rect 237378 374167 237434 374176
rect 237392 374066 237420 374167
rect 237380 374060 237432 374066
rect 237380 374002 237432 374008
rect 237378 371512 237434 371521
rect 237378 371447 237434 371456
rect 237392 371278 237420 371447
rect 237380 371272 237432 371278
rect 237380 371214 237432 371220
rect 237378 370968 237434 370977
rect 237378 370903 237434 370912
rect 237392 369918 237420 370903
rect 237380 369912 237432 369918
rect 237380 369854 237432 369860
rect 238036 366081 238064 443391
rect 238208 440972 238260 440978
rect 238208 440914 238260 440920
rect 238116 440904 238168 440910
rect 238116 440846 238168 440852
rect 238022 366072 238078 366081
rect 238022 366007 238078 366016
rect 237930 347712 237986 347721
rect 237930 347647 237986 347656
rect 237562 342136 237618 342145
rect 237562 342071 237618 342080
rect 237378 341592 237434 341601
rect 237378 341527 237434 341536
rect 237392 341222 237420 341527
rect 237576 341290 237604 342071
rect 237564 341284 237616 341290
rect 237564 341226 237616 341232
rect 237380 341216 237432 341222
rect 237380 341158 237432 341164
rect 237378 341048 237434 341057
rect 237378 340983 237434 340992
rect 237392 340950 237420 340983
rect 237380 340944 237432 340950
rect 237380 340886 237432 340892
rect 237838 340232 237894 340241
rect 237838 340167 237894 340176
rect 237378 320920 237434 320929
rect 237378 320855 237434 320864
rect 237392 316985 237420 320855
rect 237378 316976 237434 316985
rect 237378 316911 237434 316920
rect 237380 300824 237432 300830
rect 237378 300792 237380 300801
rect 237432 300792 237434 300801
rect 237378 300727 237434 300736
rect 237286 298616 237342 298625
rect 237286 298551 237342 298560
rect 237380 288380 237432 288386
rect 237380 288322 237432 288328
rect 237392 287201 237420 288322
rect 237378 287192 237434 287201
rect 237378 287127 237434 287136
rect 237380 287020 237432 287026
rect 237380 286962 237432 286968
rect 237392 286113 237420 286962
rect 237852 286657 237880 340167
rect 237944 325825 237972 347647
rect 238022 340096 238078 340105
rect 238022 340031 238078 340040
rect 237930 325816 237986 325825
rect 237930 325751 237986 325760
rect 237838 286648 237894 286657
rect 237838 286583 237894 286592
rect 237378 286104 237434 286113
rect 237378 286039 237434 286048
rect 237380 285660 237432 285666
rect 237380 285602 237432 285608
rect 237392 285569 237420 285602
rect 237378 285560 237434 285569
rect 237378 285495 237434 285504
rect 238036 284481 238064 340031
rect 238128 324193 238156 440846
rect 238114 324184 238170 324193
rect 238114 324119 238170 324128
rect 238220 322017 238248 440914
rect 238312 323649 238340 443527
rect 238484 442332 238536 442338
rect 238484 442274 238536 442280
rect 238392 441040 238444 441046
rect 238392 440982 238444 440988
rect 238298 323640 238354 323649
rect 238298 323575 238354 323584
rect 238206 322008 238262 322017
rect 238206 321943 238262 321952
rect 238404 319841 238432 440982
rect 238390 319832 238446 319841
rect 238390 319767 238446 319776
rect 238496 317665 238524 442274
rect 238588 320929 238616 446655
rect 239310 445496 239366 445505
rect 239310 445431 239366 445440
rect 238666 445088 238722 445097
rect 238666 445023 238722 445032
rect 238574 320920 238630 320929
rect 238574 320855 238630 320864
rect 238680 318753 238708 445023
rect 239126 444136 239182 444145
rect 239126 444071 239182 444080
rect 239034 442640 239090 442649
rect 239034 442575 239090 442584
rect 239048 406337 239076 442575
rect 239140 431954 239168 444071
rect 239220 441720 239272 441726
rect 239220 441662 239272 441668
rect 239232 436830 239260 441662
rect 239220 436824 239272 436830
rect 239220 436766 239272 436772
rect 239140 431926 239260 431954
rect 239232 406881 239260 431926
rect 239324 407425 239352 445431
rect 239416 407969 239444 446927
rect 239508 408513 239536 454679
rect 239678 449440 239734 449449
rect 239678 449375 239734 449384
rect 239586 447944 239642 447953
rect 239586 447879 239642 447888
rect 239494 408504 239550 408513
rect 239494 408439 239550 408448
rect 239402 407960 239458 407969
rect 239402 407895 239458 407904
rect 239310 407416 239366 407425
rect 239310 407351 239366 407360
rect 239218 406872 239274 406881
rect 239218 406807 239274 406816
rect 239034 406328 239090 406337
rect 239034 406263 239090 406272
rect 239494 405240 239550 405249
rect 239494 405175 239550 405184
rect 239508 401577 239536 405175
rect 239494 401568 239550 401577
rect 239494 401503 239550 401512
rect 239600 361185 239628 447879
rect 239692 362273 239720 449375
rect 240046 444272 240102 444281
rect 240046 444207 240102 444216
rect 240060 443086 240088 444207
rect 240048 443080 240100 443086
rect 240048 443022 240100 443028
rect 240046 442504 240102 442513
rect 240046 442439 240102 442448
rect 240060 442066 240088 442439
rect 240048 442060 240100 442066
rect 240048 442002 240100 442008
rect 239864 441788 239916 441794
rect 239864 441730 239916 441736
rect 239772 439748 239824 439754
rect 239772 439690 239824 439696
rect 239784 439113 239812 439690
rect 239770 439104 239826 439113
rect 239770 439039 239826 439048
rect 239772 436824 239824 436830
rect 239772 436766 239824 436772
rect 239678 362264 239734 362273
rect 239678 362199 239734 362208
rect 239586 361176 239642 361185
rect 239586 361111 239642 361120
rect 238666 318744 238722 318753
rect 238666 318679 238722 318688
rect 238482 317656 238538 317665
rect 238482 317591 238538 317600
rect 239784 300257 239812 436766
rect 239770 300248 239826 300257
rect 239770 300183 239826 300192
rect 239876 299713 239904 441730
rect 240784 440768 240836 440774
rect 240784 440710 240836 440716
rect 240796 439892 240824 440710
rect 241808 439892 241836 478479
rect 243544 476060 243596 476066
rect 243544 476002 243596 476008
rect 243556 475289 243584 476002
rect 243818 475824 243874 475833
rect 243818 475759 243874 475768
rect 243542 475280 243598 475289
rect 243542 475215 243598 475224
rect 242808 442060 242860 442066
rect 242808 442002 242860 442008
rect 242820 439892 242848 442002
rect 243832 439892 243860 475759
rect 244844 439892 244872 479703
rect 249812 478009 249840 480148
rect 255884 478689 255912 480148
rect 255870 478680 255926 478689
rect 255870 478615 255926 478624
rect 258998 478544 259054 478553
rect 258998 478479 259054 478488
rect 249798 478000 249854 478009
rect 249798 477935 249854 477944
rect 251088 475992 251140 475998
rect 249890 475960 249946 475969
rect 251088 475934 251140 475940
rect 249890 475895 249946 475904
rect 247866 473240 247922 473249
rect 247866 473175 247922 473184
rect 247040 473136 247092 473142
rect 247040 473078 247092 473084
rect 247052 472161 247080 473078
rect 247038 472152 247094 472161
rect 247038 472087 247094 472096
rect 246854 466032 246910 466041
rect 246854 465967 246910 465976
rect 245842 464536 245898 464545
rect 245842 464471 245898 464480
rect 245856 439892 245884 464471
rect 246868 439892 246896 465967
rect 247880 439892 247908 473175
rect 248878 460320 248934 460329
rect 248878 460255 248934 460264
rect 248892 439892 248920 460255
rect 249904 439892 249932 475895
rect 251100 475153 251128 475934
rect 251086 475144 251142 475153
rect 251086 475079 251142 475088
rect 257986 474328 258042 474337
rect 257986 474263 258042 474272
rect 255320 473068 255372 473074
rect 255320 473010 255372 473016
rect 255332 472297 255360 473010
rect 256054 472424 256110 472433
rect 256054 472359 256110 472368
rect 255318 472288 255374 472297
rect 255318 472223 255374 472232
rect 251914 471472 251970 471481
rect 251914 471407 251970 471416
rect 250902 442504 250958 442513
rect 250902 442439 250958 442448
rect 250916 439892 250944 442439
rect 251086 442232 251142 442241
rect 251086 442167 251142 442176
rect 251100 441930 251128 442167
rect 251088 441924 251140 441930
rect 251088 441866 251140 441872
rect 251928 439892 251956 471407
rect 252926 463040 252982 463049
rect 252926 462975 252982 462984
rect 252940 439892 252968 462975
rect 256068 451274 256096 472359
rect 256974 467528 257030 467537
rect 256974 467463 257030 467472
rect 255976 451246 256096 451274
rect 254030 442776 254086 442785
rect 254030 442711 254086 442720
rect 253938 442368 253994 442377
rect 253938 442303 253994 442312
rect 253952 441998 253980 442303
rect 254044 442066 254072 442711
rect 254398 442504 254454 442513
rect 254398 442439 254454 442448
rect 254032 442060 254084 442066
rect 254032 442002 254084 442008
rect 253940 441992 253992 441998
rect 253940 441934 253992 441940
rect 254412 441614 254440 442439
rect 254950 442368 255006 442377
rect 254950 442303 255006 442312
rect 254320 441586 254440 441614
rect 254320 439906 254348 441586
rect 253966 439878 254348 439906
rect 254964 439892 254992 442303
rect 255976 439892 256004 451246
rect 256988 439892 257016 467463
rect 258000 439892 258028 474263
rect 259012 439892 259040 478479
rect 260010 476912 260066 476921
rect 260010 476847 260066 476856
rect 260024 439892 260052 476847
rect 261022 459096 261078 459105
rect 261022 459031 261078 459040
rect 261036 439892 261064 459031
rect 261956 442649 261984 480148
rect 264058 479904 264114 479913
rect 264058 479839 264114 479848
rect 262034 478680 262090 478689
rect 262034 478615 262090 478624
rect 261942 442640 261998 442649
rect 261942 442575 261998 442584
rect 262048 439892 262076 478615
rect 263046 476096 263102 476105
rect 263046 476031 263102 476040
rect 262864 475856 262916 475862
rect 262864 475798 262916 475804
rect 262876 475017 262904 475798
rect 262862 475008 262918 475017
rect 262862 474943 262918 474952
rect 263060 439892 263088 476031
rect 264072 439892 264100 479839
rect 267094 478816 267150 478825
rect 267094 478751 267150 478760
rect 265070 442776 265126 442785
rect 265070 442711 265126 442720
rect 264978 442096 265034 442105
rect 264978 442031 265034 442040
rect 264992 441862 265020 442031
rect 264980 441856 265032 441862
rect 264980 441798 265032 441804
rect 265084 439892 265112 442711
rect 266082 442640 266138 442649
rect 266082 442575 266138 442584
rect 266096 439892 266124 442575
rect 267108 439892 267136 478751
rect 268028 444145 268056 480148
rect 268106 480040 268162 480049
rect 268106 479975 268162 479984
rect 268014 444136 268070 444145
rect 268014 444071 268070 444080
rect 267740 442128 267792 442134
rect 267740 442070 267792 442076
rect 267752 441590 267780 442070
rect 267740 441584 267792 441590
rect 267740 441526 267792 441532
rect 268120 439892 268148 479975
rect 271234 477048 271290 477057
rect 271234 476983 271290 476992
rect 271142 475280 271198 475289
rect 271142 475215 271198 475224
rect 269118 474464 269174 474473
rect 269118 474399 269174 474408
rect 269132 439892 269160 474399
rect 270130 442912 270186 442921
rect 270130 442847 270186 442856
rect 270144 439892 270172 442847
rect 270408 442128 270460 442134
rect 270408 442070 270460 442076
rect 270420 441969 270448 442070
rect 270406 441960 270462 441969
rect 270406 441895 270462 441904
rect 271156 439892 271184 475215
rect 271248 442921 271276 476983
rect 271788 475788 271840 475794
rect 271788 475730 271840 475736
rect 271800 474881 271828 475730
rect 271786 474872 271842 474881
rect 271786 474807 271842 474816
rect 273166 471608 273222 471617
rect 273166 471543 273222 471552
rect 271234 442912 271290 442921
rect 271234 442847 271290 442856
rect 272154 442912 272210 442921
rect 272154 442847 272210 442856
rect 272168 439892 272196 442847
rect 273180 439892 273208 471543
rect 274100 445505 274128 480148
rect 278226 480111 278282 480120
rect 276202 478000 276258 478009
rect 276202 477935 276258 477944
rect 275190 468752 275246 468761
rect 275190 468687 275246 468696
rect 274086 445496 274142 445505
rect 274086 445431 274142 445440
rect 274178 442096 274234 442105
rect 274178 442031 274234 442040
rect 273258 441824 273314 441833
rect 273258 441759 273314 441768
rect 273272 441658 273300 441759
rect 273260 441652 273312 441658
rect 273260 441594 273312 441600
rect 274192 439892 274220 442031
rect 275204 439892 275232 468687
rect 276216 439892 276244 477935
rect 277216 442400 277268 442406
rect 277216 442342 277268 442348
rect 277228 439892 277256 442342
rect 278240 439892 278268 480111
rect 279238 456240 279294 456249
rect 279238 456175 279294 456184
rect 279252 439892 279280 456175
rect 280172 447001 280200 480148
rect 286244 454753 286272 480148
rect 286230 454744 286286 454753
rect 286230 454679 286286 454688
rect 283010 453384 283066 453393
rect 283010 453319 283066 453328
rect 280158 446992 280214 447001
rect 280158 446927 280214 446936
rect 280436 442060 280488 442066
rect 280436 442002 280488 442008
rect 280448 441614 280476 442002
rect 280712 441992 280764 441998
rect 280712 441934 280764 441940
rect 280724 441614 280752 441934
rect 282920 441924 282972 441930
rect 282920 441866 282972 441872
rect 281080 441856 281132 441862
rect 281080 441798 281132 441804
rect 281092 441614 281120 441798
rect 280356 441586 280476 441614
rect 280540 441586 280752 441614
rect 280816 441586 281120 441614
rect 280252 440428 280304 440434
rect 280252 440370 280304 440376
rect 280160 439680 280212 439686
rect 280160 439622 280212 439628
rect 280068 439544 280120 439550
rect 280068 439486 280120 439492
rect 280080 397633 280108 439486
rect 280172 398993 280200 439622
rect 280264 400353 280292 440370
rect 280356 401713 280384 441586
rect 280540 440450 280568 441586
rect 280448 440422 280568 440450
rect 280448 403073 280476 440422
rect 280528 440360 280580 440366
rect 280528 440302 280580 440308
rect 280540 405793 280568 440302
rect 280620 439612 280672 439618
rect 280620 439554 280672 439560
rect 280526 405784 280582 405793
rect 280526 405719 280582 405728
rect 280632 404433 280660 439554
rect 280816 436778 280844 441586
rect 281906 441552 281962 441561
rect 281906 441487 281962 441496
rect 281080 440632 281132 440638
rect 281080 440574 281132 440580
rect 281630 440600 281686 440609
rect 280988 440496 281040 440502
rect 280988 440438 281040 440444
rect 280896 439476 280948 439482
rect 280896 439418 280948 439424
rect 280724 436750 280844 436778
rect 280724 407153 280752 436750
rect 280908 436642 280936 439418
rect 280816 436614 280936 436642
rect 280816 412593 280844 436614
rect 280896 436552 280948 436558
rect 280896 436494 280948 436500
rect 280908 413953 280936 436494
rect 281000 416673 281028 440438
rect 281092 436558 281120 440574
rect 281630 440535 281686 440544
rect 281538 440464 281594 440473
rect 281538 440399 281594 440408
rect 281080 436552 281132 436558
rect 281080 436494 281132 436500
rect 281552 434353 281580 440399
rect 281644 435713 281672 440535
rect 281722 440056 281778 440065
rect 281722 439991 281778 440000
rect 281630 435704 281686 435713
rect 281630 435639 281686 435648
rect 281632 435600 281684 435606
rect 281632 435542 281684 435548
rect 281538 434344 281594 434353
rect 281538 434279 281594 434288
rect 281540 434240 281592 434246
rect 281540 434182 281592 434188
rect 280986 416664 281042 416673
rect 280986 416599 281042 416608
rect 281552 415313 281580 434182
rect 281644 418033 281672 435542
rect 281736 419393 281764 439991
rect 281816 439408 281868 439414
rect 281816 439350 281868 439356
rect 281828 420753 281856 439350
rect 281920 432993 281948 441487
rect 282366 441416 282422 441425
rect 282366 441351 282422 441360
rect 282274 440872 282330 440881
rect 282274 440807 282330 440816
rect 282092 440700 282144 440706
rect 282092 440642 282144 440648
rect 282000 440564 282052 440570
rect 282000 440506 282052 440512
rect 282012 434246 282040 440506
rect 282104 435606 282132 440642
rect 282092 435600 282144 435606
rect 282092 435542 282144 435548
rect 282288 435282 282316 440807
rect 282104 435254 282316 435282
rect 282000 434240 282052 434246
rect 282000 434182 282052 434188
rect 282104 434058 282132 435254
rect 282012 434030 282132 434058
rect 281906 432984 281962 432993
rect 281906 432919 281962 432928
rect 282012 431954 282040 434030
rect 282380 433786 282408 441351
rect 282458 440192 282514 440201
rect 282458 440127 282514 440136
rect 281920 431926 282040 431954
rect 282104 433758 282408 433786
rect 281920 422113 281948 431926
rect 282104 424833 282132 433758
rect 282472 431954 282500 440127
rect 282196 431926 282500 431954
rect 282196 427553 282224 431926
rect 282182 427544 282238 427553
rect 282182 427479 282238 427488
rect 282090 424824 282146 424833
rect 282090 424759 282146 424768
rect 281906 422104 281962 422113
rect 281906 422039 281962 422048
rect 281814 420744 281870 420753
rect 281814 420679 281870 420688
rect 281722 419384 281778 419393
rect 281722 419319 281778 419328
rect 281630 418024 281686 418033
rect 281630 417959 281686 417968
rect 281538 415304 281594 415313
rect 281538 415239 281594 415248
rect 280894 413944 280950 413953
rect 280894 413879 280950 413888
rect 280802 412584 280858 412593
rect 280802 412519 280858 412528
rect 281906 409864 281962 409873
rect 281906 409799 281908 409808
rect 281960 409799 281962 409808
rect 281908 409770 281960 409776
rect 281906 408504 281962 408513
rect 281906 408439 281908 408448
rect 281960 408439 281962 408448
rect 281908 408410 281960 408416
rect 280710 407144 280766 407153
rect 280710 407079 280766 407088
rect 280618 404424 280674 404433
rect 280618 404359 280674 404368
rect 280434 403064 280490 403073
rect 280434 402999 280490 403008
rect 280342 401704 280398 401713
rect 280342 401639 280398 401648
rect 280250 400344 280306 400353
rect 280250 400279 280306 400288
rect 280158 398984 280214 398993
rect 280158 398919 280214 398928
rect 280066 397624 280122 397633
rect 280066 397559 280122 397568
rect 282826 395720 282882 395729
rect 282932 395706 282960 441866
rect 282882 395678 282960 395706
rect 282826 395655 282882 395664
rect 281816 394664 281868 394670
rect 281816 394606 281868 394612
rect 281828 393553 281856 394606
rect 281814 393544 281870 393553
rect 281814 393479 281870 393488
rect 280158 389464 280214 389473
rect 280158 389399 280214 389408
rect 239862 299704 239918 299713
rect 239862 299639 239918 299648
rect 280066 296984 280122 296993
rect 280066 296919 280122 296928
rect 239862 289368 239918 289377
rect 239862 289303 239918 289312
rect 239770 288824 239826 288833
rect 239770 288759 239826 288768
rect 238022 284472 238078 284481
rect 238022 284407 238078 284416
rect 237380 282872 237432 282878
rect 237380 282814 237432 282820
rect 237392 282305 237420 282814
rect 237378 282296 237434 282305
rect 237378 282231 237434 282240
rect 237564 281512 237616 281518
rect 237564 281454 237616 281460
rect 238666 281480 238722 281489
rect 237380 281444 237432 281450
rect 237380 281386 237432 281392
rect 237392 281217 237420 281386
rect 237378 281208 237434 281217
rect 237378 281143 237434 281152
rect 237576 280673 237604 281454
rect 238666 281415 238722 281424
rect 237562 280664 237618 280673
rect 237562 280599 237618 280608
rect 237380 280152 237432 280158
rect 237378 280120 237380 280129
rect 237432 280120 237434 280129
rect 237378 280055 237434 280064
rect 235906 277400 235962 277409
rect 235906 277335 235962 277344
rect 229834 269784 229890 269793
rect 229834 269719 229890 269728
rect 238680 240281 238708 281415
rect 238666 240272 238722 240281
rect 238666 240207 238722 240216
rect 236000 239964 236052 239970
rect 236000 239906 236052 239912
rect 236012 239057 236040 239906
rect 237472 239896 237524 239902
rect 237472 239838 237524 239844
rect 237380 239760 237432 239766
rect 237380 239702 237432 239708
rect 237010 239592 237066 239601
rect 237010 239527 237066 239536
rect 235998 239048 236054 239057
rect 235998 238983 236054 238992
rect 233422 237144 233478 237153
rect 233422 237079 233478 237088
rect 229834 228576 229890 228585
rect 229834 228511 229890 228520
rect 228362 33960 228418 33969
rect 228362 33895 228418 33904
rect 229848 480 229876 228511
rect 233436 480 233464 237079
rect 237024 480 237052 239527
rect 237392 239465 237420 239702
rect 237378 239456 237434 239465
rect 237378 239391 237434 239400
rect 237484 239193 237512 239838
rect 237564 239828 237616 239834
rect 237564 239770 237616 239776
rect 237470 239184 237526 239193
rect 237470 239119 237526 239128
rect 237576 238921 237604 239770
rect 237562 238912 237618 238921
rect 237562 238847 237618 238856
rect 239784 236609 239812 288759
rect 239770 236600 239826 236609
rect 239770 236535 239826 236544
rect 239876 235249 239904 289303
rect 280080 241913 280108 296919
rect 280066 241904 280122 241913
rect 280066 241839 280122 241848
rect 280066 241768 280122 241777
rect 280066 241703 280122 241712
rect 239862 235240 239918 235249
rect 239862 235175 239918 235184
rect 241440 5001 241468 240108
rect 242636 6225 242664 240108
rect 243832 238746 243860 240108
rect 243820 238740 243872 238746
rect 243820 238682 243872 238688
rect 245028 238678 245056 240108
rect 245016 238672 245068 238678
rect 245016 238614 245068 238620
rect 246224 237969 246252 240108
rect 247420 238105 247448 240108
rect 248616 238241 248644 240108
rect 249812 238377 249840 240108
rect 251008 238513 251036 240108
rect 252204 238649 252232 240108
rect 252190 238640 252246 238649
rect 252190 238575 252246 238584
rect 250994 238504 251050 238513
rect 250994 238439 251050 238448
rect 249798 238368 249854 238377
rect 249798 238303 249854 238312
rect 248602 238232 248658 238241
rect 248602 238167 248658 238176
rect 251178 238232 251234 238241
rect 251178 238167 251234 238176
rect 247406 238096 247462 238105
rect 247406 238031 247462 238040
rect 246210 237960 246266 237969
rect 246210 237895 246266 237904
rect 247590 237960 247646 237969
rect 247590 237895 247646 237904
rect 246302 69456 246358 69465
rect 246302 69391 246358 69400
rect 242622 6216 242678 6225
rect 242622 6151 242678 6160
rect 246316 5001 246344 69391
rect 241426 4992 241482 5001
rect 241426 4927 241482 4936
rect 246302 4992 246358 5001
rect 246302 4927 246358 4936
rect 243544 4140 243596 4146
rect 243544 4082 243596 4088
rect 240506 3904 240562 3913
rect 240506 3839 240562 3848
rect 240520 480 240548 3839
rect 243556 2961 243584 4082
rect 244094 4040 244150 4049
rect 244094 3975 244150 3984
rect 243542 2952 243598 2961
rect 243542 2887 243598 2896
rect 244108 480 244136 3975
rect 247604 480 247632 237895
rect 250442 78976 250498 78985
rect 250442 78911 250498 78920
rect 250456 50425 250484 78911
rect 250442 50416 250498 50425
rect 250442 50351 250498 50360
rect 251192 480 251220 238167
rect 253400 6361 253428 240108
rect 254596 38049 254624 240108
rect 254674 238096 254730 238105
rect 254674 238031 254730 238040
rect 254582 38040 254638 38049
rect 254582 37975 254638 37984
rect 253386 6352 253442 6361
rect 253386 6287 253442 6296
rect 254688 480 254716 238031
rect 255792 6497 255820 240108
rect 256988 6633 257016 240108
rect 258184 6769 258212 240108
rect 259276 239692 259328 239698
rect 259276 239634 259328 239640
rect 258262 239456 258318 239465
rect 258262 239391 258318 239400
rect 258170 6760 258226 6769
rect 258170 6695 258226 6704
rect 256974 6624 257030 6633
rect 256974 6559 257030 6568
rect 255778 6488 255834 6497
rect 255778 6423 255834 6432
rect 258276 480 258304 239391
rect 259288 238785 259316 239634
rect 259274 238776 259330 238785
rect 259274 238711 259330 238720
rect 259380 24313 259408 240108
rect 259366 24304 259422 24313
rect 259366 24239 259422 24248
rect 260576 20097 260604 240108
rect 261772 238754 261800 240108
rect 261680 238726 261800 238754
rect 260562 20088 260618 20097
rect 260562 20023 260618 20032
rect 261680 6905 261708 238726
rect 261758 238368 261814 238377
rect 261758 238303 261814 238312
rect 261666 6896 261722 6905
rect 261666 6831 261722 6840
rect 261772 480 261800 238303
rect 262968 6089 262996 240108
rect 264164 25673 264192 240108
rect 264980 239624 265032 239630
rect 264980 239566 265032 239572
rect 264992 239329 265020 239566
rect 264978 239320 265034 239329
rect 265360 239306 265388 240108
rect 264978 239255 265034 239264
rect 265268 239278 265388 239306
rect 265268 50561 265296 239278
rect 265346 239184 265402 239193
rect 265346 239119 265402 239128
rect 265254 50552 265310 50561
rect 265254 50487 265310 50496
rect 264150 25664 264206 25673
rect 264150 25599 264206 25608
rect 262954 6080 263010 6089
rect 262954 6015 263010 6024
rect 265360 480 265388 239119
rect 266556 91769 266584 240108
rect 267752 213217 267780 240108
rect 267738 213208 267794 213217
rect 267738 213143 267794 213152
rect 268948 211857 268976 240108
rect 268934 211848 268990 211857
rect 268934 211783 268990 211792
rect 270144 210361 270172 240108
rect 270130 210352 270186 210361
rect 270130 210287 270186 210296
rect 271340 177313 271368 240108
rect 272536 209001 272564 240108
rect 272522 208992 272578 209001
rect 272522 208927 272578 208936
rect 273732 178673 273760 240108
rect 273718 178664 273774 178673
rect 273718 178599 273774 178608
rect 271326 177304 271382 177313
rect 271326 177239 271382 177248
rect 274928 93129 274956 240108
rect 276124 238754 276152 240108
rect 275296 238726 276152 238754
rect 275296 207641 275324 238726
rect 275282 207632 275338 207641
rect 275282 207567 275338 207576
rect 277320 206281 277348 240108
rect 278516 237833 278544 240108
rect 278502 237824 278558 237833
rect 278502 237759 278558 237768
rect 277306 206272 277362 206281
rect 277306 206207 277362 206216
rect 274914 93120 274970 93129
rect 274914 93055 274970 93064
rect 266542 91760 266598 91769
rect 266542 91695 266598 91704
rect 275282 86048 275338 86057
rect 275282 85983 275338 85992
rect 271142 85912 271198 85921
rect 271142 85847 271198 85856
rect 268842 49056 268898 49065
rect 268842 48991 268898 49000
rect 268856 480 268884 48991
rect 271156 3369 271184 85847
rect 273902 54496 273958 54505
rect 273902 54431 273958 54440
rect 273916 5137 273944 54431
rect 275296 16574 275324 85983
rect 278042 21448 278098 21457
rect 278042 21383 278098 21392
rect 275296 16546 275968 16574
rect 273902 5128 273958 5137
rect 273902 5063 273958 5072
rect 271788 4072 271840 4078
rect 271788 4014 271840 4020
rect 271142 3360 271198 3369
rect 271142 3295 271198 3304
rect 271800 2825 271828 4014
rect 272430 3360 272486 3369
rect 272430 3295 272486 3304
rect 271786 2816 271842 2825
rect 271786 2751 271842 2760
rect 272444 480 272472 3295
rect 275940 3074 275968 16546
rect 278056 3369 278084 21383
rect 278042 3360 278098 3369
rect 278042 3295 278098 3304
rect 279514 3360 279570 3369
rect 279514 3295 279570 3304
rect 275940 3046 276060 3074
rect 276032 480 276060 3046
rect 279528 480 279556 3295
rect 280080 3233 280108 241703
rect 280172 239193 280200 389399
rect 280250 384024 280306 384033
rect 280250 383959 280306 383968
rect 280158 239184 280214 239193
rect 280158 239119 280214 239128
rect 280264 238241 280292 383959
rect 281722 382664 281778 382673
rect 281722 382599 281778 382608
rect 281630 381304 281686 381313
rect 281630 381239 281686 381248
rect 281538 379944 281594 379953
rect 281538 379879 281594 379888
rect 280434 378584 280490 378593
rect 280434 378519 280490 378528
rect 280342 373144 280398 373153
rect 280342 373079 280398 373088
rect 280250 238232 280306 238241
rect 280250 238167 280306 238176
rect 280356 230081 280384 373079
rect 280448 239601 280476 378519
rect 280526 367704 280582 367713
rect 280526 367639 280582 367648
rect 280434 239592 280490 239601
rect 280434 239527 280490 239536
rect 280540 232801 280568 367639
rect 280618 362264 280674 362273
rect 280618 362199 280674 362208
rect 280526 232792 280582 232801
rect 280526 232727 280582 232736
rect 280632 231305 280660 362199
rect 280710 358184 280766 358193
rect 280710 358119 280766 358128
rect 280724 235657 280752 358119
rect 280894 355464 280950 355473
rect 280894 355399 280950 355408
rect 280802 311944 280858 311953
rect 280802 311879 280858 311888
rect 280710 235648 280766 235657
rect 280710 235583 280766 235592
rect 280618 231296 280674 231305
rect 280618 231231 280674 231240
rect 280342 230072 280398 230081
rect 280342 230007 280398 230016
rect 280816 3913 280844 311879
rect 280908 239766 280936 355399
rect 281446 312080 281502 312089
rect 281446 312015 281502 312024
rect 281460 311794 281488 312015
rect 281552 311953 281580 379879
rect 281538 311944 281594 311953
rect 281538 311879 281594 311888
rect 281460 311766 281580 311794
rect 280986 299432 281042 299441
rect 280986 299367 281042 299376
rect 280896 239760 280948 239766
rect 280896 239702 280948 239708
rect 281000 4049 281028 299367
rect 281552 18737 281580 311766
rect 281644 299441 281672 381239
rect 281630 299432 281686 299441
rect 281630 299367 281686 299376
rect 281736 237969 281764 382599
rect 282826 369064 282882 369073
rect 282826 368999 282882 369008
rect 282840 368558 282868 368999
rect 282828 368552 282880 368558
rect 282828 368494 282880 368500
rect 281998 364984 282054 364993
rect 281998 364919 282054 364928
rect 281906 360904 281962 360913
rect 281906 360839 281962 360848
rect 281814 305144 281870 305153
rect 281814 305079 281870 305088
rect 281722 237960 281778 237969
rect 281722 237895 281778 237904
rect 281828 174593 281856 305079
rect 281920 229945 281948 360839
rect 282012 237017 282040 364919
rect 282826 359544 282882 359553
rect 282826 359479 282882 359488
rect 282840 358834 282868 359479
rect 282828 358828 282880 358834
rect 282828 358770 282880 358776
rect 282826 356824 282882 356833
rect 282826 356759 282882 356768
rect 282840 356114 282868 356759
rect 282828 356108 282880 356114
rect 282828 356050 282880 356056
rect 282826 354104 282882 354113
rect 282826 354039 282882 354048
rect 282840 353326 282868 354039
rect 282828 353320 282880 353326
rect 282828 353262 282880 353268
rect 282826 348664 282882 348673
rect 282826 348599 282882 348608
rect 282840 347818 282868 348599
rect 282828 347812 282880 347818
rect 282828 347754 282880 347760
rect 282826 344584 282882 344593
rect 282826 344519 282882 344528
rect 282840 343670 282868 344519
rect 282828 343664 282880 343670
rect 282828 343606 282880 343612
rect 282918 316024 282974 316033
rect 282918 315959 282974 315968
rect 282274 313304 282330 313313
rect 282274 313239 282330 313248
rect 282182 309224 282238 309233
rect 282182 309159 282238 309168
rect 282090 298344 282146 298353
rect 282090 298279 282146 298288
rect 281998 237008 282054 237017
rect 281998 236943 282054 236952
rect 281906 229936 281962 229945
rect 281906 229871 281962 229880
rect 282104 203561 282132 298279
rect 282196 214577 282224 309159
rect 282288 241074 282316 313239
rect 282366 310584 282422 310593
rect 282366 310519 282422 310528
rect 282380 241777 282408 310519
rect 282550 306504 282606 306513
rect 282550 306439 282606 306448
rect 282366 241768 282422 241777
rect 282366 241703 282422 241712
rect 282288 241046 282408 241074
rect 282274 240952 282330 240961
rect 282274 240887 282330 240896
rect 282288 240417 282316 240887
rect 282274 240408 282330 240417
rect 282274 240343 282330 240352
rect 282380 240106 282408 241046
rect 282368 240100 282420 240106
rect 282368 240042 282420 240048
rect 282182 214568 282238 214577
rect 282182 214503 282238 214512
rect 282090 203552 282146 203561
rect 282090 203487 282146 203496
rect 281814 174584 281870 174593
rect 281814 174519 281870 174528
rect 282564 36689 282592 306439
rect 282826 295624 282882 295633
rect 282826 295559 282882 295568
rect 282840 295390 282868 295559
rect 282828 295384 282880 295390
rect 282828 295326 282880 295332
rect 282828 281512 282880 281518
rect 282828 281454 282880 281460
rect 282840 280673 282868 281454
rect 282826 280664 282882 280673
rect 282826 280599 282882 280608
rect 282828 274644 282880 274650
rect 282828 274586 282880 274592
rect 282840 273873 282868 274586
rect 282826 273864 282882 273873
rect 282826 273799 282882 273808
rect 282828 273216 282880 273222
rect 282828 273158 282880 273164
rect 282840 272513 282868 273158
rect 282826 272504 282882 272513
rect 282826 272439 282882 272448
rect 282550 36680 282606 36689
rect 282550 36615 282606 36624
rect 282932 28393 282960 315959
rect 283024 275233 283052 453319
rect 288716 443080 288768 443086
rect 283102 443048 283158 443057
rect 288716 443022 288768 443028
rect 283102 442983 283158 442992
rect 288624 443012 288676 443018
rect 283116 411233 283144 442983
rect 288624 442954 288676 442960
rect 284484 442128 284536 442134
rect 284484 442070 284536 442076
rect 284392 441652 284444 441658
rect 284392 441594 284444 441600
rect 284300 440292 284352 440298
rect 284300 440234 284352 440240
rect 283102 411224 283158 411233
rect 283102 411159 283158 411168
rect 284312 394670 284340 440234
rect 284404 408474 284432 441594
rect 284496 409834 284524 442070
rect 287704 440768 287756 440774
rect 287704 440710 287756 440716
rect 284484 409828 284536 409834
rect 284484 409770 284536 409776
rect 284392 408468 284444 408474
rect 284392 408410 284444 408416
rect 284300 394664 284352 394670
rect 284300 394606 284352 394612
rect 283102 388104 283158 388113
rect 283102 388039 283158 388048
rect 283010 275224 283066 275233
rect 283010 275159 283066 275168
rect 283116 238377 283144 388039
rect 284482 385384 284538 385393
rect 284482 385319 284538 385328
rect 284390 374504 284446 374513
rect 284390 374439 284446 374448
rect 284298 371784 284354 371793
rect 284298 371719 284354 371728
rect 283286 366344 283342 366353
rect 283286 366279 283342 366288
rect 283194 345944 283250 345953
rect 283194 345879 283250 345888
rect 283102 238368 283158 238377
rect 283102 238303 283158 238312
rect 283208 196625 283236 345879
rect 283300 223009 283328 366279
rect 283378 363624 283434 363633
rect 283378 363559 283434 363568
rect 283392 234161 283420 363559
rect 283470 351384 283526 351393
rect 283470 351319 283526 351328
rect 283378 234152 283434 234161
rect 283378 234087 283434 234096
rect 283484 228449 283512 351319
rect 283562 350024 283618 350033
rect 283562 349959 283618 349968
rect 283576 236881 283604 349959
rect 283654 337784 283710 337793
rect 283654 337719 283710 337728
rect 283562 236872 283618 236881
rect 283562 236807 283618 236816
rect 283470 228440 283526 228449
rect 283470 228375 283526 228384
rect 283668 225729 283696 337719
rect 283746 336424 283802 336433
rect 283746 336359 283802 336368
rect 283760 232665 283788 336359
rect 283838 274680 283894 274689
rect 283838 274615 283894 274624
rect 283746 232656 283802 232665
rect 283746 232591 283802 232600
rect 283654 225720 283710 225729
rect 283654 225655 283710 225664
rect 283286 223000 283342 223009
rect 283286 222935 283342 222944
rect 283194 196616 283250 196625
rect 283194 196551 283250 196560
rect 282918 28384 282974 28393
rect 282918 28319 282974 28328
rect 281538 18728 281594 18737
rect 281538 18663 281594 18672
rect 283102 5128 283158 5137
rect 283102 5063 283158 5072
rect 280986 4040 281042 4049
rect 280986 3975 281042 3984
rect 280802 3904 280858 3913
rect 280802 3839 280858 3848
rect 280066 3224 280122 3233
rect 280066 3159 280122 3168
rect 283116 480 283144 5063
rect 283852 4078 283880 274615
rect 284312 203697 284340 371719
rect 284404 221649 284432 374439
rect 284496 243438 284524 385319
rect 284850 377224 284906 377233
rect 284850 377159 284906 377168
rect 284574 375864 284630 375873
rect 284574 375799 284630 375808
rect 284484 243432 284536 243438
rect 284484 243374 284536 243380
rect 284482 240136 284538 240145
rect 284482 240071 284538 240080
rect 284496 239426 284524 240071
rect 284484 239420 284536 239426
rect 284484 239362 284536 239368
rect 284588 228585 284616 375799
rect 284666 370424 284722 370433
rect 284666 370359 284722 370368
rect 284574 228576 284630 228585
rect 284574 228511 284630 228520
rect 284680 224369 284708 370359
rect 284758 343224 284814 343233
rect 284758 343159 284814 343168
rect 284666 224360 284722 224369
rect 284666 224295 284722 224304
rect 284390 221640 284446 221649
rect 284390 221575 284446 221584
rect 284298 203688 284354 203697
rect 284298 203623 284354 203632
rect 284772 197985 284800 343159
rect 284864 243574 284892 377159
rect 287152 368552 287204 368558
rect 287152 368494 287204 368500
rect 287058 352744 287114 352753
rect 287058 352679 287114 352688
rect 285034 347304 285090 347313
rect 285034 347239 285090 347248
rect 284942 340504 284998 340513
rect 284942 340439 284998 340448
rect 284852 243568 284904 243574
rect 284852 243510 284904 243516
rect 284852 243432 284904 243438
rect 284852 243374 284904 243380
rect 284864 238105 284892 243374
rect 284850 238096 284906 238105
rect 284850 238031 284906 238040
rect 284956 200705 284984 340439
rect 285048 231169 285076 347239
rect 285126 341864 285182 341873
rect 285126 341799 285182 341808
rect 285140 248414 285168 341799
rect 286138 333704 286194 333713
rect 286138 333639 286194 333648
rect 285862 329624 285918 329633
rect 285862 329559 285918 329568
rect 285678 321464 285734 321473
rect 285678 321399 285734 321408
rect 285140 248386 285260 248414
rect 285128 243568 285180 243574
rect 285128 243510 285180 243516
rect 285140 237153 285168 243510
rect 285126 237144 285182 237153
rect 285126 237079 285182 237088
rect 285232 235521 285260 248386
rect 285218 235512 285274 235521
rect 285218 235447 285274 235456
rect 285034 231160 285090 231169
rect 285034 231095 285090 231104
rect 284942 200696 284998 200705
rect 284942 200631 284998 200640
rect 284758 197976 284814 197985
rect 284758 197911 284814 197920
rect 285692 89049 285720 321399
rect 285770 320104 285826 320113
rect 285770 320039 285826 320048
rect 285784 204921 285812 320039
rect 285876 222873 285904 329559
rect 285954 324184 286010 324193
rect 285954 324119 286010 324128
rect 285862 222864 285918 222873
rect 285862 222799 285918 222808
rect 285968 221513 285996 324119
rect 286046 322824 286102 322833
rect 286046 322759 286102 322768
rect 285954 221504 286010 221513
rect 285954 221439 286010 221448
rect 286060 220153 286088 322759
rect 286152 232529 286180 333639
rect 286506 330984 286562 330993
rect 286506 330919 286562 330928
rect 286414 328264 286470 328273
rect 286414 328199 286470 328208
rect 286230 326904 286286 326913
rect 286230 326839 286286 326848
rect 286138 232520 286194 232529
rect 286138 232455 286194 232464
rect 286244 226953 286272 326839
rect 286322 325544 286378 325553
rect 286322 325479 286378 325488
rect 286336 229809 286364 325479
rect 286428 234025 286456 328199
rect 286520 236745 286548 330919
rect 286506 236736 286562 236745
rect 286506 236671 286562 236680
rect 286414 234016 286470 234025
rect 286414 233951 286470 233960
rect 286322 229800 286378 229809
rect 286322 229735 286378 229744
rect 286230 226944 286286 226953
rect 286230 226879 286286 226888
rect 286046 220144 286102 220153
rect 286046 220079 286102 220088
rect 285770 204912 285826 204921
rect 285770 204847 285826 204856
rect 285678 89040 285734 89049
rect 285678 88975 285734 88984
rect 284942 83464 284998 83473
rect 284942 83399 284998 83408
rect 283840 4072 283892 4078
rect 283840 4014 283892 4020
rect 284956 3369 284984 83399
rect 286598 4992 286654 5001
rect 286598 4927 286654 4936
rect 284942 3360 284998 3369
rect 284942 3295 284998 3304
rect 286612 480 286640 4927
rect 287072 3777 287100 352679
rect 287164 239630 287192 368494
rect 287244 356108 287296 356114
rect 287244 356050 287296 356056
rect 287256 239834 287284 356050
rect 287336 343664 287388 343670
rect 287336 343606 287388 343612
rect 287348 240038 287376 343606
rect 287426 288824 287482 288833
rect 287426 288759 287482 288768
rect 287440 241505 287468 288759
rect 287610 282976 287666 282985
rect 287610 282911 287666 282920
rect 287518 281888 287574 281897
rect 287518 281823 287574 281832
rect 287532 279313 287560 281823
rect 287518 279304 287574 279313
rect 287518 279239 287574 279248
rect 287624 277953 287652 282911
rect 287610 277944 287666 277953
rect 287610 277879 287666 277888
rect 287426 241496 287482 241505
rect 287426 241431 287482 241440
rect 287336 240032 287388 240038
rect 287336 239974 287388 239980
rect 287244 239828 287296 239834
rect 287244 239770 287296 239776
rect 287152 239624 287204 239630
rect 287152 239566 287204 239572
rect 287716 6866 287744 440710
rect 288438 332344 288494 332353
rect 288438 332279 288494 332288
rect 287704 6860 287756 6866
rect 287704 6802 287756 6808
rect 287058 3768 287114 3777
rect 287058 3703 287114 3712
rect 288452 3505 288480 332279
rect 288532 295384 288584 295390
rect 288532 295326 288584 295332
rect 288544 4146 288572 295326
rect 288636 273222 288664 442954
rect 288728 274650 288756 443022
rect 289004 442921 289032 480247
rect 289188 475969 289216 489886
rect 289464 485194 289492 491263
rect 289280 485166 289492 485194
rect 289174 475960 289230 475969
rect 289174 475895 289230 475904
rect 289280 464545 289308 485166
rect 289450 481128 289506 481137
rect 289450 481063 289506 481072
rect 289266 464536 289322 464545
rect 289266 464471 289322 464480
rect 288990 442912 289046 442921
rect 288990 442847 289046 442856
rect 289464 442406 289492 481063
rect 289556 473249 289584 499695
rect 289634 481536 289690 481545
rect 289634 481471 289690 481480
rect 289542 473240 289598 473249
rect 289542 473175 289598 473184
rect 289452 442400 289504 442406
rect 289452 442342 289504 442348
rect 288808 442196 288860 442202
rect 288808 442138 288860 442144
rect 288820 281518 288848 442138
rect 289648 442105 289676 481471
rect 289832 459105 289860 552327
rect 289924 479913 289952 564431
rect 290002 556200 290058 556209
rect 290002 556135 290058 556144
rect 289910 479904 289966 479913
rect 289910 479839 289966 479848
rect 290016 478689 290044 556135
rect 290094 548856 290150 548865
rect 290094 548791 290150 548800
rect 290002 478680 290058 478689
rect 290002 478615 290058 478624
rect 290108 476921 290136 548791
rect 290370 544776 290426 544785
rect 290370 544711 290426 544720
rect 290278 540696 290334 540705
rect 290278 540631 290334 540640
rect 290186 536616 290242 536625
rect 290186 536551 290242 536560
rect 290094 476912 290150 476921
rect 290094 476847 290150 476856
rect 290200 467537 290228 536551
rect 290292 474337 290320 540631
rect 290384 478553 290412 544711
rect 290462 532536 290518 532545
rect 290462 532471 290518 532480
rect 290370 478544 290426 478553
rect 290370 478479 290426 478488
rect 290278 474328 290334 474337
rect 290278 474263 290334 474272
rect 290476 472433 290504 532471
rect 291198 512136 291254 512145
rect 291198 512071 291254 512080
rect 291212 495530 291240 512071
rect 290568 495502 291240 495530
rect 290462 472424 290518 472433
rect 290462 472359 290518 472368
rect 290186 467528 290242 467537
rect 290186 467463 290242 467472
rect 289818 459096 289874 459105
rect 289818 459031 289874 459040
rect 289726 442912 289782 442921
rect 289726 442847 289782 442856
rect 289634 442096 289690 442105
rect 289634 442031 289690 442040
rect 289634 441960 289690 441969
rect 289634 441895 289690 441904
rect 289648 441726 289676 441895
rect 289740 441794 289768 442847
rect 290568 442241 290596 495502
rect 291198 495408 291254 495417
rect 291198 495343 291254 495352
rect 290646 487656 290702 487665
rect 290646 487591 290702 487600
rect 290660 479777 290688 487591
rect 290646 479768 290702 479777
rect 290646 479703 290702 479712
rect 291212 466041 291240 495343
rect 291304 481545 291332 605911
rect 291934 601896 291990 601905
rect 291934 601831 291990 601840
rect 291474 597816 291530 597825
rect 291474 597751 291530 597760
rect 291382 593736 291438 593745
rect 291382 593671 291438 593680
rect 291290 481536 291346 481545
rect 291290 481471 291346 481480
rect 291396 475289 291424 593671
rect 291488 480321 291516 597751
rect 291566 589656 291622 589665
rect 291566 589591 291622 589600
rect 291474 480312 291530 480321
rect 291474 480247 291530 480256
rect 291580 477057 291608 589591
rect 291658 585576 291714 585585
rect 291658 585511 291714 585520
rect 291566 477048 291622 477057
rect 291566 476983 291622 476992
rect 291382 475280 291438 475289
rect 291382 475215 291438 475224
rect 291672 474473 291700 585511
rect 291750 577416 291806 577425
rect 291750 577351 291806 577360
rect 291764 478825 291792 577351
rect 291842 520296 291898 520305
rect 291842 520231 291898 520240
rect 291750 478816 291806 478825
rect 291750 478751 291806 478760
rect 291658 474464 291714 474473
rect 291658 474399 291714 474408
rect 291198 466032 291254 466041
rect 291198 465967 291254 465976
rect 291856 463049 291884 520231
rect 291948 471617 291976 601831
rect 292026 503976 292082 503985
rect 292026 503911 292082 503920
rect 291934 471608 291990 471617
rect 291934 471543 291990 471552
rect 291842 463040 291898 463049
rect 291842 462975 291898 462984
rect 292040 460329 292068 503911
rect 292026 460320 292082 460329
rect 292026 460255 292082 460264
rect 290554 442232 290610 442241
rect 290554 442167 290610 442176
rect 289728 441788 289780 441794
rect 289728 441730 289780 441736
rect 289636 441720 289688 441726
rect 289636 441662 289688 441668
rect 288898 386744 288954 386753
rect 288898 386679 288954 386688
rect 288808 281512 288860 281518
rect 288808 281454 288860 281460
rect 288716 274644 288768 274650
rect 288716 274586 288768 274592
rect 288624 273216 288676 273222
rect 288624 273158 288676 273164
rect 288912 239465 288940 386679
rect 288992 358828 289044 358834
rect 288992 358770 289044 358776
rect 289004 239698 289032 358770
rect 289084 353320 289136 353326
rect 289084 353262 289136 353268
rect 289096 239902 289124 353262
rect 291292 347812 291344 347818
rect 291292 347754 291344 347760
rect 291198 335064 291254 335073
rect 291198 334999 291254 335008
rect 289084 239896 289136 239902
rect 289084 239838 289136 239844
rect 288992 239692 289044 239698
rect 288992 239634 289044 239640
rect 288898 239456 288954 239465
rect 288898 239391 288954 239400
rect 289084 87100 289136 87106
rect 289084 87042 289136 87048
rect 289096 7614 289124 87042
rect 289084 7608 289136 7614
rect 289084 7550 289136 7556
rect 290186 4856 290242 4865
rect 290186 4791 290242 4800
rect 288532 4140 288584 4146
rect 288532 4082 288584 4088
rect 288438 3496 288494 3505
rect 288438 3431 288494 3440
rect 290200 480 290228 4791
rect 291212 3641 291240 334999
rect 291304 239970 291332 347754
rect 292592 269793 292620 700567
rect 292776 442921 292804 700703
rect 292868 475697 292896 700975
rect 294050 700904 294106 700913
rect 294050 700839 294106 700848
rect 293222 700496 293278 700505
rect 293222 700431 293278 700440
rect 292946 633312 293002 633321
rect 292946 633247 293002 633256
rect 292960 478417 292988 633247
rect 293040 632256 293092 632262
rect 293040 632198 293092 632204
rect 293052 478718 293080 632198
rect 293130 524376 293186 524385
rect 293130 524311 293186 524320
rect 293040 478712 293092 478718
rect 293040 478654 293092 478660
rect 292946 478408 293002 478417
rect 292946 478343 293002 478352
rect 292854 475688 292910 475697
rect 292854 475623 292910 475632
rect 292762 442912 292818 442921
rect 292762 442847 292818 442856
rect 293144 442513 293172 524311
rect 293130 442504 293186 442513
rect 293130 442439 293186 442448
rect 293236 441969 293264 700431
rect 293958 700224 294014 700233
rect 293958 700159 294014 700168
rect 293222 441960 293278 441969
rect 293222 441895 293278 441904
rect 292578 269784 292634 269793
rect 292578 269719 292634 269728
rect 293972 267073 294000 700159
rect 294064 268433 294092 700839
rect 298742 700496 298798 700505
rect 298742 700431 298798 700440
rect 295338 700360 295394 700369
rect 295338 700295 295394 700304
rect 295982 700360 296038 700369
rect 295982 700295 296038 700304
rect 294144 632324 294196 632330
rect 294144 632266 294196 632272
rect 294156 478786 294184 632266
rect 294328 632188 294380 632194
rect 294328 632130 294380 632136
rect 294234 632088 294290 632097
rect 294234 632023 294290 632032
rect 294144 478780 294196 478786
rect 294144 478722 294196 478728
rect 294248 478281 294276 632023
rect 294340 478650 294368 632130
rect 294418 528456 294474 528465
rect 294418 528391 294474 528400
rect 294328 478644 294380 478650
rect 294328 478586 294380 478592
rect 294234 478272 294290 478281
rect 294234 478207 294290 478216
rect 294432 442377 294460 528391
rect 294510 483576 294566 483585
rect 294510 483511 294566 483520
rect 294524 475833 294552 483511
rect 294510 475824 294566 475833
rect 294510 475759 294566 475768
rect 294418 442368 294474 442377
rect 294418 442303 294474 442312
rect 295352 271153 295380 700295
rect 295430 569256 295486 569265
rect 295430 569191 295486 569200
rect 295444 442785 295472 569191
rect 295430 442776 295486 442785
rect 295430 442711 295486 442720
rect 295338 271144 295394 271153
rect 295338 271079 295394 271088
rect 294050 268424 294106 268433
rect 294050 268359 294106 268368
rect 293958 267064 294014 267073
rect 293958 266999 294014 267008
rect 295996 262993 296024 700295
rect 296718 573336 296774 573345
rect 296718 573271 296774 573280
rect 296732 442649 296760 573271
rect 296810 561096 296866 561105
rect 296810 561031 296866 561040
rect 296824 476105 296852 561031
rect 296810 476096 296866 476105
rect 296810 476031 296866 476040
rect 296718 442640 296774 442649
rect 296718 442575 296774 442584
rect 298756 264353 298784 700431
rect 300136 657257 300164 703520
rect 302882 700632 302938 700641
rect 302882 700567 302938 700576
rect 300122 657248 300178 657257
rect 300122 657183 300178 657192
rect 300136 635497 300164 657183
rect 300122 635488 300178 635497
rect 300122 635423 300178 635432
rect 300122 598224 300178 598233
rect 300122 598159 300178 598168
rect 300136 443465 300164 598159
rect 300122 443456 300178 443465
rect 300122 443391 300178 443400
rect 302896 265713 302924 700567
rect 332520 450809 332548 703520
rect 348804 700641 348832 703520
rect 348790 700632 348846 700641
rect 348790 700567 348846 700576
rect 353942 658880 353998 658889
rect 353942 658815 353998 658824
rect 332506 450800 332562 450809
rect 332506 450735 332562 450744
rect 302882 265704 302938 265713
rect 302882 265639 302938 265648
rect 298742 264344 298798 264353
rect 298742 264279 298798 264288
rect 295982 262984 296038 262993
rect 295982 262919 296038 262928
rect 353956 261633 353984 658815
rect 364996 657393 365024 703520
rect 364982 657384 365038 657393
rect 364982 657319 365038 657328
rect 364996 652089 365024 657319
rect 364982 652080 365038 652089
rect 364982 652015 365038 652024
rect 397472 449585 397500 703520
rect 413664 700505 413692 703520
rect 413650 700496 413706 700505
rect 413650 700431 413706 700440
rect 429856 657665 429884 703520
rect 429842 657656 429898 657665
rect 429842 657591 429898 657600
rect 429856 634273 429884 657591
rect 429842 634264 429898 634273
rect 429842 634199 429898 634208
rect 462332 475726 462360 703520
rect 478524 700369 478552 703520
rect 478510 700360 478566 700369
rect 478510 700295 478566 700304
rect 485044 700324 485096 700330
rect 485044 700266 485096 700272
rect 474646 657792 474702 657801
rect 474646 657727 474702 657736
rect 474660 634814 474688 657727
rect 474660 634786 474780 634814
rect 474752 634137 474780 634786
rect 474738 634128 474794 634137
rect 474738 634063 474794 634072
rect 462320 475720 462372 475726
rect 462320 475662 462372 475668
rect 397458 449576 397514 449585
rect 397458 449511 397514 449520
rect 474752 441590 474780 634063
rect 485056 475930 485084 700266
rect 494808 663794 494836 703520
rect 508502 700360 508558 700369
rect 527192 700330 527220 703520
rect 508502 700295 508558 700304
rect 527180 700324 527232 700330
rect 507122 670712 507178 670721
rect 507122 670647 507178 670656
rect 494624 663766 494836 663794
rect 489366 658064 489422 658073
rect 489366 657999 489422 658008
rect 487158 657792 487214 657801
rect 487158 657727 487214 657736
rect 486884 657416 486936 657422
rect 486884 657358 486936 657364
rect 486896 632874 486924 657358
rect 487172 657354 487200 657727
rect 487804 657552 487856 657558
rect 487804 657494 487856 657500
rect 487160 657348 487212 657354
rect 487160 657290 487212 657296
rect 487068 657008 487120 657014
rect 487068 656950 487120 656956
rect 486976 656940 487028 656946
rect 486976 656882 487028 656888
rect 486988 633418 487016 656882
rect 486976 633412 487028 633418
rect 486976 633354 487028 633360
rect 486884 632868 486936 632874
rect 486884 632810 486936 632816
rect 486896 632330 486924 632810
rect 486884 632324 486936 632330
rect 486884 632266 486936 632272
rect 486988 632194 487016 633354
rect 487080 632738 487108 656950
rect 487816 636857 487844 657494
rect 487896 657484 487948 657490
rect 487896 657426 487948 657432
rect 487908 642394 487936 657426
rect 489184 657144 489236 657150
rect 489184 657086 489236 657092
rect 488448 657076 488500 657082
rect 488448 657018 488500 657024
rect 487896 642388 487948 642394
rect 487896 642330 487948 642336
rect 488170 641200 488226 641209
rect 488170 641135 488226 641144
rect 487802 636848 487858 636857
rect 487802 636783 487858 636792
rect 487068 632732 487120 632738
rect 487068 632674 487120 632680
rect 487080 632262 487108 632674
rect 488080 632324 488132 632330
rect 488080 632266 488132 632272
rect 487068 632256 487120 632262
rect 487068 632198 487120 632204
rect 487988 632256 488040 632262
rect 487988 632198 488040 632204
rect 486976 632188 487028 632194
rect 486976 632130 487028 632136
rect 487896 632188 487948 632194
rect 487896 632130 487948 632136
rect 487802 613728 487858 613737
rect 487802 613663 487858 613672
rect 485044 475924 485096 475930
rect 485044 475866 485096 475872
rect 487816 472569 487844 613663
rect 487802 472560 487858 472569
rect 487802 472495 487858 472504
rect 474740 441584 474792 441590
rect 474740 441526 474792 441532
rect 474752 440298 474780 441526
rect 474740 440292 474792 440298
rect 474740 440234 474792 440240
rect 475384 440292 475436 440298
rect 475384 440234 475436 440240
rect 475396 344350 475424 440234
rect 475384 344344 475436 344350
rect 475384 344286 475436 344292
rect 353942 261624 353998 261633
rect 353942 261559 353998 261568
rect 291292 239964 291344 239970
rect 291292 239906 291344 239912
rect 291844 87304 291896 87310
rect 291844 87246 291896 87252
rect 291856 4826 291884 87246
rect 487908 86970 487936 632130
rect 488000 167006 488028 632198
rect 488092 245614 488120 632266
rect 488184 442950 488212 641135
rect 488460 632806 488488 657018
rect 489196 647902 489224 657086
rect 489276 655648 489328 655654
rect 489276 655590 489328 655596
rect 489184 647896 489236 647902
rect 489184 647838 489236 647844
rect 488448 632800 488500 632806
rect 488448 632742 488500 632748
rect 488460 632194 488488 632742
rect 488448 632188 488500 632194
rect 488448 632130 488500 632136
rect 489184 632188 489236 632194
rect 489184 632130 489236 632136
rect 488172 442944 488224 442950
rect 488172 442886 488224 442892
rect 488080 245608 488132 245614
rect 488080 245550 488132 245556
rect 489196 206990 489224 632130
rect 489288 442270 489316 655590
rect 489380 649233 489408 657999
rect 494624 657801 494652 663766
rect 505098 658064 505154 658073
rect 505098 657999 505154 658008
rect 494702 657928 494758 657937
rect 494702 657863 494758 657872
rect 494610 657792 494666 657801
rect 494610 657727 494666 657736
rect 490380 657280 490432 657286
rect 490380 657222 490432 657228
rect 490392 650690 490420 657222
rect 490472 657212 490524 657218
rect 490472 657154 490524 657160
rect 490484 653721 490512 657154
rect 493508 657008 493560 657014
rect 493508 656950 493560 656956
rect 492128 656940 492180 656946
rect 492128 656882 492180 656888
rect 492140 654908 492168 656882
rect 493520 654908 493548 656950
rect 494624 654809 494652 657727
rect 494716 656946 494744 657863
rect 496268 657416 496320 657422
rect 496268 657358 496320 657364
rect 503168 657416 503220 657422
rect 503168 657358 503220 657364
rect 494888 657076 494940 657082
rect 494888 657018 494940 657024
rect 494704 656940 494756 656946
rect 494704 656882 494756 656888
rect 494900 654908 494928 657018
rect 496280 654908 496308 657358
rect 497648 657348 497700 657354
rect 497648 657290 497700 657296
rect 497660 654908 497688 657290
rect 503180 656198 503208 657358
rect 505112 657354 505140 657999
rect 505100 657348 505152 657354
rect 505100 657290 505152 657296
rect 504548 656940 504600 656946
rect 504548 656882 504600 656888
rect 503168 656192 503220 656198
rect 503168 656134 503220 656140
rect 500408 655716 500460 655722
rect 500408 655658 500460 655664
rect 499028 655648 499080 655654
rect 499028 655590 499080 655596
rect 499040 654908 499068 655590
rect 500420 654945 500448 655658
rect 501788 655648 501840 655654
rect 501786 655616 501788 655625
rect 501840 655616 501842 655625
rect 501786 655551 501842 655560
rect 500406 654936 500462 654945
rect 501800 654908 501828 655551
rect 503180 654908 503208 656134
rect 504560 655790 504588 656882
rect 505926 656568 505982 656577
rect 505926 656503 505982 656512
rect 504548 655784 504600 655790
rect 504548 655726 504600 655732
rect 504560 654908 504588 655726
rect 505940 654908 505968 656503
rect 507136 655761 507164 670647
rect 508516 655897 508544 700295
rect 527180 700266 527232 700272
rect 543476 658889 543504 703520
rect 559668 700369 559696 703520
rect 559654 700360 559710 700369
rect 559654 700295 559710 700304
rect 580262 697232 580318 697241
rect 580262 697167 580318 697176
rect 543462 658880 543518 658889
rect 543462 658815 543518 658824
rect 510066 657792 510122 657801
rect 510066 657727 510122 657736
rect 508502 655888 508558 655897
rect 508502 655823 508558 655832
rect 507122 655752 507178 655761
rect 507122 655687 507178 655696
rect 507136 654922 507164 655687
rect 508516 654922 508544 655823
rect 507136 654894 507334 654922
rect 508516 654894 508714 654922
rect 510080 654908 510108 657727
rect 511446 657656 511502 657665
rect 511446 657591 511502 657600
rect 511460 654908 511488 657591
rect 534908 657552 534960 657558
rect 515586 657520 515642 657529
rect 534908 657494 534960 657500
rect 515586 657455 515642 657464
rect 512826 657384 512882 657393
rect 512826 657319 512882 657328
rect 512840 654908 512868 657319
rect 514206 657248 514262 657257
rect 514206 657183 514262 657192
rect 514220 654908 514248 657183
rect 514760 656940 514812 656946
rect 514760 656882 514812 656888
rect 500406 654871 500462 654880
rect 514772 654838 514800 656882
rect 515600 654908 515628 657455
rect 530768 657348 530820 657354
rect 530768 657290 530820 657296
rect 529388 657280 529440 657286
rect 529388 657222 529440 657228
rect 516966 657112 517022 657121
rect 516966 657047 517022 657056
rect 516980 654908 517008 657047
rect 526628 656940 526680 656946
rect 526628 656882 526680 656888
rect 525246 656432 525302 656441
rect 525246 656367 525302 656376
rect 522486 656296 522542 656305
rect 522486 656231 522542 656240
rect 519726 656160 519782 656169
rect 519726 656095 519782 656104
rect 518346 656024 518402 656033
rect 518346 655959 518402 655968
rect 518360 654908 518388 655959
rect 519740 654908 519768 656095
rect 522500 654908 522528 656231
rect 525260 654908 525288 656367
rect 526640 654908 526668 656882
rect 528008 655580 528060 655586
rect 528008 655522 528060 655528
rect 528020 654908 528048 655522
rect 529400 654908 529428 657222
rect 530780 654908 530808 657290
rect 533528 657212 533580 657218
rect 533528 657154 533580 657160
rect 532148 657144 532200 657150
rect 532148 657086 532200 657092
rect 532160 654908 532188 657086
rect 533540 654908 533568 657154
rect 534920 654908 534948 657494
rect 537668 657484 537720 657490
rect 537668 657426 537720 657432
rect 537680 654908 537708 657426
rect 577504 655716 577556 655722
rect 577504 655658 577556 655664
rect 514760 654832 514812 654838
rect 494610 654800 494666 654809
rect 514760 654774 514812 654780
rect 494610 654735 494666 654744
rect 523866 654664 523922 654673
rect 523866 654599 523922 654608
rect 536012 654560 536064 654566
rect 521106 654528 521162 654537
rect 536064 654508 536314 654514
rect 536012 654502 536314 654508
rect 536024 654486 536314 654502
rect 538784 654498 539074 654514
rect 538772 654492 539074 654498
rect 521106 654463 521162 654472
rect 538824 654486 539074 654492
rect 538772 654434 538824 654440
rect 490576 654214 490774 654242
rect 490470 653712 490526 653721
rect 490470 653647 490526 653656
rect 490380 650684 490432 650690
rect 490380 650626 490432 650632
rect 489366 649224 489422 649233
rect 489366 649159 489422 649168
rect 490576 632126 490604 654214
rect 540150 651264 540206 651273
rect 540150 651199 540206 651208
rect 539782 642560 539838 642569
rect 539782 642495 539838 642504
rect 539598 637800 539654 637809
rect 539598 637735 539654 637744
rect 490564 632120 490616 632126
rect 490564 632062 490616 632068
rect 490576 594114 490604 632062
rect 490564 594108 490616 594114
rect 490564 594050 490616 594056
rect 490760 475561 490788 600100
rect 490746 475552 490802 475561
rect 490746 475487 490802 475496
rect 492140 462913 492168 600100
rect 493520 465905 493548 600100
rect 493506 465896 493562 465905
rect 493506 465831 493562 465840
rect 492126 462904 492182 462913
rect 492126 462839 492182 462848
rect 494900 448225 494928 600100
rect 496280 468625 496308 600100
rect 496266 468616 496322 468625
rect 496266 468551 496322 468560
rect 494886 448216 494942 448225
rect 494886 448151 494942 448160
rect 497660 446865 497688 600100
rect 497646 446856 497702 446865
rect 497646 446791 497702 446800
rect 499040 443873 499068 600100
rect 500420 448089 500448 600100
rect 500406 448080 500462 448089
rect 500406 448015 500462 448024
rect 501800 445369 501828 600100
rect 503180 473113 503208 600100
rect 504560 475425 504588 600100
rect 505940 475794 505968 600100
rect 507320 475862 507348 600100
rect 508700 475998 508728 600100
rect 508688 475992 508740 475998
rect 508688 475934 508740 475940
rect 507308 475856 507360 475862
rect 507308 475798 507360 475804
rect 505928 475788 505980 475794
rect 505928 475730 505980 475736
rect 504546 475416 504602 475425
rect 504546 475351 504602 475360
rect 503166 473104 503222 473113
rect 503166 473039 503222 473048
rect 510080 472977 510108 600100
rect 511264 594108 511316 594114
rect 511264 594050 511316 594056
rect 510066 472968 510122 472977
rect 510066 472903 510122 472912
rect 501786 445360 501842 445369
rect 501786 445295 501842 445304
rect 499026 443864 499082 443873
rect 499026 443799 499082 443808
rect 489276 442264 489328 442270
rect 489276 442206 489328 442212
rect 489288 366382 489316 442206
rect 489276 366376 489328 366382
rect 489276 366318 489328 366324
rect 498844 366376 498896 366382
rect 498844 366318 498896 366324
rect 498856 353258 498884 366318
rect 498844 353252 498896 353258
rect 498844 353194 498896 353200
rect 497464 344344 497516 344350
rect 497464 344286 497516 344292
rect 497476 299470 497504 344286
rect 497464 299464 497516 299470
rect 497464 299406 497516 299412
rect 489184 206984 489236 206990
rect 489184 206926 489236 206932
rect 487988 167000 488040 167006
rect 487988 166942 488040 166948
rect 487896 86964 487948 86970
rect 487896 86906 487948 86912
rect 311438 86184 311494 86193
rect 311438 86119 311494 86128
rect 304354 51776 304410 51785
rect 304354 51711 304410 51720
rect 293682 46336 293738 46345
rect 293682 46271 293738 46280
rect 291844 4820 291896 4826
rect 291844 4762 291896 4768
rect 291198 3632 291254 3641
rect 291198 3567 291254 3576
rect 293696 480 293724 46271
rect 297270 43616 297326 43625
rect 297270 43551 297326 43560
rect 297284 480 297312 43551
rect 300766 42256 300822 42265
rect 300766 42191 300822 42200
rect 300780 480 300808 42191
rect 304368 480 304396 51711
rect 307942 50280 307998 50289
rect 307942 50215 307998 50224
rect 307956 480 307984 50215
rect 311452 480 311480 86119
rect 322110 85776 322166 85785
rect 322110 85711 322166 85720
rect 318522 80744 318578 80753
rect 318522 80679 318578 80688
rect 315026 53136 315082 53145
rect 315026 53071 315082 53080
rect 315040 480 315068 53071
rect 318536 480 318564 80679
rect 322124 480 322152 85711
rect 336278 85640 336334 85649
rect 336278 85575 336334 85584
rect 325606 69592 325662 69601
rect 325606 69527 325662 69536
rect 325620 480 325648 69527
rect 329194 54632 329250 54641
rect 329194 54567 329250 54576
rect 329208 480 329236 54567
rect 332690 9072 332746 9081
rect 332690 9007 332746 9016
rect 332704 480 332732 9007
rect 336292 480 336320 85575
rect 368202 84960 368258 84969
rect 368202 84895 368258 84904
rect 357530 84824 357586 84833
rect 357530 84759 357586 84768
rect 343362 84688 343418 84697
rect 343362 84623 343418 84632
rect 339868 83496 339920 83502
rect 339868 83438 339920 83444
rect 339880 480 339908 83438
rect 343376 480 343404 84623
rect 353942 57216 353998 57225
rect 353942 57151 353998 57160
rect 351182 55856 351238 55865
rect 351182 55791 351238 55800
rect 350448 51740 350500 51746
rect 350448 51682 350500 51688
rect 346952 4820 347004 4826
rect 346952 4762 347004 4768
rect 346964 480 346992 4762
rect 350460 480 350488 51682
rect 351196 4865 351224 55791
rect 353956 7585 353984 57151
rect 354036 7608 354088 7614
rect 353942 7576 353998 7585
rect 354036 7550 354088 7556
rect 353942 7511 353998 7520
rect 351182 4856 351238 4865
rect 351182 4791 351238 4800
rect 354048 480 354076 7550
rect 357544 480 357572 84759
rect 361118 84552 361174 84561
rect 361118 84487 361174 84496
rect 361132 480 361160 84487
rect 364616 79348 364668 79354
rect 364616 79290 364668 79296
rect 364628 480 364656 79290
rect 368216 480 368244 84895
rect 435362 83056 435418 83065
rect 435362 82991 435418 83000
rect 432602 81696 432658 81705
rect 432602 81631 432658 81640
rect 428554 80336 428610 80345
rect 428554 80271 428610 80280
rect 421562 77616 421618 77625
rect 421562 77551 421618 77560
rect 417422 76256 417478 76265
rect 417422 76191 417478 76200
rect 414662 74896 414718 74905
rect 414662 74831 414718 74840
rect 406382 64016 406438 64025
rect 406382 63951 406438 63960
rect 400126 40760 400182 40769
rect 400126 40695 400182 40704
rect 378874 21312 378930 21321
rect 378874 21247 378930 21256
rect 375286 10432 375342 10441
rect 375286 10367 375342 10376
rect 371698 3360 371754 3369
rect 371698 3295 371754 3304
rect 371712 480 371740 3295
rect 375300 480 375328 10367
rect 378888 480 378916 21247
rect 396538 17368 396594 17377
rect 396538 17303 396594 17312
rect 393042 16008 393098 16017
rect 393042 15943 393098 15952
rect 389454 14648 389510 14657
rect 389454 14583 389510 14592
rect 385958 13152 386014 13161
rect 385958 13087 386014 13096
rect 382370 11792 382426 11801
rect 382370 11727 382426 11736
rect 382384 480 382412 11727
rect 385972 480 386000 13087
rect 389468 480 389496 14583
rect 393056 480 393084 15943
rect 396552 480 396580 17303
rect 400140 480 400168 40695
rect 403622 22808 403678 22817
rect 403622 22743 403678 22752
rect 403636 480 403664 22743
rect 406396 7721 406424 63951
rect 411902 58576 411958 58585
rect 411902 58511 411958 58520
rect 407210 39400 407266 39409
rect 407210 39335 407266 39344
rect 406382 7712 406438 7721
rect 406382 7647 406438 7656
rect 407224 480 407252 39335
rect 411916 4865 411944 58511
rect 414294 7576 414350 7585
rect 414294 7511 414350 7520
rect 410798 4856 410854 4865
rect 410798 4791 410854 4800
rect 411902 4856 411958 4865
rect 411902 4791 411958 4800
rect 410812 480 410840 4791
rect 414308 480 414336 7511
rect 414676 3097 414704 74831
rect 417436 3505 417464 76191
rect 418802 59936 418858 59945
rect 418802 59871 418858 59880
rect 417882 4856 417938 4865
rect 417882 4791 417938 4800
rect 417422 3496 417478 3505
rect 417422 3431 417478 3440
rect 414662 3088 414718 3097
rect 414662 3023 414718 3032
rect 417896 480 417924 4791
rect 418816 4185 418844 59871
rect 418802 4176 418858 4185
rect 418802 4111 418858 4120
rect 421378 4176 421434 4185
rect 421378 4111 421434 4120
rect 421392 480 421420 4111
rect 421576 3913 421604 77551
rect 425702 62656 425758 62665
rect 425702 62591 425758 62600
rect 422942 61296 422998 61305
rect 422942 61231 422998 61240
rect 422956 4185 422984 61231
rect 425716 4185 425744 62591
rect 422942 4176 422998 4185
rect 422942 4111 422998 4120
rect 424966 4176 425022 4185
rect 424966 4111 425022 4120
rect 425702 4176 425758 4185
rect 425702 4111 425758 4120
rect 428462 4176 428518 4185
rect 428462 4111 428518 4120
rect 421562 3904 421618 3913
rect 421562 3839 421618 3848
rect 424980 480 425008 4111
rect 428476 480 428504 4111
rect 428568 3777 428596 80271
rect 431222 68096 431278 68105
rect 431222 68031 431278 68040
rect 429842 65376 429898 65385
rect 429842 65311 429898 65320
rect 429856 4865 429884 65311
rect 431236 7585 431264 68031
rect 432050 7712 432106 7721
rect 432050 7647 432106 7656
rect 431222 7576 431278 7585
rect 431222 7511 431278 7520
rect 429842 4856 429898 4865
rect 429842 4791 429898 4800
rect 428554 3768 428610 3777
rect 428554 3703 428610 3712
rect 432064 480 432092 7647
rect 432616 3233 432644 81631
rect 435376 3641 435404 82991
rect 450542 73536 450598 73545
rect 450542 73471 450598 73480
rect 447782 72176 447838 72185
rect 447782 72111 447838 72120
rect 443642 70816 443698 70825
rect 443642 70751 443698 70760
rect 436742 66736 436798 66745
rect 436742 66671 436798 66680
rect 435546 4856 435602 4865
rect 435546 4791 435602 4800
rect 435362 3632 435418 3641
rect 435362 3567 435418 3576
rect 432602 3224 432658 3233
rect 432602 3159 432658 3168
rect 435560 480 435588 4791
rect 436756 4185 436784 66671
rect 439502 47832 439558 47841
rect 439502 47767 439558 47776
rect 436742 4176 436798 4185
rect 436742 4111 436798 4120
rect 439134 4176 439190 4185
rect 439134 4111 439190 4120
rect 439148 480 439176 4111
rect 439516 4049 439544 47767
rect 442262 47696 442318 47705
rect 442262 47631 442318 47640
rect 439502 4040 439558 4049
rect 439502 3975 439558 3984
rect 442276 3369 442304 47631
rect 442630 7576 442686 7585
rect 442630 7511 442686 7520
rect 442262 3360 442318 3369
rect 442262 3295 442318 3304
rect 442644 480 442672 7511
rect 443656 4185 443684 70751
rect 446402 47560 446458 47569
rect 446402 47495 446458 47504
rect 443642 4176 443698 4185
rect 443642 4111 443698 4120
rect 446218 4176 446274 4185
rect 446218 4111 446274 4120
rect 442906 4040 442962 4049
rect 442906 3975 442962 3984
rect 442920 2854 442948 3975
rect 442908 2848 442960 2854
rect 442908 2790 442960 2796
rect 446232 480 446260 4111
rect 446416 3466 446444 47495
rect 447796 4185 447824 72111
rect 450556 4865 450584 73471
rect 467470 50416 467526 50425
rect 467470 50351 467526 50360
rect 450542 4856 450598 4865
rect 450542 4791 450598 4800
rect 453302 4856 453358 4865
rect 453302 4791 453358 4800
rect 447782 4176 447838 4185
rect 447782 4111 447838 4120
rect 449806 4176 449862 4185
rect 449806 4111 449862 4120
rect 446404 3460 446456 3466
rect 446404 3402 446456 3408
rect 449820 480 449848 4111
rect 453316 480 453344 4791
rect 463974 3904 464030 3913
rect 463974 3839 464030 3848
rect 460386 3496 460442 3505
rect 460386 3431 460442 3440
rect 456890 3088 456946 3097
rect 456890 3023 456946 3032
rect 456904 480 456932 3023
rect 460400 480 460428 3431
rect 463988 480 464016 3839
rect 467484 480 467512 50351
rect 511276 46918 511304 594050
rect 511460 464409 511488 600100
rect 512840 471345 512868 600100
rect 512826 471336 512882 471345
rect 512826 471271 512882 471280
rect 511446 464400 511502 464409
rect 511446 464335 511502 464344
rect 514220 460193 514248 600100
rect 514206 460184 514262 460193
rect 514206 460119 514262 460128
rect 515600 447817 515628 600100
rect 515586 447808 515642 447817
rect 515586 447743 515642 447752
rect 516980 443737 517008 600100
rect 518360 447953 518388 600100
rect 519740 472841 519768 600100
rect 519726 472832 519782 472841
rect 519726 472767 519782 472776
rect 521120 449449 521148 600100
rect 521106 449440 521162 449449
rect 521106 449375 521162 449384
rect 518346 447944 518402 447953
rect 518346 447879 518402 447888
rect 522500 445233 522528 600100
rect 523880 472705 523908 600100
rect 525260 473074 525288 600100
rect 526640 473142 526668 600100
rect 526628 473136 526680 473142
rect 526628 473078 526680 473084
rect 525248 473068 525300 473074
rect 525248 473010 525300 473016
rect 523866 472696 523922 472705
rect 523866 472631 523922 472640
rect 528020 458969 528048 600100
rect 528006 458960 528062 458969
rect 528006 458895 528062 458904
rect 529400 450673 529428 600100
rect 530780 598233 530808 600100
rect 530766 598224 530822 598233
rect 530766 598159 530822 598168
rect 532160 474201 532188 600100
rect 532146 474192 532202 474201
rect 532146 474127 532202 474136
rect 533540 467265 533568 600100
rect 533526 467256 533582 467265
rect 533526 467191 533582 467200
rect 534920 467129 534948 600100
rect 534906 467120 534962 467129
rect 534906 467055 534962 467064
rect 536300 453257 536328 600100
rect 536286 453248 536342 453257
rect 536286 453183 536342 453192
rect 529386 450664 529442 450673
rect 529386 450599 529442 450608
rect 537680 446593 537708 600100
rect 539060 472666 539088 600100
rect 539048 472660 539100 472666
rect 539048 472602 539100 472608
rect 537666 446584 537722 446593
rect 537666 446519 537722 446528
rect 522486 445224 522542 445233
rect 522486 445159 522542 445168
rect 516966 443728 517022 443737
rect 516966 443663 517022 443672
rect 539612 443601 539640 637735
rect 539690 633312 539746 633321
rect 539690 633247 539746 633256
rect 539598 443592 539654 443601
rect 539598 443527 539654 443536
rect 539704 440978 539732 633247
rect 539796 449313 539824 642495
rect 539966 631000 540022 631009
rect 539966 630935 540022 630944
rect 539874 627872 539930 627881
rect 539874 627807 539930 627816
rect 539782 449304 539838 449313
rect 539782 449239 539838 449248
rect 539888 441046 539916 627807
rect 539980 446729 540008 630935
rect 540058 625560 540114 625569
rect 540058 625495 540114 625504
rect 539966 446720 540022 446729
rect 539966 446655 540022 446664
rect 540072 445097 540100 625495
rect 540164 478378 540192 651199
rect 546498 649904 546554 649913
rect 546498 649839 546554 649848
rect 543738 648544 543794 648553
rect 543738 648479 543794 648488
rect 542634 640384 542690 640393
rect 542634 640319 542690 640328
rect 540978 639024 541034 639033
rect 540978 638959 541034 638968
rect 540152 478372 540204 478378
rect 540152 478314 540204 478320
rect 540058 445088 540114 445097
rect 540058 445023 540114 445032
rect 539876 441040 539928 441046
rect 539876 440982 539928 440988
rect 539692 440972 539744 440978
rect 539692 440914 539744 440920
rect 540992 440910 541020 638959
rect 541070 622704 541126 622713
rect 541070 622639 541126 622648
rect 541084 442338 541112 622639
rect 541162 621344 541218 621353
rect 541162 621279 541218 621288
rect 541176 473210 541204 621279
rect 542450 615904 542506 615913
rect 542450 615839 542506 615848
rect 542358 613184 542414 613193
rect 542358 613119 542414 613128
rect 541164 473204 541216 473210
rect 541164 473146 541216 473152
rect 542372 446457 542400 613119
rect 542464 449177 542492 615839
rect 542542 610464 542598 610473
rect 542542 610399 542598 610408
rect 542450 449168 542506 449177
rect 542450 449103 542506 449112
rect 542358 446448 542414 446457
rect 542358 446383 542414 446392
rect 542556 444961 542584 610399
rect 542648 475454 542676 640319
rect 542726 634944 542782 634953
rect 542726 634879 542782 634888
rect 542740 476066 542768 634879
rect 543002 632224 543058 632233
rect 543002 632159 543058 632168
rect 542910 614544 542966 614553
rect 542910 614479 542966 614488
rect 542818 609104 542874 609113
rect 542818 609039 542874 609048
rect 542728 476060 542780 476066
rect 542728 476002 542780 476008
rect 542636 475448 542688 475454
rect 542636 475390 542688 475396
rect 542832 451897 542860 609039
rect 542924 458833 542952 614479
rect 543016 478310 543044 632159
rect 543094 629504 543150 629513
rect 543094 629439 543150 629448
rect 543108 479641 543136 629439
rect 543186 611824 543242 611833
rect 543186 611759 543242 611768
rect 543094 479632 543150 479641
rect 543094 479567 543150 479576
rect 543004 478304 543056 478310
rect 543004 478246 543056 478252
rect 543200 471209 543228 611759
rect 543186 471200 543242 471209
rect 543186 471135 543242 471144
rect 543752 469849 543780 648479
rect 545118 647184 545174 647193
rect 545118 647119 545174 647128
rect 543830 645824 543886 645833
rect 543830 645759 543886 645768
rect 543738 469840 543794 469849
rect 543738 469775 543794 469784
rect 543844 469713 543872 645759
rect 543922 641744 543978 641753
rect 543922 641679 543978 641688
rect 543936 470393 543964 641679
rect 544106 624064 544162 624073
rect 544106 623999 544162 624008
rect 544014 619984 544070 619993
rect 544014 619919 544070 619928
rect 544028 473278 544056 619919
rect 544120 478854 544148 623999
rect 544198 617264 544254 617273
rect 544198 617199 544254 617208
rect 544108 478848 544160 478854
rect 544108 478790 544160 478796
rect 544212 473346 544240 617199
rect 544200 473340 544252 473346
rect 544200 473282 544252 473288
rect 544016 473272 544068 473278
rect 544016 473214 544068 473220
rect 543922 470384 543978 470393
rect 543922 470319 543978 470328
rect 545132 470121 545160 647119
rect 545210 644464 545266 644473
rect 545210 644399 545266 644408
rect 545224 470529 545252 644399
rect 545302 626784 545358 626793
rect 545302 626719 545358 626728
rect 545210 470520 545266 470529
rect 545210 470455 545266 470464
rect 545316 470257 545344 626719
rect 545302 470248 545358 470257
rect 545302 470183 545358 470192
rect 545118 470112 545174 470121
rect 545118 470047 545174 470056
rect 546512 469985 546540 649839
rect 546498 469976 546554 469985
rect 546498 469911 546554 469920
rect 543830 469704 543886 469713
rect 543830 469639 543886 469648
rect 542910 458824 542966 458833
rect 542910 458759 542966 458768
rect 542818 451888 542874 451897
rect 542818 451823 542874 451832
rect 542542 444952 542598 444961
rect 542542 444887 542598 444896
rect 541072 442332 541124 442338
rect 541072 442274 541124 442280
rect 540980 440904 541032 440910
rect 540980 440846 541032 440852
rect 577516 405686 577544 655658
rect 577596 643136 577648 643142
rect 577596 643078 577648 643084
rect 577608 475386 577636 643078
rect 577596 475380 577648 475386
rect 577596 475322 577648 475328
rect 580276 465769 580304 697167
rect 580448 657416 580500 657422
rect 580448 657358 580500 657364
rect 580356 655648 580408 655654
rect 580356 655590 580408 655596
rect 580262 465760 580318 465769
rect 580262 465695 580318 465704
rect 580368 458153 580396 655590
rect 580460 511329 580488 657358
rect 580538 656976 580594 656985
rect 580538 656911 580594 656920
rect 580552 617545 580580 656911
rect 580632 655784 580684 655790
rect 580632 655726 580684 655732
rect 580538 617536 580594 617545
rect 580538 617471 580594 617480
rect 580538 591016 580594 591025
rect 580538 590951 580594 590960
rect 580446 511320 580502 511329
rect 580446 511255 580502 511264
rect 580552 478242 580580 590951
rect 580644 564369 580672 655726
rect 580722 644056 580778 644065
rect 580722 643991 580778 644000
rect 580736 643142 580764 643991
rect 580724 643136 580776 643142
rect 580724 643078 580776 643084
rect 580630 564360 580686 564369
rect 580630 564295 580686 564304
rect 580630 537840 580686 537849
rect 580630 537775 580686 537784
rect 580540 478236 580592 478242
rect 580540 478178 580592 478184
rect 580644 478174 580672 537775
rect 580632 478168 580684 478174
rect 580632 478110 580684 478116
rect 580354 458144 580410 458153
rect 580354 458079 580410 458088
rect 580264 439748 580316 439754
rect 580264 439690 580316 439696
rect 580276 431633 580304 439690
rect 580262 431624 580318 431633
rect 580262 431559 580318 431568
rect 577504 405680 577556 405686
rect 577504 405622 577556 405628
rect 579712 405680 579764 405686
rect 579712 405622 579764 405628
rect 579724 404977 579752 405622
rect 579710 404968 579766 404977
rect 579710 404903 579766 404912
rect 580262 378448 580318 378457
rect 580262 378383 580318 378392
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580276 240281 580304 378383
rect 580262 240272 580318 240281
rect 580262 240207 580318 240216
rect 580262 236600 580318 236609
rect 580262 236535 580318 236544
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 520738 48920 520794 48929
rect 520738 48855 520794 48864
rect 511264 46912 511316 46918
rect 511264 46854 511316 46860
rect 481730 46200 481786 46209
rect 481730 46135 481786 46144
rect 471058 3768 471114 3777
rect 471058 3703 471114 3712
rect 471072 480 471100 3703
rect 478142 3632 478198 3641
rect 478142 3567 478198 3576
rect 474554 3224 474610 3233
rect 474554 3159 474610 3168
rect 474568 480 474596 3159
rect 478156 480 478184 3567
rect 481744 480 481772 46135
rect 502982 43480 503038 43489
rect 502982 43415 503038 43424
rect 499394 14512 499450 14521
rect 499394 14447 499450 14456
rect 495898 13016 495954 13025
rect 495898 12951 495954 12960
rect 492310 11656 492366 11665
rect 492310 11591 492366 11600
rect 488814 10296 488870 10305
rect 488814 10231 488870 10240
rect 485226 8936 485282 8945
rect 485226 8871 485282 8880
rect 485240 480 485268 8871
rect 488828 480 488856 10231
rect 492324 480 492352 11591
rect 495912 480 495940 12951
rect 499408 480 499436 14447
rect 502996 480 503024 43415
rect 508502 42120 508558 42129
rect 508502 42055 508558 42064
rect 506478 15872 506534 15881
rect 506478 15807 506534 15816
rect 506492 480 506520 15807
rect 508516 4049 508544 42055
rect 512642 40624 512698 40633
rect 512642 40559 512698 40568
rect 508502 4040 508558 4049
rect 508502 3975 508558 3984
rect 510066 4040 510122 4049
rect 510066 3975 510122 3984
rect 510080 480 510108 3975
rect 512656 3505 512684 40559
rect 517150 25528 517206 25537
rect 517150 25463 517206 25472
rect 512642 3496 512698 3505
rect 512642 3431 512698 3440
rect 513562 3496 513618 3505
rect 513562 3431 513618 3440
rect 513576 480 513604 3431
rect 517164 480 517192 25463
rect 520752 480 520780 48855
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 549074 44840 549130 44849
rect 549074 44775 549130 44784
rect 524234 39264 524290 39273
rect 524234 39199 524290 39208
rect 524248 480 524276 39199
rect 531318 37904 531374 37913
rect 531318 37839 531374 37848
rect 527822 17232 527878 17241
rect 527822 17167 527878 17176
rect 527836 480 527864 17167
rect 531332 480 531360 37839
rect 534906 36544 534962 36553
rect 534906 36479 534962 36488
rect 534920 480 534948 36479
rect 538402 35184 538458 35193
rect 538402 35119 538458 35128
rect 538416 480 538444 35119
rect 541990 33824 542046 33833
rect 541990 33759 542046 33768
rect 542004 480 542032 33759
rect 545486 32464 545542 32473
rect 545486 32399 545542 32408
rect 545500 480 545528 32399
rect 549088 480 549116 44775
rect 580276 33153 580304 236535
rect 580354 235240 580410 235249
rect 580354 235175 580410 235184
rect 580368 73001 580396 235175
rect 580354 72992 580410 73001
rect 580354 72927 580410 72936
rect 580262 33144 580318 33153
rect 580262 33079 580318 33088
rect 552662 30968 552718 30977
rect 552662 30903 552718 30912
rect 552676 480 552704 30903
rect 556158 29608 556214 29617
rect 556158 29543 556214 29552
rect 556172 480 556200 29543
rect 562322 28248 562378 28257
rect 562322 28183 562378 28192
rect 559746 18592 559802 18601
rect 559746 18527 559802 18536
rect 559760 480 559788 18527
rect 562336 3505 562364 28183
rect 566830 26888 566886 26897
rect 566830 26823 566886 26832
rect 562322 3496 562378 3505
rect 562322 3431 562378 3440
rect 563242 3496 563298 3505
rect 563242 3431 563298 3440
rect 563256 480 563284 3431
rect 566844 480 566872 26823
rect 570326 24168 570382 24177
rect 570326 24103 570382 24112
rect 570340 480 570368 24103
rect 573914 22672 573970 22681
rect 573914 22607 573970 22616
rect 573928 480 573956 22607
rect 576122 19952 576178 19961
rect 576122 19887 576178 19896
rect 576136 4049 576164 19887
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 576122 4040 576178 4049
rect 576122 3975 576178 3984
rect 577410 4040 577466 4049
rect 577410 3975 577466 3984
rect 577424 480 577452 3975
rect 583392 3460 583444 3466
rect 583392 3402 583444 3408
rect 582194 3360 582250 3369
rect 582194 3295 582250 3304
rect 581000 2848 581052 2854
rect 581000 2790 581052 2796
rect 581012 480 581040 2790
rect 582208 480 582236 3295
rect 583404 480 583432 3402
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 4066 553424 4122 553480
rect 3422 527856 3478 527912
rect 3974 502288 4030 502344
rect 3422 475632 3478 475688
rect 3974 474000 4030 474056
rect 4066 453328 4122 453384
rect 3422 423580 3424 423600
rect 3424 423580 3476 423600
rect 3476 423580 3478 423600
rect 3422 423544 3478 423580
rect 3422 371320 3478 371376
rect 24306 700440 24362 700496
rect 60002 700440 60058 700496
rect 40498 700304 40554 700360
rect 52642 632168 52698 632224
rect 48134 442448 48190 442504
rect 8114 364928 8170 364984
rect 5262 349152 5318 349208
rect 3422 319232 3478 319288
rect 3422 267144 3478 267200
rect 3422 214920 3478 214976
rect 3422 162832 3478 162888
rect 3422 110608 3478 110664
rect 4066 94424 4122 94480
rect 3422 71576 3478 71632
rect 570 51720 626 51776
rect 3422 32408 3478 32464
rect 2870 18808 2926 18864
rect 1674 3984 1730 4040
rect 6458 348064 6514 348120
rect 8758 95784 8814 95840
rect 7562 40840 7618 40896
rect 7654 4936 7710 4992
rect 7562 3984 7618 4040
rect 14738 235320 14794 235376
rect 12346 6160 12402 6216
rect 9954 3304 10010 3360
rect 13542 3576 13598 3632
rect 18234 269728 18290 269784
rect 17038 237496 17094 237552
rect 23018 268368 23074 268424
rect 21822 237360 21878 237416
rect 19430 2896 19486 2952
rect 31298 264152 31354 264208
rect 30102 238040 30158 238096
rect 26514 237904 26570 237960
rect 24214 225528 24270 225584
rect 25502 218592 25558 218648
rect 25502 3304 25558 3360
rect 27710 102720 27766 102776
rect 28906 3440 28962 3496
rect 34794 244840 34850 244896
rect 33598 238176 33654 238232
rect 32402 203496 32458 203552
rect 32402 3440 32458 3496
rect 32402 2760 32458 2816
rect 35990 238720 36046 238776
rect 37186 238312 37242 238368
rect 40682 238448 40738 238504
rect 39578 233824 39634 233880
rect 38382 104080 38438 104136
rect 43074 228248 43130 228304
rect 41878 105440 41934 105496
rect 50618 367648 50674 367704
rect 48226 340040 48282 340096
rect 48134 324944 48190 325000
rect 48226 295024 48282 295080
rect 44270 238584 44326 238640
rect 44178 237496 44234 237552
rect 46662 174528 46718 174584
rect 45466 106800 45522 106856
rect 48042 81640 48098 81696
rect 47582 63960 47638 64016
rect 47490 57160 47546 57216
rect 47950 62600 48006 62656
rect 47858 61240 47914 61296
rect 47766 59880 47822 59936
rect 47674 58520 47730 58576
rect 47674 28192 47730 28248
rect 47766 26832 47822 26888
rect 47858 24112 47914 24168
rect 48134 80280 48190 80336
rect 69938 633120 69994 633176
rect 69846 632848 69902 632904
rect 64786 632576 64842 632632
rect 60646 632032 60702 632088
rect 60554 579944 60610 580000
rect 60554 579536 60610 579592
rect 60002 444080 60058 444136
rect 62026 631488 62082 631544
rect 61934 629720 61990 629776
rect 61842 629584 61898 629640
rect 60738 527196 60794 527232
rect 60738 527176 60740 527196
rect 60740 527176 60792 527196
rect 60792 527176 60794 527196
rect 61750 527176 61806 527232
rect 60646 343032 60702 343088
rect 60554 342896 60610 342952
rect 61750 343576 61806 343632
rect 63406 631216 63462 631272
rect 63222 630264 63278 630320
rect 63130 630128 63186 630184
rect 62026 344120 62082 344176
rect 61934 343168 61990 343224
rect 64694 629856 64750 629912
rect 64602 629448 64658 629504
rect 63130 342624 63186 342680
rect 64694 343440 64750 343496
rect 66074 632440 66130 632496
rect 65798 492632 65854 492688
rect 64786 342760 64842 342816
rect 65982 629312 66038 629368
rect 65982 478080 66038 478136
rect 66166 631352 66222 631408
rect 69202 630808 69258 630864
rect 68926 630264 68982 630320
rect 67362 629992 67418 630048
rect 66902 629312 66958 629368
rect 66074 477808 66130 477864
rect 66902 527176 66958 527232
rect 67454 629584 67510 629640
rect 68282 629584 68338 629640
rect 67546 629448 67602 629504
rect 67454 540912 67510 540968
rect 67362 478624 67418 478680
rect 67454 344528 67510 344584
rect 66166 343576 66222 343632
rect 66074 343304 66130 343360
rect 67454 342080 67510 342136
rect 68742 604424 68798 604480
rect 68650 601024 68706 601080
rect 68282 579536 68338 579592
rect 68098 531256 68154 531312
rect 67914 522960 67970 523016
rect 68466 525816 68522 525872
rect 68190 517520 68246 517576
rect 68282 507864 68338 507920
rect 68190 479440 68246 479496
rect 68558 500792 68614 500848
rect 68282 468424 68338 468480
rect 68650 476720 68706 476776
rect 68834 513984 68890 514040
rect 68742 475360 68798 475416
rect 68558 446392 68614 446448
rect 68926 482976 68982 483032
rect 68834 351056 68890 351112
rect 68926 340720 68982 340776
rect 69570 571240 69626 571296
rect 69754 487328 69810 487384
rect 69754 478488 69810 478544
rect 69846 478352 69902 478408
rect 70030 632712 70086 632768
rect 69938 478216 69994 478272
rect 86222 700304 86278 700360
rect 89166 700304 89222 700360
rect 79782 632168 79838 632224
rect 72974 631488 73030 631544
rect 70214 630944 70270 631000
rect 70122 496304 70178 496360
rect 70030 477536 70086 477592
rect 68926 340040 68982 340096
rect 69570 340176 69626 340232
rect 70582 630672 70638 630728
rect 70306 342080 70362 342136
rect 70214 341944 70270 342000
rect 70490 341808 70546 341864
rect 70490 341400 70546 341456
rect 70122 340040 70178 340096
rect 86222 632304 86278 632360
rect 104070 634072 104126 634128
rect 88246 633120 88302 633176
rect 86866 632168 86922 632224
rect 87602 632168 87658 632224
rect 86222 631352 86278 631408
rect 87602 631216 87658 631272
rect 218978 700848 219034 700904
rect 170310 700712 170366 700768
rect 189722 700712 189778 700768
rect 202786 700712 202842 700768
rect 154118 700576 154174 700632
rect 137834 700440 137890 700496
rect 134430 657872 134486 657928
rect 129002 655560 129058 655616
rect 122286 653520 122342 653576
rect 116214 653384 116270 653440
rect 105450 633256 105506 633312
rect 110142 630944 110198 631000
rect 183006 657464 183062 657520
rect 140042 656512 140098 656568
rect 152462 655832 152518 655888
rect 146942 655696 146998 655752
rect 140134 630808 140190 630864
rect 140502 630808 140558 630864
rect 159362 654744 159418 654800
rect 152646 632712 152702 632768
rect 146942 630672 146998 630728
rect 170862 652024 170918 652080
rect 164790 634208 164846 634264
rect 158718 632576 158774 632632
rect 159362 632576 159418 632632
rect 164790 632440 164846 632496
rect 176934 635432 176990 635488
rect 170862 630128 170918 630184
rect 176658 629992 176714 630048
rect 267646 700984 267702 701040
rect 292854 700984 292910 701040
rect 292762 700712 292818 700768
rect 292578 700576 292634 700632
rect 283838 700168 283894 700224
rect 235170 657464 235226 657520
rect 189078 657056 189134 657112
rect 189722 657056 189778 657112
rect 183006 629856 183062 629912
rect 225510 656376 225566 656432
rect 213182 656240 213238 656296
rect 200762 656104 200818 656160
rect 195242 655968 195298 656024
rect 207662 654472 207718 654528
rect 195242 633256 195298 633312
rect 200854 632304 200910 632360
rect 201222 632304 201278 632360
rect 207662 632168 207718 632224
rect 224958 655560 225014 655616
rect 219438 654608 219494 654664
rect 213182 632032 213238 632088
rect 189078 629720 189134 629776
rect 219438 629584 219494 629640
rect 225510 629448 225566 629504
rect 262126 653656 262182 653712
rect 249798 649168 249854 649224
rect 268014 632168 268070 632224
rect 289818 636792 289874 636848
rect 289818 633256 289874 633312
rect 262126 632032 262182 632088
rect 249798 629584 249854 629640
rect 291290 605920 291346 605976
rect 289910 564440 289966 564496
rect 289818 552336 289874 552392
rect 289358 507864 289414 507920
rect 289542 499704 289598 499760
rect 289450 491272 289506 491328
rect 288990 480256 289046 480312
rect 72514 477536 72570 477592
rect 70674 341400 70730 341456
rect 70674 340992 70730 341048
rect 79138 478624 79194 478680
rect 75826 477808 75882 477864
rect 73710 389408 73766 389464
rect 73710 342760 73766 342816
rect 77298 342624 77354 342680
rect 84106 478352 84162 478408
rect 79782 389952 79838 390008
rect 80334 343440 80390 343496
rect 81990 343168 82046 343224
rect 91926 391040 91982 391096
rect 85854 390496 85910 390552
rect 85578 343304 85634 343360
rect 88614 343032 88670 343088
rect 90270 342896 90326 342952
rect 99378 478216 99434 478272
rect 102322 478216 102378 478272
rect 99010 478080 99066 478136
rect 97998 391584 98054 391640
rect 104162 478352 104218 478408
rect 104070 392128 104126 392184
rect 105542 477944 105598 478000
rect 108302 477808 108358 477864
rect 106922 477672 106978 477728
rect 110142 454688 110198 454744
rect 112994 440680 113050 440736
rect 111062 388320 111118 388376
rect 54574 278704 54630 278760
rect 56230 278568 56286 278624
rect 52918 277344 52974 277400
rect 57702 277072 57758 277128
rect 59266 276936 59322 276992
rect 61198 276800 61254 276856
rect 64510 277888 64566 277944
rect 69156 280064 69212 280120
rect 71134 279656 71190 279712
rect 67546 279112 67602 279168
rect 74124 280064 74180 280120
rect 75826 279248 75882 279304
rect 72790 278976 72846 279032
rect 78954 279928 79010 279984
rect 79414 279520 79470 279576
rect 78586 279112 78642 279168
rect 80748 279792 80804 279848
rect 81438 279656 81494 279712
rect 83002 279656 83058 279712
rect 83094 279384 83150 279440
rect 83370 279384 83426 279440
rect 80058 278976 80114 279032
rect 77758 278840 77814 278896
rect 84106 278024 84162 278080
rect 86038 277752 86094 277808
rect 89718 278588 89774 278624
rect 89718 278568 89720 278588
rect 89720 278568 89772 278588
rect 89772 278568 89774 278588
rect 89350 278432 89406 278488
rect 91098 278704 91154 278760
rect 92386 278704 92442 278760
rect 91006 278296 91062 278352
rect 96526 280064 96582 280120
rect 95974 279112 96030 279168
rect 94318 278160 94374 278216
rect 97906 278024 97962 278080
rect 95146 277888 95202 277944
rect 97630 277888 97686 277944
rect 100620 280064 100676 280120
rect 99378 279520 99434 279576
rect 102138 278432 102194 278488
rect 99286 278024 99342 278080
rect 98642 277752 98698 277808
rect 87694 277616 87750 277672
rect 104254 278432 104310 278488
rect 107382 278704 107438 278760
rect 107566 278704 107622 278760
rect 106186 278332 106188 278352
rect 106188 278332 106240 278352
rect 106240 278332 106242 278352
rect 106186 278296 106242 278332
rect 111246 386688 111302 386744
rect 111062 278704 111118 278760
rect 108946 278568 109002 278624
rect 108302 278160 108358 278216
rect 105910 277752 105966 277808
rect 104806 277616 104862 277672
rect 111430 385600 111486 385656
rect 111338 379072 111394 379128
rect 111338 279792 111394 279848
rect 112626 384512 112682 384568
rect 112626 279112 112682 279168
rect 113086 439048 113142 439104
rect 112994 339360 113050 339416
rect 116214 431160 116270 431216
rect 123482 479440 123538 479496
rect 122286 393760 122342 393816
rect 116582 387776 116638 387832
rect 115202 386144 115258 386200
rect 114006 380160 114062 380216
rect 113822 379616 113878 379672
rect 113086 322904 113142 322960
rect 113822 279928 113878 279984
rect 115202 280064 115258 280120
rect 114006 279656 114062 279712
rect 116398 318008 116454 318064
rect 111430 278024 111486 278080
rect 102598 277480 102654 277536
rect 111246 277480 111302 277536
rect 66166 277208 66222 277264
rect 62854 276664 62910 276720
rect 98642 272584 98698 272640
rect 87970 224168 88026 224224
rect 85670 204856 85726 204912
rect 52918 87760 52974 87816
rect 50986 85856 51042 85912
rect 63866 87624 63922 87680
rect 59266 87488 59322 87544
rect 57610 87216 57666 87272
rect 54666 87080 54722 87136
rect 56506 86128 56562 86184
rect 62026 87352 62082 87408
rect 60646 85720 60702 85776
rect 84934 87488 84990 87544
rect 65614 86944 65670 87000
rect 68650 85992 68706 86048
rect 66994 85584 67050 85640
rect 82312 84904 82368 84960
rect 77620 84768 77676 84824
rect 71364 84632 71420 84688
rect 79184 84496 79240 84552
rect 84290 83408 84346 83464
rect 84934 80688 84990 80744
rect 49330 78920 49386 78976
rect 49238 69400 49294 69456
rect 49054 68040 49110 68096
rect 48226 51448 48282 51504
rect 48134 49000 48190 49056
rect 49146 54440 49202 54496
rect 49054 48864 49110 48920
rect 48042 42200 48098 42256
rect 49606 77560 49662 77616
rect 49514 74840 49570 74896
rect 49422 72120 49478 72176
rect 49330 44784 49386 44840
rect 49238 39208 49294 39264
rect 49422 37848 49478 37904
rect 49514 35128 49570 35184
rect 50250 75928 50306 75984
rect 50158 70352 50214 70408
rect 50066 52536 50122 52592
rect 50066 43560 50122 43616
rect 49606 32408 49662 32464
rect 49146 30912 49202 30968
rect 47950 22616 48006 22672
rect 47582 19896 47638 19952
rect 47490 18536 47546 18592
rect 50434 73208 50490 73264
rect 50342 66272 50398 66328
rect 50250 33768 50306 33824
rect 50618 65048 50674 65104
rect 50526 55528 50582 55584
rect 50434 36488 50490 36544
rect 84658 53216 84714 53272
rect 83278 50496 83334 50552
rect 50986 47776 51042 47832
rect 52366 47640 52422 47696
rect 53746 47504 53802 47560
rect 50618 46280 50674 46336
rect 51354 37984 51410 38040
rect 50526 29552 50582 29608
rect 50342 25472 50398 25528
rect 50158 17176 50214 17232
rect 48962 7792 49018 7848
rect 47858 6296 47914 6352
rect 50158 3440 50214 3496
rect 51722 36624 51778 36680
rect 52550 27104 52606 27160
rect 51722 3440 51778 3496
rect 53746 26968 53802 27024
rect 54942 6432 54998 6488
rect 56506 46144 56562 46200
rect 56046 29824 56102 29880
rect 55034 4800 55090 4856
rect 59634 28464 59690 28520
rect 59174 10240 59230 10296
rect 58622 8880 58678 8936
rect 58438 6568 58494 6624
rect 57242 3440 57298 3496
rect 63222 31048 63278 31104
rect 61934 12960 61990 13016
rect 60554 11600 60610 11656
rect 62026 6704 62082 6760
rect 60830 3304 60886 3360
rect 64694 43424 64750 43480
rect 65522 24248 65578 24304
rect 64326 18672 64382 18728
rect 63314 14456 63370 14512
rect 67454 42064 67510 42120
rect 68834 40568 68890 40624
rect 66718 32680 66774 32736
rect 66074 15816 66130 15872
rect 70306 34040 70362 34096
rect 70214 21392 70270 21448
rect 69110 20032 69166 20088
rect 67914 3712 67970 3768
rect 71502 32544 71558 32600
rect 74446 46960 74502 47016
rect 75182 46960 75238 47016
rect 73802 35264 73858 35320
rect 72974 21256 73030 21312
rect 71594 10376 71650 10432
rect 72606 6840 72662 6896
rect 74998 28328 75054 28384
rect 77390 36760 77446 36816
rect 77114 14592 77170 14648
rect 76562 13096 76618 13152
rect 75182 11736 75238 11792
rect 76194 6024 76250 6080
rect 79690 25608 79746 25664
rect 79322 15952 79378 16008
rect 78586 7656 78642 7712
rect 82726 47912 82782 47968
rect 81254 40704 81310 40760
rect 80886 33904 80942 33960
rect 79874 17312 79930 17368
rect 82082 29688 82138 29744
rect 83462 47912 83518 47968
rect 84014 39344 84070 39400
rect 83462 22752 83518 22808
rect 86866 91704 86922 91760
rect 86222 87760 86278 87816
rect 86406 87216 86462 87272
rect 86406 53080 86462 53136
rect 86222 51720 86278 51776
rect 87602 90344 87658 90400
rect 87878 87624 87934 87680
rect 87694 87080 87750 87136
rect 86958 52536 87014 52592
rect 87602 52536 87658 52592
rect 87878 54576 87934 54632
rect 87694 50224 87750 50280
rect 86958 40840 87014 40896
rect 96250 221448 96306 221504
rect 92754 220088 92810 220144
rect 91742 214512 91798 214568
rect 90362 213152 90418 213208
rect 89166 88984 89222 89040
rect 91558 97144 91614 97200
rect 90638 87352 90694 87408
rect 90454 86944 90510 87000
rect 90638 69536 90694 69592
rect 90454 9016 90510 9072
rect 91742 3440 91798 3496
rect 93950 211792 94006 211848
rect 95146 98640 95202 98696
rect 97446 210296 97502 210352
rect 105726 243480 105782 243536
rect 101402 239536 101458 239592
rect 99838 229744 99894 229800
rect 101034 177248 101090 177304
rect 103334 226888 103390 226944
rect 102230 100000 102286 100056
rect 101402 3712 101458 3768
rect 104530 208936 104586 208992
rect 114006 236680 114062 236736
rect 106922 233960 106978 234016
rect 110510 222808 110566 222864
rect 108118 178608 108174 178664
rect 109314 5072 109370 5128
rect 112810 101360 112866 101416
rect 111614 93064 111670 93120
rect 115202 207576 115258 207632
rect 119434 387232 119490 387288
rect 117962 385056 118018 385112
rect 119342 331200 119398 331256
rect 117962 277888 118018 277944
rect 116582 277752 116638 277808
rect 118790 3848 118846 3904
rect 117594 3440 117650 3496
rect 120722 378528 120778 378584
rect 122102 373632 122158 373688
rect 120722 279248 120778 279304
rect 119434 278432 119490 278488
rect 123482 284960 123538 285016
rect 123666 373088 123722 373144
rect 134430 394848 134486 394904
rect 128358 394304 128414 394360
rect 126334 388864 126390 388920
rect 127714 372544 127770 372600
rect 126334 278568 126390 278624
rect 130382 372000 130438 372056
rect 134522 370368 134578 370424
rect 140502 395392 140558 395448
rect 140042 374720 140098 374776
rect 134522 277344 134578 277400
rect 142802 339360 142858 339416
rect 140042 277208 140098 277264
rect 130382 277072 130438 277128
rect 127714 276936 127770 276992
rect 123666 276800 123722 276856
rect 122102 276664 122158 276720
rect 123482 265512 123538 265568
rect 122286 237768 122342 237824
rect 121458 237360 121514 237416
rect 121090 232464 121146 232520
rect 119894 3712 119950 3768
rect 119342 3576 119398 3632
rect 141238 235456 141294 235512
rect 126978 232600 127034 232656
rect 126242 206216 126298 206272
rect 126242 3848 126298 3904
rect 124678 3576 124734 3632
rect 130566 225664 130622 225720
rect 134154 220224 134210 220280
rect 137650 200640 137706 200696
rect 151174 474000 151230 474056
rect 146574 395936 146630 395992
rect 146942 345344 146998 345400
rect 144734 197920 144790 197976
rect 142802 34040 142858 34096
rect 151082 336640 151138 336696
rect 148322 239264 148378 239320
rect 146942 5072 146998 5128
rect 155222 468424 155278 468480
rect 152646 396480 152702 396536
rect 151174 301824 151230 301880
rect 164790 464344 164846 464400
rect 189078 474000 189134 474056
rect 199474 446392 199530 446448
rect 195150 400288 195206 400344
rect 183006 399200 183062 399256
rect 176934 398656 176990 398712
rect 170862 398112 170918 398168
rect 158718 397024 158774 397080
rect 159362 349696 159418 349752
rect 155222 275712 155278 275768
rect 158902 238992 158958 239048
rect 155406 231104 155462 231160
rect 151818 196560 151874 196616
rect 151082 27104 151138 27160
rect 163502 346976 163558 347032
rect 162490 236816 162546 236872
rect 159362 18808 159418 18864
rect 174542 343168 174598 343224
rect 173162 239128 173218 239184
rect 166078 228384 166134 228440
rect 163502 3712 163558 3768
rect 169574 3712 169630 3768
rect 175922 338816 175978 338872
rect 174542 98640 174598 98696
rect 178682 337728 178738 337784
rect 176658 239400 176714 239456
rect 175922 32680 175978 32736
rect 188342 337184 188398 337240
rect 184202 335552 184258 335608
rect 180246 238856 180302 238912
rect 179418 238720 179474 238776
rect 178682 28464 178738 28520
rect 183742 235592 183798 235648
rect 186962 333920 187018 333976
rect 186962 244840 187018 244896
rect 186318 239536 186374 239592
rect 187330 238720 187386 238776
rect 184202 106800 184258 106856
rect 191102 335008 191158 335064
rect 190826 229880 190882 229936
rect 188342 29824 188398 29880
rect 199382 345888 199438 345944
rect 195242 340448 195298 340504
rect 194414 231240 194470 231296
rect 191102 105440 191158 105496
rect 198002 334464 198058 334520
rect 197910 234096 197966 234152
rect 195242 36760 195298 36816
rect 198002 104080 198058 104136
rect 211802 431160 211858 431216
rect 207294 401376 207350 401432
rect 201222 400832 201278 400888
rect 214654 475360 214710 475416
rect 213366 401920 213422 401976
rect 211802 393216 211858 393272
rect 210422 348608 210478 348664
rect 202142 344800 202198 344856
rect 199474 275168 199530 275224
rect 203522 338272 203578 338328
rect 202142 243480 202198 243536
rect 201498 236952 201554 237008
rect 199382 101360 199438 101416
rect 206282 336096 206338 336152
rect 205086 222944 205142 223000
rect 203522 31048 203578 31104
rect 209042 332832 209098 332888
rect 208582 232736 208638 232792
rect 206282 7792 206338 7848
rect 209042 102720 209098 102776
rect 211802 342624 211858 342680
rect 212446 239264 212502 239320
rect 212722 239264 212778 239320
rect 211802 97144 211858 97200
rect 210422 94424 210478 94480
rect 214562 330112 214618 330168
rect 215942 474000 215998 474056
rect 218702 442992 218758 443048
rect 215942 399744 215998 399800
rect 214654 288224 214710 288280
rect 215666 224304 215722 224360
rect 214562 90344 214618 90400
rect 213182 53216 213238 53272
rect 216126 347520 216182 347576
rect 217322 344256 217378 344312
rect 216678 344120 216734 344176
rect 216126 265512 216182 265568
rect 215942 224168 215998 224224
rect 224774 477536 224830 477592
rect 224222 476720 224278 476776
rect 222106 469784 222162 469840
rect 222014 440816 222070 440872
rect 219438 402464 219494 402520
rect 220082 339904 220138 339960
rect 218702 305904 218758 305960
rect 219254 203632 219310 203688
rect 217322 100000 217378 100056
rect 222842 343712 222898 343768
rect 222106 327936 222162 327992
rect 222014 299376 222070 299432
rect 224866 470056 224922 470112
rect 224774 409944 224830 410000
rect 224314 332288 224370 332344
rect 224222 287680 224278 287736
rect 222842 272584 222898 272640
rect 231214 478760 231270 478816
rect 228454 478624 228510 478680
rect 227718 477536 227774 477592
rect 227626 475632 227682 475688
rect 227534 474952 227590 475008
rect 227442 473048 227498 473104
rect 227350 472912 227406 472968
rect 227258 472232 227314 472288
rect 226062 470328 226118 470384
rect 225970 469920 226026 469976
rect 225510 403008 225566 403064
rect 225602 344936 225658 344992
rect 225418 344392 225474 344448
rect 224866 327392 224922 327448
rect 225418 283328 225474 283384
rect 225786 343984 225842 344040
rect 225694 333376 225750 333432
rect 225602 271904 225658 271960
rect 224314 268368 224370 268424
rect 225786 283872 225842 283928
rect 225970 328480 226026 328536
rect 226246 470192 226302 470248
rect 226154 442176 226210 442232
rect 226062 325216 226118 325272
rect 226982 454688 227038 454744
rect 226890 444080 226946 444136
rect 226890 443808 226946 443864
rect 227166 440292 227222 440328
rect 227166 440272 227168 440292
rect 227168 440272 227220 440292
rect 227220 440272 227222 440292
rect 226982 392672 227038 392728
rect 227258 363840 227314 363896
rect 227350 357856 227406 357912
rect 227534 356768 227590 356824
rect 227442 355136 227498 355192
rect 227074 351056 227130 351112
rect 226982 330656 227038 330712
rect 226246 319232 226302 319288
rect 226154 295296 226210 295352
rect 225694 264152 225750 264208
rect 222750 230016 222806 230072
rect 220082 35264 220138 35320
rect 226338 221584 226394 221640
rect 227166 346432 227222 346488
rect 227166 318008 227222 318064
rect 228178 475224 228234 475280
rect 227626 299104 227682 299160
rect 228362 470464 228418 470520
rect 228270 442720 228326 442776
rect 228362 406000 228418 406056
rect 228822 475088 228878 475144
rect 228638 472640 228694 472696
rect 228546 472096 228602 472152
rect 228454 405728 228510 405784
rect 228546 364384 228602 364440
rect 228730 439184 228786 439240
rect 228638 363296 228694 363352
rect 228454 344528 228510 344584
rect 228178 297472 228234 297528
rect 227074 276256 227130 276312
rect 226982 95784 227038 95840
rect 228454 281696 228510 281752
rect 230386 475360 230442 475416
rect 230202 474816 230258 474872
rect 229742 472504 229798 472560
rect 229006 442040 229062 442096
rect 229650 442040 229706 442096
rect 229650 441632 229706 441688
rect 229006 440816 229062 440872
rect 229650 440680 229706 440736
rect 228914 440272 228970 440328
rect 228914 440136 228970 440192
rect 228822 357312 228878 357368
rect 228730 331336 228786 331392
rect 229650 440000 229706 440056
rect 229374 439592 229430 439648
rect 229650 439592 229706 439648
rect 229006 439320 229062 439376
rect 229650 439048 229706 439104
rect 230110 472776 230166 472832
rect 230018 439884 230074 439920
rect 230018 439864 230020 439884
rect 230020 439864 230072 439884
rect 230072 439864 230074 439884
rect 230110 361664 230166 361720
rect 230386 472368 230442 472424
rect 230294 471960 230350 472016
rect 230202 356224 230258 356280
rect 229742 340720 229798 340776
rect 230294 334056 230350 334112
rect 229834 331744 229890 331800
rect 229742 329704 229798 329760
rect 228914 304000 228970 304056
rect 231122 464344 231178 464400
rect 230478 440580 230480 440600
rect 230480 440580 230532 440600
rect 230532 440580 230534 440600
rect 230478 440544 230534 440580
rect 231030 439048 231086 439104
rect 231490 475496 231546 475552
rect 231306 474136 231362 474192
rect 231214 404640 231270 404696
rect 231122 397568 231178 397624
rect 231398 440272 231454 440328
rect 231306 366560 231362 366616
rect 231214 364928 231270 364984
rect 230938 341944 230994 342000
rect 230386 296928 230442 296984
rect 231122 341264 231178 341320
rect 230938 278976 230994 279032
rect 231306 341808 231362 341864
rect 231214 301280 231270 301336
rect 231122 278432 231178 278488
rect 234526 479576 234582 479632
rect 231766 477808 231822 477864
rect 233146 477672 233202 477728
rect 231858 475360 231914 475416
rect 232870 475360 232926 475416
rect 231582 403552 231638 403608
rect 231582 369824 231638 369880
rect 231582 367648 231638 367704
rect 231490 350240 231546 350296
rect 231490 341128 231546 341184
rect 231398 324400 231454 324456
rect 231674 329024 231730 329080
rect 232686 440272 232742 440328
rect 232778 369280 232834 369336
rect 232962 469648 233018 469704
rect 232870 355680 232926 355736
rect 232962 326848 233018 326904
rect 231766 320864 231822 320920
rect 233882 475224 233938 475280
rect 234250 475224 234306 475280
rect 233146 465704 233202 465760
rect 233054 313248 233110 313304
rect 234158 451832 234214 451888
rect 233790 449112 233846 449168
rect 233882 446392 233938 446448
rect 233974 444896 234030 444952
rect 233974 441632 234030 441688
rect 233882 313792 233938 313848
rect 234066 314880 234122 314936
rect 233974 312704 234030 312760
rect 234250 322496 234306 322552
rect 234434 471144 234490 471200
rect 234342 321408 234398 321464
rect 235446 458904 235502 458960
rect 235078 453192 235134 453248
rect 234986 448160 235042 448216
rect 234894 440136 234950 440192
rect 234894 439320 234950 439376
rect 235170 450608 235226 450664
rect 235078 368192 235134 368248
rect 235354 445304 235410 445360
rect 235262 443536 235318 443592
rect 235170 365472 235226 365528
rect 235538 446800 235594 446856
rect 235446 364928 235502 364984
rect 235354 354592 235410 354648
rect 235262 353504 235318 353560
rect 237102 471280 237158 471336
rect 235814 467200 235870 467256
rect 235722 467064 235778 467120
rect 235630 444080 235686 444136
rect 235722 367648 235778 367704
rect 235906 465840 235962 465896
rect 235814 367104 235870 367160
rect 235538 352960 235594 353016
rect 234986 351872 235042 351928
rect 236918 464344 236974 464400
rect 236826 460128 236882 460184
rect 236734 448024 236790 448080
rect 236642 447752 236698 447808
rect 236458 445168 236514 445224
rect 236550 443672 236606 443728
rect 236458 362752 236514 362808
rect 236550 360576 236606 360632
rect 236642 360032 236698 360088
rect 236826 359488 236882 359544
rect 237010 462848 237066 462904
rect 236918 358400 236974 358456
rect 236734 354048 236790 354104
rect 235906 351328 235962 351384
rect 237194 468560 237250 468616
rect 237102 358944 237158 359000
rect 237286 450744 237342 450800
rect 237194 352416 237250 352472
rect 237010 350784 237066 350840
rect 234526 320320 234582 320376
rect 234434 313248 234490 313304
rect 234158 312160 234214 312216
rect 235814 340992 235870 341048
rect 235906 340856 235962 340912
rect 235814 324672 235870 324728
rect 235906 314336 235962 314392
rect 235906 307672 235962 307728
rect 233146 296384 233202 296440
rect 231490 279520 231546 279576
rect 231306 277888 231362 277944
rect 237378 443808 237434 443864
rect 237562 443808 237618 443864
rect 237562 443536 237618 443592
rect 244830 479712 244886 479768
rect 243726 478760 243782 478816
rect 241794 478488 241850 478544
rect 241426 477944 241482 478000
rect 238482 471960 238538 472016
rect 239494 454688 239550 454744
rect 239402 446936 239458 446992
rect 238574 446664 238630 446720
rect 238298 443536 238354 443592
rect 238022 443400 238078 443456
rect 237654 404096 237710 404152
rect 237378 383968 237434 384024
rect 237378 383424 237434 383480
rect 237470 382880 237526 382936
rect 237378 382356 237434 382392
rect 237378 382336 237380 382356
rect 237380 382336 237432 382356
rect 237432 382336 237434 382356
rect 237562 381792 237618 381848
rect 237378 381248 237434 381304
rect 237378 380704 237434 380760
rect 237746 377984 237802 378040
rect 237562 377440 237618 377496
rect 237378 376916 237434 376952
rect 237378 376896 237380 376916
rect 237380 376896 237432 376916
rect 237432 376896 237434 376916
rect 237562 376352 237618 376408
rect 237378 375808 237434 375864
rect 237378 375264 237434 375320
rect 237378 374176 237434 374232
rect 237378 371456 237434 371512
rect 237378 370912 237434 370968
rect 238022 366016 238078 366072
rect 237930 347656 237986 347712
rect 237562 342080 237618 342136
rect 237378 341536 237434 341592
rect 237378 340992 237434 341048
rect 237838 340176 237894 340232
rect 237378 320864 237434 320920
rect 237378 316920 237434 316976
rect 237378 300772 237380 300792
rect 237380 300772 237432 300792
rect 237432 300772 237434 300792
rect 237378 300736 237434 300772
rect 237286 298560 237342 298616
rect 237378 287136 237434 287192
rect 238022 340040 238078 340096
rect 237930 325760 237986 325816
rect 237838 286592 237894 286648
rect 237378 286048 237434 286104
rect 237378 285504 237434 285560
rect 238114 324128 238170 324184
rect 238298 323584 238354 323640
rect 238206 321952 238262 322008
rect 238390 319776 238446 319832
rect 239310 445440 239366 445496
rect 238666 445032 238722 445088
rect 238574 320864 238630 320920
rect 239126 444080 239182 444136
rect 239034 442584 239090 442640
rect 239678 449384 239734 449440
rect 239586 447888 239642 447944
rect 239494 408448 239550 408504
rect 239402 407904 239458 407960
rect 239310 407360 239366 407416
rect 239218 406816 239274 406872
rect 239034 406272 239090 406328
rect 239494 405184 239550 405240
rect 239494 401512 239550 401568
rect 240046 444216 240102 444272
rect 240046 442448 240102 442504
rect 239770 439048 239826 439104
rect 239678 362208 239734 362264
rect 239586 361120 239642 361176
rect 238666 318688 238722 318744
rect 238482 317600 238538 317656
rect 239770 300192 239826 300248
rect 243818 475768 243874 475824
rect 243542 475224 243598 475280
rect 255870 478624 255926 478680
rect 258998 478488 259054 478544
rect 249798 477944 249854 478000
rect 249890 475904 249946 475960
rect 247866 473184 247922 473240
rect 247038 472096 247094 472152
rect 246854 465976 246910 466032
rect 245842 464480 245898 464536
rect 248878 460264 248934 460320
rect 251086 475088 251142 475144
rect 257986 474272 258042 474328
rect 256054 472368 256110 472424
rect 255318 472232 255374 472288
rect 251914 471416 251970 471472
rect 250902 442448 250958 442504
rect 251086 442176 251142 442232
rect 252926 462984 252982 463040
rect 256974 467472 257030 467528
rect 254030 442720 254086 442776
rect 253938 442312 253994 442368
rect 254398 442448 254454 442504
rect 254950 442312 255006 442368
rect 260010 476856 260066 476912
rect 261022 459040 261078 459096
rect 264058 479848 264114 479904
rect 262034 478624 262090 478680
rect 261942 442584 261998 442640
rect 263046 476040 263102 476096
rect 262862 474952 262918 475008
rect 267094 478760 267150 478816
rect 265070 442720 265126 442776
rect 264978 442040 265034 442096
rect 266082 442584 266138 442640
rect 268106 479984 268162 480040
rect 268014 444080 268070 444136
rect 271234 476992 271290 477048
rect 271142 475224 271198 475280
rect 269118 474408 269174 474464
rect 270130 442856 270186 442912
rect 270406 441904 270462 441960
rect 271786 474816 271842 474872
rect 273166 471552 273222 471608
rect 271234 442856 271290 442912
rect 272154 442856 272210 442912
rect 278226 480120 278282 480176
rect 276202 477944 276258 478000
rect 275190 468696 275246 468752
rect 274086 445440 274142 445496
rect 274178 442040 274234 442096
rect 273258 441768 273314 441824
rect 279238 456184 279294 456240
rect 286230 454688 286286 454744
rect 283010 453328 283066 453384
rect 280158 446936 280214 446992
rect 280526 405728 280582 405784
rect 281906 441496 281962 441552
rect 281630 440544 281686 440600
rect 281538 440408 281594 440464
rect 281722 440000 281778 440056
rect 281630 435648 281686 435704
rect 281538 434288 281594 434344
rect 280986 416608 281042 416664
rect 282366 441360 282422 441416
rect 282274 440816 282330 440872
rect 281906 432928 281962 432984
rect 282458 440136 282514 440192
rect 282182 427488 282238 427544
rect 282090 424768 282146 424824
rect 281906 422048 281962 422104
rect 281814 420688 281870 420744
rect 281722 419328 281778 419384
rect 281630 417968 281686 418024
rect 281538 415248 281594 415304
rect 280894 413888 280950 413944
rect 280802 412528 280858 412584
rect 281906 409828 281962 409864
rect 281906 409808 281908 409828
rect 281908 409808 281960 409828
rect 281960 409808 281962 409828
rect 281906 408468 281962 408504
rect 281906 408448 281908 408468
rect 281908 408448 281960 408468
rect 281960 408448 281962 408468
rect 280710 407088 280766 407144
rect 280618 404368 280674 404424
rect 280434 403008 280490 403064
rect 280342 401648 280398 401704
rect 280250 400288 280306 400344
rect 280158 398928 280214 398984
rect 280066 397568 280122 397624
rect 282826 395664 282882 395720
rect 281814 393488 281870 393544
rect 280158 389408 280214 389464
rect 239862 299648 239918 299704
rect 280066 296928 280122 296984
rect 239862 289312 239918 289368
rect 239770 288768 239826 288824
rect 238022 284416 238078 284472
rect 237378 282240 237434 282296
rect 237378 281152 237434 281208
rect 238666 281424 238722 281480
rect 237562 280608 237618 280664
rect 237378 280100 237380 280120
rect 237380 280100 237432 280120
rect 237432 280100 237434 280120
rect 237378 280064 237434 280100
rect 235906 277344 235962 277400
rect 229834 269728 229890 269784
rect 238666 240216 238722 240272
rect 237010 239536 237066 239592
rect 235998 238992 236054 239048
rect 233422 237088 233478 237144
rect 229834 228520 229890 228576
rect 228362 33904 228418 33960
rect 237378 239400 237434 239456
rect 237470 239128 237526 239184
rect 237562 238856 237618 238912
rect 239770 236544 239826 236600
rect 280066 241848 280122 241904
rect 280066 241712 280122 241768
rect 239862 235184 239918 235240
rect 252190 238584 252246 238640
rect 250994 238448 251050 238504
rect 249798 238312 249854 238368
rect 248602 238176 248658 238232
rect 251178 238176 251234 238232
rect 247406 238040 247462 238096
rect 246210 237904 246266 237960
rect 247590 237904 247646 237960
rect 246302 69400 246358 69456
rect 242622 6160 242678 6216
rect 241426 4936 241482 4992
rect 246302 4936 246358 4992
rect 240506 3848 240562 3904
rect 244094 3984 244150 4040
rect 243542 2896 243598 2952
rect 250442 78920 250498 78976
rect 250442 50360 250498 50416
rect 254674 238040 254730 238096
rect 254582 37984 254638 38040
rect 253386 6296 253442 6352
rect 258262 239400 258318 239456
rect 258170 6704 258226 6760
rect 256974 6568 257030 6624
rect 255778 6432 255834 6488
rect 259274 238720 259330 238776
rect 259366 24248 259422 24304
rect 260562 20032 260618 20088
rect 261758 238312 261814 238368
rect 261666 6840 261722 6896
rect 264978 239264 265034 239320
rect 265346 239128 265402 239184
rect 265254 50496 265310 50552
rect 264150 25608 264206 25664
rect 262954 6024 263010 6080
rect 267738 213152 267794 213208
rect 268934 211792 268990 211848
rect 270130 210296 270186 210352
rect 272522 208936 272578 208992
rect 273718 178608 273774 178664
rect 271326 177248 271382 177304
rect 275282 207576 275338 207632
rect 278502 237768 278558 237824
rect 277306 206216 277362 206272
rect 274914 93064 274970 93120
rect 266542 91704 266598 91760
rect 275282 85992 275338 86048
rect 271142 85856 271198 85912
rect 268842 49000 268898 49056
rect 273902 54440 273958 54496
rect 278042 21392 278098 21448
rect 273902 5072 273958 5128
rect 271142 3304 271198 3360
rect 272430 3304 272486 3360
rect 271786 2760 271842 2816
rect 278042 3304 278098 3360
rect 279514 3304 279570 3360
rect 280250 383968 280306 384024
rect 280158 239128 280214 239184
rect 281722 382608 281778 382664
rect 281630 381248 281686 381304
rect 281538 379888 281594 379944
rect 280434 378528 280490 378584
rect 280342 373088 280398 373144
rect 280250 238176 280306 238232
rect 280526 367648 280582 367704
rect 280434 239536 280490 239592
rect 280618 362208 280674 362264
rect 280526 232736 280582 232792
rect 280710 358128 280766 358184
rect 280894 355408 280950 355464
rect 280802 311888 280858 311944
rect 280710 235592 280766 235648
rect 280618 231240 280674 231296
rect 280342 230016 280398 230072
rect 281446 312024 281502 312080
rect 281538 311888 281594 311944
rect 280986 299376 281042 299432
rect 281630 299376 281686 299432
rect 282826 369008 282882 369064
rect 281998 364928 282054 364984
rect 281906 360848 281962 360904
rect 281814 305088 281870 305144
rect 281722 237904 281778 237960
rect 282826 359488 282882 359544
rect 282826 356768 282882 356824
rect 282826 354048 282882 354104
rect 282826 348608 282882 348664
rect 282826 344528 282882 344584
rect 282918 315968 282974 316024
rect 282274 313248 282330 313304
rect 282182 309168 282238 309224
rect 282090 298288 282146 298344
rect 281998 236952 282054 237008
rect 281906 229880 281962 229936
rect 282366 310528 282422 310584
rect 282550 306448 282606 306504
rect 282366 241712 282422 241768
rect 282274 240896 282330 240952
rect 282274 240352 282330 240408
rect 282182 214512 282238 214568
rect 282090 203496 282146 203552
rect 281814 174528 281870 174584
rect 282826 295568 282882 295624
rect 282826 280608 282882 280664
rect 282826 273808 282882 273864
rect 282826 272448 282882 272504
rect 282550 36624 282606 36680
rect 283102 442992 283158 443048
rect 283102 411168 283158 411224
rect 283102 388048 283158 388104
rect 283010 275168 283066 275224
rect 284482 385328 284538 385384
rect 284390 374448 284446 374504
rect 284298 371728 284354 371784
rect 283286 366288 283342 366344
rect 283194 345888 283250 345944
rect 283102 238312 283158 238368
rect 283378 363568 283434 363624
rect 283470 351328 283526 351384
rect 283378 234096 283434 234152
rect 283562 349968 283618 350024
rect 283654 337728 283710 337784
rect 283562 236816 283618 236872
rect 283470 228384 283526 228440
rect 283746 336368 283802 336424
rect 283838 274624 283894 274680
rect 283746 232600 283802 232656
rect 283654 225664 283710 225720
rect 283286 222944 283342 223000
rect 283194 196560 283250 196616
rect 282918 28328 282974 28384
rect 281538 18672 281594 18728
rect 283102 5072 283158 5128
rect 280986 3984 281042 4040
rect 280802 3848 280858 3904
rect 280066 3168 280122 3224
rect 284850 377168 284906 377224
rect 284574 375808 284630 375864
rect 284482 240080 284538 240136
rect 284666 370368 284722 370424
rect 284574 228520 284630 228576
rect 284758 343168 284814 343224
rect 284666 224304 284722 224360
rect 284390 221584 284446 221640
rect 284298 203632 284354 203688
rect 287058 352688 287114 352744
rect 285034 347248 285090 347304
rect 284942 340448 284998 340504
rect 284850 238040 284906 238096
rect 285126 341808 285182 341864
rect 286138 333648 286194 333704
rect 285862 329568 285918 329624
rect 285678 321408 285734 321464
rect 285126 237088 285182 237144
rect 285218 235456 285274 235512
rect 285034 231104 285090 231160
rect 284942 200640 284998 200696
rect 284758 197920 284814 197976
rect 285770 320048 285826 320104
rect 285954 324128 286010 324184
rect 285862 222808 285918 222864
rect 286046 322768 286102 322824
rect 285954 221448 286010 221504
rect 286506 330928 286562 330984
rect 286414 328208 286470 328264
rect 286230 326848 286286 326904
rect 286138 232464 286194 232520
rect 286322 325488 286378 325544
rect 286506 236680 286562 236736
rect 286414 233960 286470 234016
rect 286322 229744 286378 229800
rect 286230 226888 286286 226944
rect 286046 220088 286102 220144
rect 285770 204856 285826 204912
rect 285678 88984 285734 89040
rect 284942 83408 284998 83464
rect 286598 4936 286654 4992
rect 284942 3304 284998 3360
rect 287426 288768 287482 288824
rect 287610 282920 287666 282976
rect 287518 281832 287574 281888
rect 287518 279248 287574 279304
rect 287610 277888 287666 277944
rect 287426 241440 287482 241496
rect 288438 332288 288494 332344
rect 287058 3712 287114 3768
rect 289174 475904 289230 475960
rect 289450 481072 289506 481128
rect 289266 464480 289322 464536
rect 288990 442856 289046 442912
rect 289634 481480 289690 481536
rect 289542 473184 289598 473240
rect 290002 556144 290058 556200
rect 289910 479848 289966 479904
rect 290094 548800 290150 548856
rect 290002 478624 290058 478680
rect 290370 544720 290426 544776
rect 290278 540640 290334 540696
rect 290186 536560 290242 536616
rect 290094 476856 290150 476912
rect 290462 532480 290518 532536
rect 290370 478488 290426 478544
rect 290278 474272 290334 474328
rect 291198 512080 291254 512136
rect 290462 472368 290518 472424
rect 290186 467472 290242 467528
rect 289818 459040 289874 459096
rect 289726 442856 289782 442912
rect 289634 442040 289690 442096
rect 289634 441904 289690 441960
rect 291198 495352 291254 495408
rect 290646 487600 290702 487656
rect 290646 479712 290702 479768
rect 291934 601840 291990 601896
rect 291474 597760 291530 597816
rect 291382 593680 291438 593736
rect 291290 481480 291346 481536
rect 291566 589600 291622 589656
rect 291474 480256 291530 480312
rect 291658 585520 291714 585576
rect 291566 476992 291622 477048
rect 291382 475224 291438 475280
rect 291750 577360 291806 577416
rect 291842 520240 291898 520296
rect 291750 478760 291806 478816
rect 291658 474408 291714 474464
rect 291198 465976 291254 466032
rect 292026 503920 292082 503976
rect 291934 471552 291990 471608
rect 291842 462984 291898 463040
rect 292026 460264 292082 460320
rect 290554 442176 290610 442232
rect 288898 386688 288954 386744
rect 291198 335008 291254 335064
rect 288898 239400 288954 239456
rect 290186 4800 290242 4856
rect 288438 3440 288494 3496
rect 294050 700848 294106 700904
rect 293222 700440 293278 700496
rect 292946 633256 293002 633312
rect 293130 524320 293186 524376
rect 292946 478352 293002 478408
rect 292854 475632 292910 475688
rect 292762 442856 292818 442912
rect 293130 442448 293186 442504
rect 293958 700168 294014 700224
rect 293222 441904 293278 441960
rect 292578 269728 292634 269784
rect 298742 700440 298798 700496
rect 295338 700304 295394 700360
rect 295982 700304 296038 700360
rect 294234 632032 294290 632088
rect 294418 528400 294474 528456
rect 294234 478216 294290 478272
rect 294510 483520 294566 483576
rect 294510 475768 294566 475824
rect 294418 442312 294474 442368
rect 295430 569200 295486 569256
rect 295430 442720 295486 442776
rect 295338 271088 295394 271144
rect 294050 268368 294106 268424
rect 293958 267008 294014 267064
rect 296718 573280 296774 573336
rect 296810 561040 296866 561096
rect 296810 476040 296866 476096
rect 296718 442584 296774 442640
rect 302882 700576 302938 700632
rect 300122 657192 300178 657248
rect 300122 635432 300178 635488
rect 300122 598168 300178 598224
rect 300122 443400 300178 443456
rect 348790 700576 348846 700632
rect 353942 658824 353998 658880
rect 332506 450744 332562 450800
rect 302882 265648 302938 265704
rect 298742 264288 298798 264344
rect 295982 262928 296038 262984
rect 364982 657328 365038 657384
rect 364982 652024 365038 652080
rect 413650 700440 413706 700496
rect 429842 657600 429898 657656
rect 429842 634208 429898 634264
rect 478510 700304 478566 700360
rect 474646 657736 474702 657792
rect 474738 634072 474794 634128
rect 397458 449520 397514 449576
rect 508502 700304 508558 700360
rect 507122 670656 507178 670712
rect 489366 658008 489422 658064
rect 487158 657736 487214 657792
rect 488170 641144 488226 641200
rect 487802 636792 487858 636848
rect 487802 613672 487858 613728
rect 487802 472504 487858 472560
rect 353942 261568 353998 261624
rect 505098 658008 505154 658064
rect 494702 657872 494758 657928
rect 494610 657736 494666 657792
rect 501786 655596 501788 655616
rect 501788 655596 501840 655616
rect 501840 655596 501842 655616
rect 501786 655560 501842 655596
rect 500406 654880 500462 654936
rect 505926 656512 505982 656568
rect 559654 700304 559710 700360
rect 580262 697176 580318 697232
rect 543462 658824 543518 658880
rect 510066 657736 510122 657792
rect 508502 655832 508558 655888
rect 507122 655696 507178 655752
rect 511446 657600 511502 657656
rect 515586 657464 515642 657520
rect 512826 657328 512882 657384
rect 514206 657192 514262 657248
rect 516966 657056 517022 657112
rect 525246 656376 525302 656432
rect 522486 656240 522542 656296
rect 519726 656104 519782 656160
rect 518346 655968 518402 656024
rect 494610 654744 494666 654800
rect 523866 654608 523922 654664
rect 521106 654472 521162 654528
rect 490470 653656 490526 653712
rect 489366 649168 489422 649224
rect 540150 651208 540206 651264
rect 539782 642504 539838 642560
rect 539598 637744 539654 637800
rect 490746 475496 490802 475552
rect 493506 465840 493562 465896
rect 492126 462848 492182 462904
rect 496266 468560 496322 468616
rect 494886 448160 494942 448216
rect 497646 446800 497702 446856
rect 500406 448024 500462 448080
rect 504546 475360 504602 475416
rect 503166 473048 503222 473104
rect 510066 472912 510122 472968
rect 501786 445304 501842 445360
rect 499026 443808 499082 443864
rect 311438 86128 311494 86184
rect 304354 51720 304410 51776
rect 293682 46280 293738 46336
rect 291198 3576 291254 3632
rect 297270 43560 297326 43616
rect 300766 42200 300822 42256
rect 307942 50224 307998 50280
rect 322110 85720 322166 85776
rect 318522 80688 318578 80744
rect 315026 53080 315082 53136
rect 336278 85584 336334 85640
rect 325606 69536 325662 69592
rect 329194 54576 329250 54632
rect 332690 9016 332746 9072
rect 368202 84904 368258 84960
rect 357530 84768 357586 84824
rect 343362 84632 343418 84688
rect 353942 57160 353998 57216
rect 351182 55800 351238 55856
rect 353942 7520 353998 7576
rect 351182 4800 351238 4856
rect 361118 84496 361174 84552
rect 435362 83000 435418 83056
rect 432602 81640 432658 81696
rect 428554 80280 428610 80336
rect 421562 77560 421618 77616
rect 417422 76200 417478 76256
rect 414662 74840 414718 74896
rect 406382 63960 406438 64016
rect 400126 40704 400182 40760
rect 378874 21256 378930 21312
rect 375286 10376 375342 10432
rect 371698 3304 371754 3360
rect 396538 17312 396594 17368
rect 393042 15952 393098 16008
rect 389454 14592 389510 14648
rect 385958 13096 386014 13152
rect 382370 11736 382426 11792
rect 403622 22752 403678 22808
rect 411902 58520 411958 58576
rect 407210 39344 407266 39400
rect 406382 7656 406438 7712
rect 414294 7520 414350 7576
rect 410798 4800 410854 4856
rect 411902 4800 411958 4856
rect 418802 59880 418858 59936
rect 417882 4800 417938 4856
rect 417422 3440 417478 3496
rect 414662 3032 414718 3088
rect 418802 4120 418858 4176
rect 421378 4120 421434 4176
rect 425702 62600 425758 62656
rect 422942 61240 422998 61296
rect 422942 4120 422998 4176
rect 424966 4120 425022 4176
rect 425702 4120 425758 4176
rect 428462 4120 428518 4176
rect 421562 3848 421618 3904
rect 431222 68040 431278 68096
rect 429842 65320 429898 65376
rect 432050 7656 432106 7712
rect 431222 7520 431278 7576
rect 429842 4800 429898 4856
rect 428554 3712 428610 3768
rect 450542 73480 450598 73536
rect 447782 72120 447838 72176
rect 443642 70760 443698 70816
rect 436742 66680 436798 66736
rect 435546 4800 435602 4856
rect 435362 3576 435418 3632
rect 432602 3168 432658 3224
rect 439502 47776 439558 47832
rect 436742 4120 436798 4176
rect 439134 4120 439190 4176
rect 442262 47640 442318 47696
rect 439502 3984 439558 4040
rect 442630 7520 442686 7576
rect 442262 3304 442318 3360
rect 446402 47504 446458 47560
rect 443642 4120 443698 4176
rect 446218 4120 446274 4176
rect 442906 3984 442962 4040
rect 467470 50360 467526 50416
rect 450542 4800 450598 4856
rect 453302 4800 453358 4856
rect 447782 4120 447838 4176
rect 449806 4120 449862 4176
rect 463974 3848 464030 3904
rect 460386 3440 460442 3496
rect 456890 3032 456946 3088
rect 512826 471280 512882 471336
rect 511446 464344 511502 464400
rect 514206 460128 514262 460184
rect 515586 447752 515642 447808
rect 519726 472776 519782 472832
rect 521106 449384 521162 449440
rect 518346 447888 518402 447944
rect 523866 472640 523922 472696
rect 528006 458904 528062 458960
rect 530766 598168 530822 598224
rect 532146 474136 532202 474192
rect 533526 467200 533582 467256
rect 534906 467064 534962 467120
rect 536286 453192 536342 453248
rect 529386 450608 529442 450664
rect 537666 446528 537722 446584
rect 522486 445168 522542 445224
rect 516966 443672 517022 443728
rect 539690 633256 539746 633312
rect 539598 443536 539654 443592
rect 539966 630944 540022 631000
rect 539874 627816 539930 627872
rect 539782 449248 539838 449304
rect 540058 625504 540114 625560
rect 539966 446664 540022 446720
rect 546498 649848 546554 649904
rect 543738 648488 543794 648544
rect 542634 640328 542690 640384
rect 540978 638968 541034 639024
rect 540058 445032 540114 445088
rect 541070 622648 541126 622704
rect 541162 621288 541218 621344
rect 542450 615848 542506 615904
rect 542358 613128 542414 613184
rect 542542 610408 542598 610464
rect 542450 449112 542506 449168
rect 542358 446392 542414 446448
rect 542726 634888 542782 634944
rect 543002 632168 543058 632224
rect 542910 614488 542966 614544
rect 542818 609048 542874 609104
rect 543094 629448 543150 629504
rect 543186 611768 543242 611824
rect 543094 479576 543150 479632
rect 543186 471144 543242 471200
rect 545118 647128 545174 647184
rect 543830 645768 543886 645824
rect 543738 469784 543794 469840
rect 543922 641688 543978 641744
rect 544106 624008 544162 624064
rect 544014 619928 544070 619984
rect 544198 617208 544254 617264
rect 543922 470328 543978 470384
rect 545210 644408 545266 644464
rect 545302 626728 545358 626784
rect 545210 470464 545266 470520
rect 545302 470192 545358 470248
rect 545118 470056 545174 470112
rect 546498 469920 546554 469976
rect 543830 469648 543886 469704
rect 542910 458768 542966 458824
rect 542818 451832 542874 451888
rect 542542 444896 542598 444952
rect 580262 465704 580318 465760
rect 580538 656920 580594 656976
rect 580538 617480 580594 617536
rect 580538 590960 580594 591016
rect 580446 511264 580502 511320
rect 580722 644000 580778 644056
rect 580630 564304 580686 564360
rect 580630 537784 580686 537840
rect 580354 458088 580410 458144
rect 580262 431568 580318 431624
rect 579710 404912 579766 404968
rect 580262 378392 580318 378448
rect 580170 351872 580226 351928
rect 580170 298696 580226 298752
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580262 240216 580318 240272
rect 580262 236544 580318 236600
rect 580170 205672 580226 205728
rect 580170 165824 580226 165880
rect 580170 86128 580226 86184
rect 520738 48864 520794 48920
rect 481730 46144 481786 46200
rect 471058 3712 471114 3768
rect 478142 3576 478198 3632
rect 474554 3168 474610 3224
rect 502982 43424 503038 43480
rect 499394 14456 499450 14512
rect 495898 12960 495954 13016
rect 492310 11600 492366 11656
rect 488814 10240 488870 10296
rect 485226 8880 485282 8936
rect 508502 42064 508558 42120
rect 506478 15816 506534 15872
rect 512642 40568 512698 40624
rect 508502 3984 508558 4040
rect 510066 3984 510122 4040
rect 517150 25472 517206 25528
rect 512642 3440 512698 3496
rect 513562 3440 513618 3496
rect 580170 46280 580226 46336
rect 549074 44784 549130 44840
rect 524234 39208 524290 39264
rect 531318 37848 531374 37904
rect 527822 17176 527878 17232
rect 534906 36488 534962 36544
rect 538402 35128 538458 35184
rect 541990 33768 542046 33824
rect 545486 32408 545542 32464
rect 580354 235184 580410 235240
rect 580354 72936 580410 72992
rect 580262 33088 580318 33144
rect 552662 30912 552718 30968
rect 556158 29552 556214 29608
rect 562322 28192 562378 28248
rect 559746 18536 559802 18592
rect 566830 26832 566886 26888
rect 562322 3440 562378 3496
rect 563242 3440 563298 3496
rect 570326 24112 570382 24168
rect 573914 22616 573970 22672
rect 576122 19896 576178 19952
rect 580170 6568 580226 6624
rect 576122 3984 576178 4040
rect 577410 3984 577466 4040
rect 582194 3304 582250 3360
<< metal3 >>
rect 267641 701042 267707 701045
rect 292849 701042 292915 701045
rect 267641 701040 292915 701042
rect 267641 700984 267646 701040
rect 267702 700984 292854 701040
rect 292910 700984 292915 701040
rect 267641 700982 292915 700984
rect 267641 700979 267707 700982
rect 292849 700979 292915 700982
rect 218973 700906 219039 700909
rect 294045 700906 294111 700909
rect 218973 700904 294111 700906
rect 218973 700848 218978 700904
rect 219034 700848 294050 700904
rect 294106 700848 294111 700904
rect 218973 700846 294111 700848
rect 218973 700843 219039 700846
rect 294045 700843 294111 700846
rect 170305 700770 170371 700773
rect 189717 700770 189783 700773
rect 170305 700768 189783 700770
rect 170305 700712 170310 700768
rect 170366 700712 189722 700768
rect 189778 700712 189783 700768
rect 170305 700710 189783 700712
rect 170305 700707 170371 700710
rect 189717 700707 189783 700710
rect 202781 700770 202847 700773
rect 292757 700770 292823 700773
rect 202781 700768 292823 700770
rect 202781 700712 202786 700768
rect 202842 700712 292762 700768
rect 292818 700712 292823 700768
rect 202781 700710 292823 700712
rect 202781 700707 202847 700710
rect 292757 700707 292823 700710
rect 154113 700634 154179 700637
rect 292573 700634 292639 700637
rect 154113 700632 292639 700634
rect 154113 700576 154118 700632
rect 154174 700576 292578 700632
rect 292634 700576 292639 700632
rect 154113 700574 292639 700576
rect 154113 700571 154179 700574
rect 292573 700571 292639 700574
rect 302877 700634 302943 700637
rect 348785 700634 348851 700637
rect 302877 700632 348851 700634
rect 302877 700576 302882 700632
rect 302938 700576 348790 700632
rect 348846 700576 348851 700632
rect 302877 700574 348851 700576
rect 302877 700571 302943 700574
rect 348785 700571 348851 700574
rect 24301 700498 24367 700501
rect 59997 700498 60063 700501
rect 24301 700496 60063 700498
rect 24301 700440 24306 700496
rect 24362 700440 60002 700496
rect 60058 700440 60063 700496
rect 24301 700438 60063 700440
rect 24301 700435 24367 700438
rect 59997 700435 60063 700438
rect 137829 700498 137895 700501
rect 293217 700498 293283 700501
rect 137829 700496 293283 700498
rect 137829 700440 137834 700496
rect 137890 700440 293222 700496
rect 293278 700440 293283 700496
rect 137829 700438 293283 700440
rect 137829 700435 137895 700438
rect 293217 700435 293283 700438
rect 298737 700498 298803 700501
rect 413645 700498 413711 700501
rect 298737 700496 413711 700498
rect 298737 700440 298742 700496
rect 298798 700440 413650 700496
rect 413706 700440 413711 700496
rect 298737 700438 413711 700440
rect 298737 700435 298803 700438
rect 413645 700435 413711 700438
rect 40493 700362 40559 700365
rect 86217 700362 86283 700365
rect 40493 700360 86283 700362
rect 40493 700304 40498 700360
rect 40554 700304 86222 700360
rect 86278 700304 86283 700360
rect 40493 700302 86283 700304
rect 40493 700299 40559 700302
rect 86217 700299 86283 700302
rect 89161 700362 89227 700365
rect 295333 700362 295399 700365
rect 89161 700360 295399 700362
rect 89161 700304 89166 700360
rect 89222 700304 295338 700360
rect 295394 700304 295399 700360
rect 89161 700302 295399 700304
rect 89161 700299 89227 700302
rect 295333 700299 295399 700302
rect 295977 700362 296043 700365
rect 478505 700362 478571 700365
rect 295977 700360 478571 700362
rect 295977 700304 295982 700360
rect 296038 700304 478510 700360
rect 478566 700304 478571 700360
rect 295977 700302 478571 700304
rect 295977 700299 296043 700302
rect 478505 700299 478571 700302
rect 508497 700362 508563 700365
rect 559649 700362 559715 700365
rect 508497 700360 559715 700362
rect 508497 700304 508502 700360
rect 508558 700304 559654 700360
rect 559710 700304 559715 700360
rect 508497 700302 559715 700304
rect 508497 700299 508563 700302
rect 559649 700299 559715 700302
rect 283833 700226 283899 700229
rect 293953 700226 294019 700229
rect 283833 700224 294019 700226
rect 283833 700168 283838 700224
rect 283894 700168 293958 700224
rect 294014 700168 294019 700224
rect 283833 700166 294019 700168
rect 283833 700163 283899 700166
rect 293953 700163 294019 700166
rect -960 697220 480 697460
rect 580257 697234 580323 697237
rect 583520 697234 584960 697324
rect 580257 697232 584960 697234
rect 580257 697176 580262 697232
rect 580318 697176 584960 697232
rect 580257 697174 584960 697176
rect 580257 697171 580323 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 355174 683844 355180 683908
rect 355244 683906 355250 683908
rect 583520 683906 584960 683996
rect 355244 683846 584960 683906
rect 355244 683844 355250 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 57278 671258 57284 671260
rect -960 671198 57284 671258
rect -960 671108 480 671198
rect 57278 671196 57284 671198
rect 57348 671196 57354 671260
rect 507117 670714 507183 670717
rect 583520 670714 584960 670804
rect 507117 670712 584960 670714
rect 507117 670656 507122 670712
rect 507178 670656 584960 670712
rect 507117 670654 584960 670656
rect 507117 670651 507183 670654
rect 583520 670564 584960 670654
rect 353937 658882 354003 658885
rect 543457 658882 543523 658885
rect 353937 658880 543523 658882
rect 353937 658824 353942 658880
rect 353998 658824 543462 658880
rect 543518 658824 543523 658880
rect 353937 658822 543523 658824
rect 353937 658819 354003 658822
rect 543457 658819 543523 658822
rect -960 658202 480 658292
rect 2814 658202 2820 658204
rect -960 658142 2820 658202
rect -960 658052 480 658142
rect 2814 658140 2820 658142
rect 2884 658140 2890 658204
rect 489361 658066 489427 658069
rect 505093 658066 505159 658069
rect 489361 658064 505159 658066
rect 489361 658008 489366 658064
rect 489422 658008 505098 658064
rect 505154 658008 505159 658064
rect 489361 658006 505159 658008
rect 489361 658003 489427 658006
rect 505093 658003 505159 658006
rect 134425 657930 134491 657933
rect 494697 657930 494763 657933
rect 134425 657928 494763 657930
rect 134425 657872 134430 657928
rect 134486 657872 494702 657928
rect 494758 657872 494763 657928
rect 134425 657870 494763 657872
rect 134425 657867 134491 657870
rect 494697 657867 494763 657870
rect 474641 657794 474707 657797
rect 487153 657794 487219 657797
rect 474641 657792 487219 657794
rect 474641 657736 474646 657792
rect 474702 657736 487158 657792
rect 487214 657736 487219 657792
rect 474641 657734 487219 657736
rect 474641 657731 474707 657734
rect 487153 657731 487219 657734
rect 494605 657794 494671 657797
rect 510061 657794 510127 657797
rect 494605 657792 510127 657794
rect 494605 657736 494610 657792
rect 494666 657736 510066 657792
rect 510122 657736 510127 657792
rect 494605 657734 510127 657736
rect 494605 657731 494671 657734
rect 510061 657731 510127 657734
rect 429837 657658 429903 657661
rect 511441 657658 511507 657661
rect 429837 657656 511507 657658
rect 429837 657600 429842 657656
rect 429898 657600 511446 657656
rect 511502 657600 511507 657656
rect 429837 657598 511507 657600
rect 429837 657595 429903 657598
rect 511441 657595 511507 657598
rect 183001 657522 183067 657525
rect 235165 657522 235231 657525
rect 515581 657522 515647 657525
rect 183001 657520 515647 657522
rect 183001 657464 183006 657520
rect 183062 657464 235170 657520
rect 235226 657464 515586 657520
rect 515642 657464 515647 657520
rect 183001 657462 515647 657464
rect 183001 657459 183067 657462
rect 235165 657459 235231 657462
rect 515581 657459 515647 657462
rect 364977 657386 365043 657389
rect 512821 657386 512887 657389
rect 364977 657384 512887 657386
rect 364977 657328 364982 657384
rect 365038 657328 512826 657384
rect 512882 657328 512887 657384
rect 364977 657326 512887 657328
rect 364977 657323 365043 657326
rect 512821 657323 512887 657326
rect 300117 657250 300183 657253
rect 514201 657250 514267 657253
rect 300117 657248 514267 657250
rect 300117 657192 300122 657248
rect 300178 657192 514206 657248
rect 514262 657192 514267 657248
rect 583520 657236 584960 657476
rect 300117 657190 514267 657192
rect 300117 657187 300183 657190
rect 514201 657187 514267 657190
rect 189073 657114 189139 657117
rect 189717 657114 189783 657117
rect 516961 657114 517027 657117
rect 189073 657112 517027 657114
rect 189073 657056 189078 657112
rect 189134 657056 189722 657112
rect 189778 657056 516966 657112
rect 517022 657056 517027 657112
rect 189073 657054 517027 657056
rect 189073 657051 189139 657054
rect 189717 657051 189783 657054
rect 516961 657051 517027 657054
rect 580533 656978 580599 656981
rect 506062 656976 580599 656978
rect 506062 656920 580538 656976
rect 580594 656920 580599 656976
rect 506062 656918 580599 656920
rect 140037 656570 140103 656573
rect 505921 656570 505987 656573
rect 506062 656570 506122 656918
rect 580533 656915 580599 656918
rect 140037 656568 506122 656570
rect 140037 656512 140042 656568
rect 140098 656512 505926 656568
rect 505982 656512 506122 656568
rect 140037 656510 506122 656512
rect 140037 656507 140103 656510
rect 505921 656507 505987 656510
rect 225505 656434 225571 656437
rect 525241 656434 525307 656437
rect 225505 656432 525307 656434
rect 225505 656376 225510 656432
rect 225566 656376 525246 656432
rect 525302 656376 525307 656432
rect 225505 656374 525307 656376
rect 225505 656371 225571 656374
rect 525241 656371 525307 656374
rect 213177 656298 213243 656301
rect 522481 656298 522547 656301
rect 213177 656296 522547 656298
rect 213177 656240 213182 656296
rect 213238 656240 522486 656296
rect 522542 656240 522547 656296
rect 213177 656238 522547 656240
rect 213177 656235 213243 656238
rect 522481 656235 522547 656238
rect 200757 656162 200823 656165
rect 519721 656162 519787 656165
rect 200757 656160 519787 656162
rect 200757 656104 200762 656160
rect 200818 656104 519726 656160
rect 519782 656104 519787 656160
rect 200757 656102 519787 656104
rect 200757 656099 200823 656102
rect 519721 656099 519787 656102
rect 195237 656026 195303 656029
rect 518341 656026 518407 656029
rect 195237 656024 518407 656026
rect 195237 655968 195242 656024
rect 195298 655968 518346 656024
rect 518402 655968 518407 656024
rect 195237 655966 518407 655968
rect 195237 655963 195303 655966
rect 518341 655963 518407 655966
rect 152457 655890 152523 655893
rect 508497 655890 508563 655893
rect 152457 655888 508563 655890
rect 152457 655832 152462 655888
rect 152518 655832 508502 655888
rect 508558 655832 508563 655888
rect 152457 655830 508563 655832
rect 152457 655827 152523 655830
rect 508497 655827 508563 655830
rect 146937 655754 147003 655757
rect 507117 655754 507183 655757
rect 146937 655752 507183 655754
rect 146937 655696 146942 655752
rect 146998 655696 507122 655752
rect 507178 655696 507183 655752
rect 146937 655694 507183 655696
rect 146937 655691 147003 655694
rect 507117 655691 507183 655694
rect 128997 655618 129063 655621
rect 224953 655618 225019 655621
rect 128997 655616 225019 655618
rect 128997 655560 129002 655616
rect 129058 655560 224958 655616
rect 225014 655560 225019 655616
rect 128997 655558 225019 655560
rect 128997 655555 129063 655558
rect 224953 655555 225019 655558
rect 501638 655556 501644 655620
rect 501708 655618 501714 655620
rect 501781 655618 501847 655621
rect 501708 655616 501847 655618
rect 501708 655560 501786 655616
rect 501842 655560 501847 655616
rect 501708 655558 501847 655560
rect 501708 655556 501714 655558
rect 501781 655555 501847 655558
rect 500401 654940 500467 654941
rect 500350 654938 500356 654940
rect 500310 654878 500356 654938
rect 500420 654936 500467 654940
rect 500462 654880 500467 654936
rect 500350 654876 500356 654878
rect 500420 654876 500467 654880
rect 500401 654875 500467 654876
rect 159357 654802 159423 654805
rect 494605 654802 494671 654805
rect 159357 654800 494671 654802
rect 159357 654744 159362 654800
rect 159418 654744 494610 654800
rect 494666 654744 494671 654800
rect 159357 654742 494671 654744
rect 159357 654739 159423 654742
rect 494605 654739 494671 654742
rect 219433 654666 219499 654669
rect 523861 654666 523927 654669
rect 219433 654664 523927 654666
rect 219433 654608 219438 654664
rect 219494 654608 523866 654664
rect 523922 654608 523927 654664
rect 219433 654606 523927 654608
rect 219433 654603 219499 654606
rect 523861 654603 523927 654606
rect 207657 654530 207723 654533
rect 521101 654530 521167 654533
rect 207657 654528 521167 654530
rect 207657 654472 207662 654528
rect 207718 654472 521106 654528
rect 521162 654472 521167 654528
rect 207657 654470 521167 654472
rect 207657 654467 207723 654470
rect 521101 654467 521167 654470
rect 501638 654332 501644 654396
rect 501708 654332 501714 654396
rect 501646 654122 501706 654332
rect 499530 654062 501706 654122
rect 262121 653714 262187 653717
rect 490465 653714 490531 653717
rect 262121 653712 490531 653714
rect 262121 653656 262126 653712
rect 262182 653656 490470 653712
rect 490526 653656 490531 653712
rect 262121 653654 490531 653656
rect 262121 653651 262187 653654
rect 490465 653651 490531 653654
rect 122281 653578 122347 653581
rect 499530 653578 499590 654062
rect 122281 653576 499590 653578
rect 122281 653520 122286 653576
rect 122342 653520 499590 653576
rect 122281 653518 499590 653520
rect 122281 653515 122347 653518
rect 116209 653442 116275 653445
rect 500350 653442 500356 653444
rect 116209 653440 500356 653442
rect 116209 653384 116214 653440
rect 116270 653384 500356 653440
rect 116209 653382 500356 653384
rect 116209 653379 116275 653382
rect 500350 653380 500356 653382
rect 500420 653380 500426 653444
rect 170857 652082 170923 652085
rect 364977 652082 365043 652085
rect 170857 652080 365043 652082
rect 170857 652024 170862 652080
rect 170918 652024 364982 652080
rect 365038 652024 365043 652080
rect 170857 652022 365043 652024
rect 170857 652019 170923 652022
rect 364977 652019 365043 652022
rect 540145 651266 540211 651269
rect 539948 651264 540211 651266
rect 539948 651208 540150 651264
rect 540206 651208 540211 651264
rect 539948 651206 540211 651208
rect 540145 651203 540211 651206
rect 546493 649906 546559 649909
rect 539948 649904 546559 649906
rect 539948 649848 546498 649904
rect 546554 649848 546559 649904
rect 539948 649846 546559 649848
rect 546493 649843 546559 649846
rect 249793 649226 249859 649229
rect 489361 649226 489427 649229
rect 249793 649224 489427 649226
rect 249793 649168 249798 649224
rect 249854 649168 489366 649224
rect 489422 649168 489427 649224
rect 249793 649166 489427 649168
rect 249793 649163 249859 649166
rect 489361 649163 489427 649166
rect 543733 648546 543799 648549
rect 539948 648544 543799 648546
rect 539948 648488 543738 648544
rect 543794 648488 543799 648544
rect 539948 648486 543799 648488
rect 543733 648483 543799 648486
rect 545113 647186 545179 647189
rect 539948 647184 545179 647186
rect 539948 647128 545118 647184
rect 545174 647128 545179 647184
rect 539948 647126 545179 647128
rect 545113 647123 545179 647126
rect 543825 645826 543891 645829
rect 539948 645824 543891 645826
rect 539948 645768 543830 645824
rect 543886 645768 543891 645824
rect 539948 645766 543891 645768
rect 543825 645763 543891 645766
rect -960 644996 480 645236
rect 545205 644466 545271 644469
rect 539948 644464 545271 644466
rect 539948 644408 545210 644464
rect 545266 644408 545271 644464
rect 539948 644406 545271 644408
rect 545205 644403 545271 644406
rect 580717 644058 580783 644061
rect 583520 644058 584960 644148
rect 580717 644056 584960 644058
rect 580717 644000 580722 644056
rect 580778 644000 584960 644056
rect 580717 643998 584960 644000
rect 580717 643995 580783 643998
rect 583520 643908 584960 643998
rect 539734 642565 539794 643076
rect 539734 642560 539843 642565
rect 539734 642504 539782 642560
rect 539838 642504 539843 642560
rect 539734 642502 539843 642504
rect 539777 642499 539843 642502
rect 543917 641746 543983 641749
rect 539948 641744 543983 641746
rect 539948 641688 543922 641744
rect 543978 641688 543983 641744
rect 539948 641686 543983 641688
rect 543917 641683 543983 641686
rect 488165 641202 488231 641205
rect 488165 641200 490084 641202
rect 488165 641144 488170 641200
rect 488226 641144 490084 641200
rect 488165 641142 490084 641144
rect 488165 641139 488231 641142
rect 542629 640386 542695 640389
rect 539948 640384 542695 640386
rect 539948 640328 542634 640384
rect 542690 640328 542695 640384
rect 539948 640326 542695 640328
rect 542629 640323 542695 640326
rect 540973 639026 541039 639029
rect 539948 639024 541039 639026
rect 539948 638968 540978 639024
rect 541034 638968 541039 639024
rect 539948 638966 541039 638968
rect 540973 638963 541039 638966
rect 539593 637802 539659 637805
rect 539550 637800 539659 637802
rect 539550 637744 539598 637800
rect 539654 637744 539659 637800
rect 539550 637739 539659 637744
rect 539550 637636 539610 637739
rect 289813 636850 289879 636853
rect 487797 636850 487863 636853
rect 289813 636848 487863 636850
rect 289813 636792 289818 636848
rect 289874 636792 487802 636848
rect 487858 636792 487863 636848
rect 289813 636790 487863 636792
rect 289813 636787 289879 636790
rect 487797 636787 487863 636790
rect 542670 636306 542676 636308
rect 539948 636246 542676 636306
rect 542670 636244 542676 636246
rect 542740 636244 542746 636308
rect 176929 635490 176995 635493
rect 300117 635490 300183 635493
rect 176929 635488 300183 635490
rect 176929 635432 176934 635488
rect 176990 635432 300122 635488
rect 300178 635432 300183 635488
rect 176929 635430 300183 635432
rect 176929 635427 176995 635430
rect 300117 635427 300183 635430
rect 542721 634946 542787 634949
rect 539948 634944 542787 634946
rect 539948 634888 542726 634944
rect 542782 634888 542787 634944
rect 539948 634886 542787 634888
rect 542721 634883 542787 634886
rect 164785 634266 164851 634269
rect 429837 634266 429903 634269
rect 164785 634264 429903 634266
rect 164785 634208 164790 634264
rect 164846 634208 429842 634264
rect 429898 634208 429903 634264
rect 164785 634206 429903 634208
rect 164785 634203 164851 634206
rect 429837 634203 429903 634206
rect 104065 634130 104131 634133
rect 474733 634130 474799 634133
rect 104065 634128 474799 634130
rect 104065 634072 104070 634128
rect 104126 634072 474738 634128
rect 474794 634072 474799 634128
rect 104065 634070 474799 634072
rect 104065 634067 104131 634070
rect 474733 634067 474799 634070
rect 539734 633317 539794 633556
rect 105445 633314 105511 633317
rect 195237 633314 195303 633317
rect 289813 633314 289879 633317
rect 292941 633314 293007 633317
rect 103470 633312 195303 633314
rect 103470 633256 105450 633312
rect 105506 633256 195242 633312
rect 195298 633256 195303 633312
rect 103470 633254 195303 633256
rect 69933 633178 69999 633181
rect 88241 633178 88307 633181
rect 69933 633176 88307 633178
rect 69933 633120 69938 633176
rect 69994 633120 88246 633176
rect 88302 633120 88307 633176
rect 69933 633118 88307 633120
rect 69933 633115 69999 633118
rect 88241 633115 88307 633118
rect 69841 632906 69907 632909
rect 103470 632906 103530 633254
rect 105445 633251 105511 633254
rect 195237 633251 195303 633254
rect 277350 633312 293007 633314
rect 277350 633256 289818 633312
rect 289874 633256 292946 633312
rect 293002 633256 293007 633312
rect 277350 633254 293007 633256
rect 69841 632904 103530 632906
rect 69841 632848 69846 632904
rect 69902 632848 103530 632904
rect 69841 632846 103530 632848
rect 69841 632843 69907 632846
rect 70025 632770 70091 632773
rect 152641 632770 152707 632773
rect 70025 632768 152707 632770
rect 70025 632712 70030 632768
rect 70086 632712 152646 632768
rect 152702 632712 152707 632768
rect 70025 632710 152707 632712
rect 70025 632707 70091 632710
rect 152641 632707 152707 632710
rect 64781 632634 64847 632637
rect 158713 632634 158779 632637
rect 159357 632634 159423 632637
rect 64781 632632 159423 632634
rect 64781 632576 64786 632632
rect 64842 632576 158718 632632
rect 158774 632576 159362 632632
rect 159418 632576 159423 632632
rect 64781 632574 159423 632576
rect 64781 632571 64847 632574
rect 158713 632571 158779 632574
rect 159357 632571 159423 632574
rect 66069 632498 66135 632501
rect 164785 632498 164851 632501
rect 66069 632496 164851 632498
rect 66069 632440 66074 632496
rect 66130 632440 164790 632496
rect 164846 632440 164851 632496
rect 66069 632438 164851 632440
rect 66069 632435 66135 632438
rect 164785 632435 164851 632438
rect 86217 632362 86283 632365
rect 200849 632362 200915 632365
rect 201217 632362 201283 632365
rect 86217 632360 201283 632362
rect 86217 632304 86222 632360
rect 86278 632304 200854 632360
rect 200910 632304 201222 632360
rect 201278 632304 201283 632360
rect 86217 632302 201283 632304
rect 86217 632299 86283 632302
rect 200849 632299 200915 632302
rect 201217 632299 201283 632302
rect 52637 632226 52703 632229
rect 79777 632226 79843 632229
rect 86861 632226 86927 632229
rect 52637 632224 86927 632226
rect -960 632090 480 632180
rect 52637 632168 52642 632224
rect 52698 632168 79782 632224
rect 79838 632168 86866 632224
rect 86922 632168 86927 632224
rect 52637 632166 86927 632168
rect 52637 632163 52703 632166
rect 79777 632163 79843 632166
rect 86861 632163 86927 632166
rect 87597 632226 87663 632229
rect 207657 632226 207723 632229
rect 87597 632224 207723 632226
rect 87597 632168 87602 632224
rect 87658 632168 207662 632224
rect 207718 632168 207723 632224
rect 87597 632166 207723 632168
rect 87597 632163 87663 632166
rect 207657 632163 207723 632166
rect 268009 632226 268075 632229
rect 277350 632226 277410 633254
rect 289813 633251 289879 633254
rect 292941 633251 293007 633254
rect 539685 633312 539794 633317
rect 539685 633256 539690 633312
rect 539746 633256 539794 633312
rect 539685 633254 539794 633256
rect 539685 633251 539751 633254
rect 542997 632226 543063 632229
rect 268009 632224 277410 632226
rect 268009 632168 268014 632224
rect 268070 632168 277410 632224
rect 268009 632166 277410 632168
rect 539948 632224 543063 632226
rect 539948 632168 543002 632224
rect 543058 632168 543063 632224
rect 539948 632166 543063 632168
rect 268009 632163 268075 632166
rect 542997 632163 543063 632166
rect 60641 632090 60707 632093
rect 213177 632090 213243 632093
rect -960 632088 213243 632090
rect -960 632032 60646 632088
rect 60702 632032 213182 632088
rect 213238 632032 213243 632088
rect -960 632030 213243 632032
rect -960 631940 480 632030
rect 60641 632027 60707 632030
rect 213177 632027 213243 632030
rect 262121 632090 262187 632093
rect 294229 632090 294295 632093
rect 262121 632088 294295 632090
rect 262121 632032 262126 632088
rect 262182 632032 294234 632088
rect 294290 632032 294295 632088
rect 262121 632030 294295 632032
rect 262121 632027 262187 632030
rect 294229 632027 294295 632030
rect 62021 631546 62087 631549
rect 72969 631546 73035 631549
rect 62021 631544 73035 631546
rect 62021 631488 62026 631544
rect 62082 631488 72974 631544
rect 73030 631488 73035 631544
rect 62021 631486 73035 631488
rect 62021 631483 62087 631486
rect 72969 631483 73035 631486
rect 66161 631410 66227 631413
rect 86217 631410 86283 631413
rect 66161 631408 86283 631410
rect 66161 631352 66166 631408
rect 66222 631352 86222 631408
rect 86278 631352 86283 631408
rect 66161 631350 86283 631352
rect 66161 631347 66227 631350
rect 86217 631347 86283 631350
rect 63401 631274 63467 631277
rect 87597 631274 87663 631277
rect 63401 631272 87663 631274
rect 63401 631216 63406 631272
rect 63462 631216 87602 631272
rect 87658 631216 87663 631272
rect 63401 631214 87663 631216
rect 63401 631211 63467 631214
rect 87597 631211 87663 631214
rect 70209 631002 70275 631005
rect 110137 631002 110203 631005
rect 539961 631002 540027 631005
rect 70209 631000 110203 631002
rect 70209 630944 70214 631000
rect 70270 630944 110142 631000
rect 110198 630944 110203 631000
rect 70209 630942 110203 630944
rect 70209 630939 70275 630942
rect 110137 630939 110203 630942
rect 539918 631000 540027 631002
rect 539918 630944 539966 631000
rect 540022 630944 540027 631000
rect 539918 630939 540027 630944
rect 69197 630866 69263 630869
rect 140129 630866 140195 630869
rect 140497 630866 140563 630869
rect 69197 630864 140563 630866
rect 69197 630808 69202 630864
rect 69258 630808 140134 630864
rect 140190 630808 140502 630864
rect 140558 630808 140563 630864
rect 539918 630836 539978 630939
rect 69197 630806 140563 630808
rect 69197 630803 69263 630806
rect 140129 630803 140195 630806
rect 140497 630803 140563 630806
rect 580206 630804 580212 630868
rect 580276 630866 580282 630868
rect 583520 630866 584960 630956
rect 580276 630806 584960 630866
rect 580276 630804 580282 630806
rect 70577 630730 70643 630733
rect 146937 630730 147003 630733
rect 70577 630728 147003 630730
rect 70577 630672 70582 630728
rect 70638 630672 146942 630728
rect 146998 630672 147003 630728
rect 583520 630716 584960 630806
rect 70577 630670 147003 630672
rect 70577 630667 70643 630670
rect 146937 630667 147003 630670
rect 63217 630322 63283 630325
rect 68921 630322 68987 630325
rect 63217 630320 68987 630322
rect 63217 630264 63222 630320
rect 63278 630264 68926 630320
rect 68982 630264 68987 630320
rect 63217 630262 68987 630264
rect 63217 630259 63283 630262
rect 68921 630259 68987 630262
rect 63125 630186 63191 630189
rect 170857 630186 170923 630189
rect 63125 630184 170923 630186
rect 63125 630128 63130 630184
rect 63186 630128 170862 630184
rect 170918 630128 170923 630184
rect 63125 630126 170923 630128
rect 63125 630123 63191 630126
rect 170857 630123 170923 630126
rect 67357 630050 67423 630053
rect 176653 630050 176719 630053
rect 67357 630048 176719 630050
rect 67357 629992 67362 630048
rect 67418 629992 176658 630048
rect 176714 629992 176719 630048
rect 67357 629990 176719 629992
rect 67357 629987 67423 629990
rect 176653 629987 176719 629990
rect 64689 629914 64755 629917
rect 183001 629914 183067 629917
rect 64689 629912 183067 629914
rect 64689 629856 64694 629912
rect 64750 629856 183006 629912
rect 183062 629856 183067 629912
rect 64689 629854 183067 629856
rect 64689 629851 64755 629854
rect 183001 629851 183067 629854
rect 61929 629778 61995 629781
rect 189073 629778 189139 629781
rect 61929 629776 189139 629778
rect 61929 629720 61934 629776
rect 61990 629720 189078 629776
rect 189134 629720 189139 629776
rect 61929 629718 189139 629720
rect 61929 629715 61995 629718
rect 189073 629715 189139 629718
rect 61837 629642 61903 629645
rect 67449 629642 67515 629645
rect 61837 629640 67515 629642
rect 61837 629584 61842 629640
rect 61898 629584 67454 629640
rect 67510 629584 67515 629640
rect 61837 629582 67515 629584
rect 61837 629579 61903 629582
rect 67449 629579 67515 629582
rect 68277 629642 68343 629645
rect 219433 629642 219499 629645
rect 249793 629642 249859 629645
rect 68277 629640 219499 629642
rect 68277 629584 68282 629640
rect 68338 629584 219438 629640
rect 219494 629584 219499 629640
rect 68277 629582 219499 629584
rect 68277 629579 68343 629582
rect 219433 629579 219499 629582
rect 238710 629640 249859 629642
rect 238710 629584 249798 629640
rect 249854 629584 249859 629640
rect 238710 629582 249859 629584
rect 64597 629506 64663 629509
rect 67541 629506 67607 629509
rect 225505 629506 225571 629509
rect 64597 629504 67607 629506
rect 64597 629448 64602 629504
rect 64658 629448 67546 629504
rect 67602 629448 67607 629504
rect 64597 629446 67607 629448
rect 64597 629443 64663 629446
rect 67541 629443 67607 629446
rect 67774 629504 225571 629506
rect 67774 629448 225510 629504
rect 225566 629448 225571 629504
rect 67774 629446 225571 629448
rect 65977 629370 66043 629373
rect 66897 629370 66963 629373
rect 67774 629370 67834 629446
rect 225505 629443 225571 629446
rect 238710 629370 238770 629582
rect 249793 629579 249859 629582
rect 543089 629506 543155 629509
rect 539948 629504 543155 629506
rect 539948 629448 543094 629504
rect 543150 629448 543155 629504
rect 539948 629446 543155 629448
rect 543089 629443 543155 629446
rect 65977 629368 66730 629370
rect 65977 629312 65982 629368
rect 66038 629312 66730 629368
rect 65977 629310 66730 629312
rect 65977 629307 66043 629310
rect 66670 629234 66730 629310
rect 66897 629368 67834 629370
rect 66897 629312 66902 629368
rect 66958 629312 67834 629368
rect 66897 629310 67834 629312
rect 67958 629310 238770 629370
rect 66897 629307 66963 629310
rect 67958 629234 68018 629310
rect 66670 629174 68018 629234
rect 539918 627877 539978 628116
rect 539869 627872 539978 627877
rect 539869 627816 539874 627872
rect 539930 627816 539978 627872
rect 539869 627814 539978 627816
rect 539869 627811 539935 627814
rect 545297 626786 545363 626789
rect 539948 626784 545363 626786
rect 539948 626728 545302 626784
rect 545358 626728 545363 626784
rect 539948 626726 545363 626728
rect 545297 626723 545363 626726
rect 68502 626588 68508 626652
rect 68572 626650 68578 626652
rect 68572 626590 70196 626650
rect 68572 626588 68578 626590
rect 291142 626378 291148 626380
rect 289892 626318 291148 626378
rect 291142 626316 291148 626318
rect 291212 626316 291218 626380
rect 540053 625562 540119 625565
rect 539918 625560 540119 625562
rect 539918 625504 540058 625560
rect 540114 625504 540119 625560
rect 539918 625502 540119 625504
rect 539918 625396 539978 625502
rect 540053 625499 540119 625502
rect 544101 624066 544167 624069
rect 539948 624064 544167 624066
rect 539948 624008 544106 624064
rect 544162 624008 544167 624064
rect 539948 624006 544167 624008
rect 544101 624003 544167 624006
rect 541065 622706 541131 622709
rect 539948 622704 541131 622706
rect 539948 622648 541070 622704
rect 541126 622648 541131 622704
rect 539948 622646 541131 622648
rect 541065 622643 541131 622646
rect 68686 622236 68692 622300
rect 68756 622298 68762 622300
rect 290590 622298 290596 622300
rect 68756 622238 70196 622298
rect 289892 622238 290596 622298
rect 68756 622236 68762 622238
rect 290590 622236 290596 622238
rect 290660 622236 290666 622300
rect 541157 621346 541223 621349
rect 539948 621344 541223 621346
rect 539948 621288 541162 621344
rect 541218 621288 541223 621344
rect 539948 621286 541223 621288
rect 541157 621283 541223 621286
rect 544009 619986 544075 619989
rect 539948 619984 544075 619986
rect 539948 619928 544014 619984
rect 544070 619928 544075 619984
rect 539948 619926 544075 619928
rect 544009 619923 544075 619926
rect -960 619170 480 619260
rect 2998 619170 3004 619172
rect -960 619110 3004 619170
rect -960 619020 480 619110
rect 2998 619108 3004 619110
rect 3068 619108 3074 619172
rect 541014 618626 541020 618628
rect 539948 618566 541020 618626
rect 541014 618564 541020 618566
rect 541084 618564 541090 618628
rect 291694 618218 291700 618220
rect 289892 618158 291700 618218
rect 291694 618156 291700 618158
rect 291764 618156 291770 618220
rect 68870 617884 68876 617948
rect 68940 617946 68946 617948
rect 68940 617886 70196 617946
rect 68940 617884 68946 617886
rect 580533 617538 580599 617541
rect 583520 617538 584960 617628
rect 580533 617536 584960 617538
rect 580533 617480 580538 617536
rect 580594 617480 584960 617536
rect 580533 617478 584960 617480
rect 580533 617475 580599 617478
rect 583520 617388 584960 617478
rect 544193 617266 544259 617269
rect 539948 617264 544259 617266
rect 539948 617208 544198 617264
rect 544254 617208 544259 617264
rect 539948 617206 544259 617208
rect 544193 617203 544259 617206
rect 542445 615906 542511 615909
rect 539948 615904 542511 615906
rect 539948 615848 542450 615904
rect 542506 615848 542511 615904
rect 539948 615846 542511 615848
rect 542445 615843 542511 615846
rect 542905 614546 542971 614549
rect 539948 614544 542971 614546
rect 539948 614488 542910 614544
rect 542966 614488 542971 614544
rect 539948 614486 542971 614488
rect 542905 614483 542971 614486
rect 291510 614138 291516 614140
rect 289892 614078 291516 614138
rect 291510 614076 291516 614078
rect 291580 614076 291586 614140
rect 487797 613730 487863 613733
rect 487797 613728 490084 613730
rect 487797 613672 487802 613728
rect 487858 613672 490084 613728
rect 487797 613670 490084 613672
rect 487797 613667 487863 613670
rect 70158 613532 70164 613596
rect 70228 613532 70234 613596
rect 542353 613186 542419 613189
rect 539948 613184 542419 613186
rect 539948 613128 542358 613184
rect 542414 613128 542419 613184
rect 539948 613126 542419 613128
rect 542353 613123 542419 613126
rect 543181 611826 543247 611829
rect 539948 611824 543247 611826
rect 539948 611768 543186 611824
rect 543242 611768 543247 611824
rect 539948 611766 543247 611768
rect 543181 611763 543247 611766
rect 542537 610466 542603 610469
rect 539948 610464 542603 610466
rect 539948 610408 542542 610464
rect 542598 610408 542603 610464
rect 539948 610406 542603 610408
rect 542537 610403 542603 610406
rect 291326 610058 291332 610060
rect 289892 609998 291332 610058
rect 291326 609996 291332 609998
rect 291396 609996 291402 610060
rect 68134 609180 68140 609244
rect 68204 609242 68210 609244
rect 68204 609182 70196 609242
rect 68204 609180 68210 609182
rect 542813 609106 542879 609109
rect 539948 609104 542879 609106
rect 539948 609048 542818 609104
rect 542874 609048 542879 609104
rect 539948 609046 542879 609048
rect 542813 609043 542879 609046
rect 542854 607746 542860 607748
rect 539948 607686 542860 607746
rect 542854 607684 542860 607686
rect 542924 607684 542930 607748
rect 543038 606386 543044 606388
rect 539948 606326 543044 606386
rect 543038 606324 543044 606326
rect 543108 606324 543114 606388
rect -960 606114 480 606204
rect 3366 606114 3372 606116
rect -960 606054 3372 606114
rect -960 605964 480 606054
rect 3366 606052 3372 606054
rect 3436 606052 3442 606116
rect 291285 605978 291351 605981
rect 289892 605976 291351 605978
rect 289892 605920 291290 605976
rect 291346 605920 291351 605976
rect 289892 605918 291351 605920
rect 291285 605915 291351 605918
rect 543222 605026 543228 605028
rect 539948 604966 543228 605026
rect 543222 604964 543228 604966
rect 543292 604964 543298 605028
rect 68318 604828 68324 604892
rect 68388 604890 68394 604892
rect 68388 604830 70196 604890
rect 68388 604828 68394 604830
rect 68502 604420 68508 604484
rect 68572 604482 68578 604484
rect 68737 604482 68803 604485
rect 68572 604480 68803 604482
rect 68572 604424 68742 604480
rect 68798 604424 68803 604480
rect 68572 604422 68803 604424
rect 68572 604420 68578 604422
rect 68737 604419 68803 604422
rect 583520 604060 584960 604300
rect 539358 603604 539364 603668
rect 539428 603604 539434 603668
rect 291929 601898 291995 601901
rect 289892 601896 291995 601898
rect 289892 601840 291934 601896
rect 291990 601840 291995 601896
rect 289892 601838 291995 601840
rect 291929 601835 291995 601838
rect 68645 601084 68711 601085
rect 68645 601082 68692 601084
rect 68600 601080 68692 601082
rect 68600 601024 68650 601080
rect 68600 601022 68692 601024
rect 68645 601020 68692 601022
rect 68756 601020 68762 601084
rect 68645 601019 68711 601020
rect 68502 600476 68508 600540
rect 68572 600538 68578 600540
rect 68572 600478 70196 600538
rect 68572 600476 68578 600478
rect 300117 598226 300183 598229
rect 530761 598226 530827 598229
rect 300117 598224 530827 598226
rect 300117 598168 300122 598224
rect 300178 598168 530766 598224
rect 530822 598168 530827 598224
rect 300117 598166 530827 598168
rect 300117 598163 300183 598166
rect 530761 598163 530827 598166
rect 291469 597818 291535 597821
rect 289892 597816 291535 597818
rect 289892 597760 291474 597816
rect 291530 597760 291535 597816
rect 289892 597758 291535 597760
rect 291469 597755 291535 597758
rect 69606 596124 69612 596188
rect 69676 596186 69682 596188
rect 69676 596126 70196 596186
rect 69676 596124 69682 596126
rect 291377 593738 291443 593741
rect 289892 593736 291443 593738
rect 289892 593680 291382 593736
rect 291438 593680 291443 593736
rect 289892 593678 291443 593680
rect 291377 593675 291443 593678
rect -960 592908 480 593148
rect 63350 591772 63356 591836
rect 63420 591834 63426 591836
rect 63420 591774 70196 591834
rect 63420 591772 63426 591774
rect 306966 591228 306972 591292
rect 307036 591290 307042 591292
rect 580206 591290 580212 591292
rect 307036 591230 580212 591290
rect 307036 591228 307042 591230
rect 580206 591228 580212 591230
rect 580276 591228 580282 591292
rect 580533 591018 580599 591021
rect 583520 591018 584960 591108
rect 580533 591016 584960 591018
rect 580533 590960 580538 591016
rect 580594 590960 584960 591016
rect 580533 590958 584960 590960
rect 580533 590955 580599 590958
rect 583520 590868 584960 590958
rect 291561 589658 291627 589661
rect 289892 589656 291627 589658
rect 289892 589600 291566 589656
rect 291622 589600 291627 589656
rect 289892 589598 291627 589600
rect 291561 589595 291627 589598
rect 63166 587420 63172 587484
rect 63236 587482 63242 587484
rect 63236 587422 70196 587482
rect 63236 587420 63242 587422
rect 291653 585578 291719 585581
rect 289892 585576 291719 585578
rect 289892 585520 291658 585576
rect 291714 585520 291719 585576
rect 289892 585518 291719 585520
rect 291653 585515 291719 585518
rect 69974 582524 69980 582588
rect 70044 582586 70050 582588
rect 70166 582586 70226 583100
rect 70044 582526 70226 582586
rect 70044 582524 70050 582526
rect 290774 581498 290780 581500
rect 289892 581438 290780 581498
rect 290774 581436 290780 581438
rect 290844 581436 290850 581500
rect -960 580002 480 580092
rect 60549 580002 60615 580005
rect -960 580000 60615 580002
rect -960 579944 60554 580000
rect 60610 579944 60615 580000
rect -960 579942 60615 579944
rect -960 579852 480 579942
rect 60549 579939 60615 579942
rect 60549 579594 60615 579597
rect 68277 579594 68343 579597
rect 60549 579592 68343 579594
rect 60549 579536 60554 579592
rect 60610 579536 68282 579592
rect 68338 579536 68343 579592
rect 60549 579534 68343 579536
rect 60549 579531 60615 579534
rect 68277 579531 68343 579534
rect 69422 578716 69428 578780
rect 69492 578778 69498 578780
rect 69492 578718 70196 578778
rect 69492 578716 69498 578718
rect 313774 577628 313780 577692
rect 313844 577690 313850 577692
rect 583520 577690 584960 577780
rect 313844 577630 584960 577690
rect 313844 577628 313850 577630
rect 583520 577540 584960 577630
rect 291745 577418 291811 577421
rect 289892 577416 291811 577418
rect 289892 577360 291750 577416
rect 291806 577360 291811 577416
rect 289892 577358 291811 577360
rect 291745 577355 291811 577358
rect 66846 574364 66852 574428
rect 66916 574426 66922 574428
rect 66916 574366 70196 574426
rect 66916 574364 66922 574366
rect 296713 573338 296779 573341
rect 289892 573336 296779 573338
rect 289892 573280 296718 573336
rect 296774 573280 296779 573336
rect 289892 573278 296779 573280
rect 296713 573275 296779 573278
rect 69565 571298 69631 571301
rect 70158 571298 70164 571300
rect 69565 571296 70164 571298
rect 69565 571240 69570 571296
rect 69626 571240 70164 571296
rect 69565 571238 70164 571240
rect 69565 571235 69631 571238
rect 70158 571236 70164 571238
rect 70228 571236 70234 571300
rect 69790 570012 69796 570076
rect 69860 570074 69866 570076
rect 69860 570014 70196 570074
rect 69860 570012 69866 570014
rect 295425 569258 295491 569261
rect 289892 569256 295491 569258
rect 289892 569200 295430 569256
rect 295486 569200 295491 569256
rect 289892 569198 295491 569200
rect 295425 569195 295491 569198
rect -960 566946 480 567036
rect 3550 566946 3556 566948
rect -960 566886 3556 566946
rect -960 566796 480 566886
rect 3550 566884 3556 566886
rect 3620 566884 3626 566948
rect 65558 565660 65564 565724
rect 65628 565722 65634 565724
rect 65628 565662 70196 565722
rect 65628 565660 65634 565662
rect 289862 564501 289922 565148
rect 289862 564496 289971 564501
rect 289862 564440 289910 564496
rect 289966 564440 289971 564496
rect 289862 564438 289971 564440
rect 289905 564435 289971 564438
rect 580625 564362 580691 564365
rect 583520 564362 584960 564452
rect 580625 564360 584960 564362
rect 580625 564304 580630 564360
rect 580686 564304 584960 564360
rect 580625 564302 584960 564304
rect 580625 564299 580691 564302
rect 583520 564212 584960 564302
rect 67398 561308 67404 561372
rect 67468 561370 67474 561372
rect 67468 561310 70196 561370
rect 67468 561308 67474 561310
rect 296805 561098 296871 561101
rect 289892 561096 296871 561098
rect 289892 561040 296810 561096
rect 296866 561040 296871 561096
rect 289892 561038 296871 561040
rect 296805 561035 296871 561038
rect 67214 556956 67220 557020
rect 67284 557018 67290 557020
rect 67284 556958 70196 557018
rect 67284 556956 67290 556958
rect 289862 556202 289922 556988
rect 289997 556202 290063 556205
rect 289862 556200 290063 556202
rect 289862 556144 290002 556200
rect 290058 556144 290063 556200
rect 289862 556142 290063 556144
rect 289997 556139 290063 556142
rect -960 553890 480 553980
rect 3734 553890 3740 553892
rect -960 553830 3740 553890
rect -960 553740 480 553830
rect 3734 553828 3740 553830
rect 3804 553828 3810 553892
rect 2998 553420 3004 553484
rect 3068 553482 3074 553484
rect 4061 553482 4127 553485
rect 3068 553480 4127 553482
rect 3068 553424 4066 553480
rect 4122 553424 4127 553480
rect 3068 553422 4127 553424
rect 3068 553420 3074 553422
rect 4061 553419 4127 553422
rect 66110 552604 66116 552668
rect 66180 552666 66186 552668
rect 66180 552606 70196 552666
rect 66180 552604 66186 552606
rect 289862 552397 289922 552908
rect 289813 552392 289922 552397
rect 289813 552336 289818 552392
rect 289874 552336 289922 552392
rect 289813 552334 289922 552336
rect 289813 552331 289879 552334
rect 583520 551020 584960 551260
rect 290089 548858 290155 548861
rect 289892 548856 290155 548858
rect 289892 548800 290094 548856
rect 290150 548800 290155 548856
rect 289892 548798 290155 548800
rect 290089 548795 290155 548798
rect 67030 548252 67036 548316
rect 67100 548314 67106 548316
rect 67100 548254 70196 548314
rect 67100 548252 67106 548254
rect 290365 544778 290431 544781
rect 289892 544776 290431 544778
rect 289892 544720 290370 544776
rect 290426 544720 290431 544776
rect 289892 544718 290431 544720
rect 290365 544715 290431 544718
rect 65926 543900 65932 543964
rect 65996 543962 66002 543964
rect 65996 543902 70196 543962
rect 65996 543900 66002 543902
rect -960 540684 480 540924
rect 66846 540908 66852 540972
rect 66916 540970 66922 540972
rect 67449 540970 67515 540973
rect 66916 540968 67515 540970
rect 66916 540912 67454 540968
rect 67510 540912 67515 540968
rect 66916 540910 67515 540912
rect 66916 540908 66922 540910
rect 67449 540907 67515 540910
rect 290273 540698 290339 540701
rect 289892 540696 290339 540698
rect 289892 540640 290278 540696
rect 290334 540640 290339 540696
rect 289892 540638 290339 540640
rect 290273 540635 290339 540638
rect 66846 539548 66852 539612
rect 66916 539610 66922 539612
rect 66916 539550 70196 539610
rect 66916 539548 66922 539550
rect 580625 537842 580691 537845
rect 583520 537842 584960 537932
rect 580625 537840 584960 537842
rect 580625 537784 580630 537840
rect 580686 537784 584960 537840
rect 580625 537782 584960 537784
rect 580625 537779 580691 537782
rect 583520 537692 584960 537782
rect 290181 536618 290247 536621
rect 289892 536616 290247 536618
rect 289892 536560 290186 536616
rect 290242 536560 290247 536616
rect 289892 536558 290247 536560
rect 290181 536555 290247 536558
rect 65742 535196 65748 535260
rect 65812 535258 65818 535260
rect 65812 535198 70196 535258
rect 65812 535196 65818 535198
rect 290457 532538 290523 532541
rect 289892 532536 290523 532538
rect 289892 532480 290462 532536
rect 290518 532480 290523 532536
rect 289892 532478 290523 532480
rect 290457 532475 290523 532478
rect 68093 531314 68159 531317
rect 68870 531314 68876 531316
rect 68093 531312 68876 531314
rect 68093 531256 68098 531312
rect 68154 531256 68876 531312
rect 68093 531254 68876 531256
rect 68093 531251 68159 531254
rect 68870 531252 68876 531254
rect 68940 531252 68946 531316
rect 68686 530844 68692 530908
rect 68756 530906 68762 530908
rect 68756 530846 70196 530906
rect 68756 530844 68762 530846
rect 294413 528458 294479 528461
rect 289892 528456 294479 528458
rect 289892 528400 294418 528456
rect 294474 528400 294479 528456
rect 289892 528398 294479 528400
rect 294413 528395 294479 528398
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 60733 527234 60799 527237
rect 61745 527234 61811 527237
rect 66897 527234 66963 527237
rect 60733 527232 66963 527234
rect 60733 527176 60738 527232
rect 60794 527176 61750 527232
rect 61806 527176 66902 527232
rect 66958 527176 66963 527232
rect 60733 527174 66963 527176
rect 60733 527171 60799 527174
rect 61745 527171 61811 527174
rect 66897 527171 66963 527174
rect 68870 526492 68876 526556
rect 68940 526554 68946 526556
rect 68940 526494 70196 526554
rect 68940 526492 68946 526494
rect 68134 525812 68140 525876
rect 68204 525874 68210 525876
rect 68461 525874 68527 525877
rect 68204 525872 68527 525874
rect 68204 525816 68466 525872
rect 68522 525816 68527 525872
rect 68204 525814 68527 525816
rect 68204 525812 68210 525814
rect 68461 525811 68527 525814
rect 309726 524452 309732 524516
rect 309796 524514 309802 524516
rect 583520 524514 584960 524604
rect 309796 524454 584960 524514
rect 309796 524452 309802 524454
rect 293125 524378 293191 524381
rect 289892 524376 293191 524378
rect 289892 524320 293130 524376
rect 293186 524320 293191 524376
rect 583520 524364 584960 524454
rect 289892 524318 293191 524320
rect 293125 524315 293191 524318
rect 67909 523018 67975 523021
rect 68318 523018 68324 523020
rect 67909 523016 68324 523018
rect 67909 522960 67914 523016
rect 67970 522960 68324 523016
rect 67909 522958 68324 522960
rect 67909 522955 67975 522958
rect 68318 522956 68324 522958
rect 68388 522956 68394 523020
rect 67950 522140 67956 522204
rect 68020 522202 68026 522204
rect 68020 522142 70196 522202
rect 68020 522140 68026 522142
rect 291837 520298 291903 520301
rect 289892 520296 291903 520298
rect 289892 520240 291842 520296
rect 291898 520240 291903 520296
rect 289892 520238 291903 520240
rect 291837 520235 291903 520238
rect 68134 517788 68140 517852
rect 68204 517850 68210 517852
rect 68204 517790 70196 517850
rect 68204 517788 68210 517790
rect 68185 517578 68251 517581
rect 68502 517578 68508 517580
rect 68185 517576 68508 517578
rect 68185 517520 68190 517576
rect 68246 517520 68508 517576
rect 68185 517518 68508 517520
rect 68185 517515 68251 517518
rect 68502 517516 68508 517518
rect 68572 517516 68578 517580
rect 289302 516156 289308 516220
rect 289372 516156 289378 516220
rect -960 514858 480 514948
rect 59854 514858 59860 514860
rect -960 514798 59860 514858
rect -960 514708 480 514798
rect 59854 514796 59860 514798
rect 59924 514796 59930 514860
rect 68686 513980 68692 514044
rect 68756 514042 68762 514044
rect 68829 514042 68895 514045
rect 68756 514040 68895 514042
rect 68756 513984 68834 514040
rect 68890 513984 68895 514040
rect 68756 513982 68895 513984
rect 68756 513980 68762 513982
rect 68829 513979 68895 513982
rect 68686 513436 68692 513500
rect 68756 513498 68762 513500
rect 68756 513438 70196 513498
rect 68756 513436 68762 513438
rect 291193 512138 291259 512141
rect 289892 512136 291259 512138
rect 289892 512080 291198 512136
rect 291254 512080 291259 512136
rect 289892 512078 291259 512080
rect 291193 512075 291259 512078
rect 580441 511322 580507 511325
rect 583520 511322 584960 511412
rect 580441 511320 584960 511322
rect 580441 511264 580446 511320
rect 580502 511264 584960 511320
rect 580441 511262 584960 511264
rect 580441 511259 580507 511262
rect 583520 511172 584960 511262
rect 68502 509084 68508 509148
rect 68572 509146 68578 509148
rect 68572 509086 70196 509146
rect 68572 509084 68578 509086
rect 289310 507925 289370 508028
rect 68277 507922 68343 507925
rect 68870 507922 68876 507924
rect 68277 507920 68876 507922
rect 68277 507864 68282 507920
rect 68338 507864 68876 507920
rect 68277 507862 68876 507864
rect 68277 507859 68343 507862
rect 68870 507860 68876 507862
rect 68940 507860 68946 507924
rect 289310 507920 289419 507925
rect 289310 507864 289358 507920
rect 289414 507864 289419 507920
rect 289310 507862 289419 507864
rect 289353 507859 289419 507862
rect 62982 504732 62988 504796
rect 63052 504794 63058 504796
rect 63052 504734 70196 504794
rect 63052 504732 63058 504734
rect 292021 503978 292087 503981
rect 289892 503976 292087 503978
rect 289892 503920 292026 503976
rect 292082 503920 292087 503976
rect 289892 503918 292087 503920
rect 292021 503915 292087 503918
rect 2814 502284 2820 502348
rect 2884 502346 2890 502348
rect 3969 502346 4035 502349
rect 2884 502344 4035 502346
rect 2884 502288 3974 502344
rect 4030 502288 4035 502344
rect 2884 502286 4035 502288
rect 2884 502284 2890 502286
rect 3969 502283 4035 502286
rect -960 501802 480 501892
rect 3918 501802 3924 501804
rect -960 501742 3924 501802
rect -960 501652 480 501742
rect 3918 501740 3924 501742
rect 3988 501740 3994 501804
rect 67950 500788 67956 500852
rect 68020 500850 68026 500852
rect 68553 500850 68619 500853
rect 68020 500848 68619 500850
rect 68020 500792 68558 500848
rect 68614 500792 68619 500848
rect 68020 500790 68619 500792
rect 68020 500788 68026 500790
rect 68553 500787 68619 500790
rect 68318 500380 68324 500444
rect 68388 500442 68394 500444
rect 68388 500382 70196 500442
rect 68388 500380 68394 500382
rect 289494 499765 289554 499868
rect 289494 499760 289603 499765
rect 289494 499704 289542 499760
rect 289598 499704 289603 499760
rect 289494 499702 289603 499704
rect 289537 499699 289603 499702
rect 583520 497844 584960 498084
rect 69606 496300 69612 496364
rect 69676 496362 69682 496364
rect 70117 496362 70183 496365
rect 69676 496360 70183 496362
rect 69676 496304 70122 496360
rect 70178 496304 70183 496360
rect 69676 496302 70183 496304
rect 69676 496300 69682 496302
rect 70117 496299 70183 496302
rect 69606 496028 69612 496092
rect 69676 496090 69682 496092
rect 69676 496030 70196 496090
rect 69676 496028 69682 496030
rect 289862 495546 289922 495788
rect 289862 495486 291394 495546
rect 291193 495410 291259 495413
rect 291334 495410 291394 495486
rect 291193 495408 291394 495410
rect 291193 495352 291198 495408
rect 291254 495352 291394 495408
rect 291193 495350 291394 495352
rect 291193 495347 291259 495350
rect 65558 492628 65564 492692
rect 65628 492690 65634 492692
rect 65793 492690 65859 492693
rect 65628 492688 65859 492690
rect 65628 492632 65798 492688
rect 65854 492632 65859 492688
rect 65628 492630 65859 492632
rect 65628 492628 65634 492630
rect 65793 492627 65859 492630
rect 65558 491676 65564 491740
rect 65628 491738 65634 491740
rect 65628 491678 70196 491738
rect 65628 491676 65634 491678
rect 289494 491333 289554 491708
rect 289445 491328 289554 491333
rect 289445 491272 289450 491328
rect 289506 491272 289554 491328
rect 289445 491270 289554 491272
rect 289445 491267 289511 491270
rect -960 488596 480 488836
rect 290641 487658 290707 487661
rect 289892 487656 290707 487658
rect 289892 487600 290646 487656
rect 290702 487600 290707 487656
rect 289892 487598 290707 487600
rect 290641 487595 290707 487598
rect 69749 487386 69815 487389
rect 69749 487384 70196 487386
rect 69749 487328 69754 487384
rect 69810 487328 70196 487384
rect 69749 487326 70196 487328
rect 69749 487323 69815 487326
rect 580206 484604 580212 484668
rect 580276 484666 580282 484668
rect 583520 484666 584960 484756
rect 580276 484606 584960 484666
rect 580276 484604 580282 484606
rect 583520 484516 584960 484606
rect 294505 483578 294571 483581
rect 289892 483576 294571 483578
rect 289892 483520 294510 483576
rect 294566 483520 294571 483576
rect 289892 483518 294571 483520
rect 294505 483515 294571 483518
rect 68921 483034 68987 483037
rect 68921 483032 70196 483034
rect 68921 482976 68926 483032
rect 68982 482976 70196 483032
rect 68921 482974 70196 482976
rect 68921 482971 68987 482974
rect 289629 481538 289695 481541
rect 291285 481538 291351 481541
rect 289629 481536 291351 481538
rect 289629 481480 289634 481536
rect 289690 481480 291290 481536
rect 291346 481480 291351 481536
rect 289629 481478 291351 481480
rect 289629 481475 289695 481478
rect 291285 481475 291351 481478
rect 289445 481130 289511 481133
rect 291694 481130 291700 481132
rect 289445 481128 291700 481130
rect 289445 481072 289450 481128
rect 289506 481072 291700 481128
rect 289445 481070 291700 481072
rect 289445 481067 289511 481070
rect 291694 481068 291700 481070
rect 291764 481068 291770 481132
rect 288985 480314 289051 480317
rect 291469 480314 291535 480317
rect 288985 480312 291535 480314
rect 288985 480256 288990 480312
rect 289046 480256 291474 480312
rect 291530 480256 291535 480312
rect 288985 480254 291535 480256
rect 288985 480251 289051 480254
rect 291469 480251 291535 480254
rect 278221 480178 278287 480181
rect 290590 480178 290596 480180
rect 278221 480176 290596 480178
rect 278221 480120 278226 480176
rect 278282 480120 290596 480176
rect 278221 480118 290596 480120
rect 278221 480115 278287 480118
rect 290590 480116 290596 480118
rect 290660 480116 290666 480180
rect 268101 480042 268167 480045
rect 290774 480042 290780 480044
rect 268101 480040 290780 480042
rect 268101 479984 268106 480040
rect 268162 479984 290780 480040
rect 268101 479982 290780 479984
rect 268101 479979 268167 479982
rect 290774 479980 290780 479982
rect 290844 479980 290850 480044
rect 264053 479906 264119 479909
rect 289905 479906 289971 479909
rect 264053 479904 289971 479906
rect 264053 479848 264058 479904
rect 264114 479848 289910 479904
rect 289966 479848 289971 479904
rect 264053 479846 289971 479848
rect 264053 479843 264119 479846
rect 289905 479843 289971 479846
rect 244825 479770 244891 479773
rect 290641 479770 290707 479773
rect 244825 479768 290707 479770
rect 244825 479712 244830 479768
rect 244886 479712 290646 479768
rect 290702 479712 290707 479768
rect 244825 479710 290707 479712
rect 244825 479707 244891 479710
rect 290641 479707 290707 479710
rect 234521 479634 234587 479637
rect 543089 479634 543155 479637
rect 234521 479632 543155 479634
rect 234521 479576 234526 479632
rect 234582 479576 543094 479632
rect 543150 479576 543155 479632
rect 234521 479574 543155 479576
rect 234521 479571 234587 479574
rect 543089 479571 543155 479574
rect 68185 479498 68251 479501
rect 123477 479498 123543 479501
rect 68185 479496 123543 479498
rect 68185 479440 68190 479496
rect 68246 479440 123482 479496
rect 123538 479440 123543 479496
rect 68185 479438 123543 479440
rect 68185 479435 68251 479438
rect 123477 479435 123543 479438
rect 234470 479436 234476 479500
rect 234540 479498 234546 479500
rect 543222 479498 543228 479500
rect 234540 479438 543228 479498
rect 234540 479436 234546 479438
rect 543222 479436 543228 479438
rect 543292 479436 543298 479500
rect 231209 478818 231275 478821
rect 243721 478818 243787 478821
rect 231209 478816 243787 478818
rect 231209 478760 231214 478816
rect 231270 478760 243726 478816
rect 243782 478760 243787 478816
rect 231209 478758 243787 478760
rect 231209 478755 231275 478758
rect 243721 478755 243787 478758
rect 267089 478818 267155 478821
rect 291745 478818 291811 478821
rect 267089 478816 291811 478818
rect 267089 478760 267094 478816
rect 267150 478760 291750 478816
rect 291806 478760 291811 478816
rect 267089 478758 291811 478760
rect 267089 478755 267155 478758
rect 291745 478755 291811 478758
rect 67357 478682 67423 478685
rect 79133 478682 79199 478685
rect 67357 478680 79199 478682
rect 67357 478624 67362 478680
rect 67418 478624 79138 478680
rect 79194 478624 79199 478680
rect 67357 478622 79199 478624
rect 67357 478619 67423 478622
rect 79133 478619 79199 478622
rect 228449 478682 228515 478685
rect 255865 478682 255931 478685
rect 228449 478680 255931 478682
rect 228449 478624 228454 478680
rect 228510 478624 255870 478680
rect 255926 478624 255931 478680
rect 228449 478622 255931 478624
rect 228449 478619 228515 478622
rect 255865 478619 255931 478622
rect 262029 478682 262095 478685
rect 289997 478682 290063 478685
rect 262029 478680 290063 478682
rect 262029 478624 262034 478680
rect 262090 478624 290002 478680
rect 290058 478624 290063 478680
rect 262029 478622 290063 478624
rect 262029 478619 262095 478622
rect 289997 478619 290063 478622
rect 69749 478546 69815 478549
rect 241789 478546 241855 478549
rect 69749 478544 241855 478546
rect 69749 478488 69754 478544
rect 69810 478488 241794 478544
rect 241850 478488 241855 478544
rect 69749 478486 241855 478488
rect 69749 478483 69815 478486
rect 241789 478483 241855 478486
rect 258993 478546 259059 478549
rect 290365 478546 290431 478549
rect 258993 478544 290431 478546
rect 258993 478488 258998 478544
rect 259054 478488 290370 478544
rect 290426 478488 290431 478544
rect 258993 478486 290431 478488
rect 258993 478483 259059 478486
rect 290365 478483 290431 478486
rect 69841 478410 69907 478413
rect 84101 478410 84167 478413
rect 69841 478408 84167 478410
rect 69841 478352 69846 478408
rect 69902 478352 84106 478408
rect 84162 478352 84167 478408
rect 69841 478350 84167 478352
rect 69841 478347 69907 478350
rect 84101 478347 84167 478350
rect 104157 478410 104223 478413
rect 292941 478410 293007 478413
rect 104157 478408 293007 478410
rect 104157 478352 104162 478408
rect 104218 478352 292946 478408
rect 293002 478352 293007 478408
rect 104157 478350 293007 478352
rect 104157 478347 104223 478350
rect 292941 478347 293007 478350
rect 69933 478274 69999 478277
rect 99373 478274 99439 478277
rect 69933 478272 99439 478274
rect 69933 478216 69938 478272
rect 69994 478216 99378 478272
rect 99434 478216 99439 478272
rect 69933 478214 99439 478216
rect 69933 478211 69999 478214
rect 99373 478211 99439 478214
rect 102317 478274 102383 478277
rect 294229 478274 294295 478277
rect 102317 478272 294295 478274
rect 102317 478216 102322 478272
rect 102378 478216 294234 478272
rect 294290 478216 294295 478272
rect 102317 478214 294295 478216
rect 102317 478211 102383 478214
rect 294229 478211 294295 478214
rect 65977 478138 66043 478141
rect 99005 478138 99071 478141
rect 65977 478136 99071 478138
rect 65977 478080 65982 478136
rect 66038 478080 99010 478136
rect 99066 478080 99071 478136
rect 65977 478078 99071 478080
rect 65977 478075 66043 478078
rect 99005 478075 99071 478078
rect 232262 478076 232268 478140
rect 232332 478138 232338 478140
rect 580206 478138 580212 478140
rect 232332 478078 580212 478138
rect 232332 478076 232338 478078
rect 580206 478076 580212 478078
rect 580276 478076 580282 478140
rect 105537 478002 105603 478005
rect 241421 478002 241487 478005
rect 249793 478002 249859 478005
rect 105537 478000 241487 478002
rect 105537 477944 105542 478000
rect 105598 477944 241426 478000
rect 241482 477944 241487 478000
rect 105537 477942 241487 477944
rect 105537 477939 105603 477942
rect 241421 477939 241487 477942
rect 248370 478000 249859 478002
rect 248370 477944 249798 478000
rect 249854 477944 249859 478000
rect 248370 477942 249859 477944
rect 66069 477866 66135 477869
rect 75821 477866 75887 477869
rect 66069 477864 75887 477866
rect 66069 477808 66074 477864
rect 66130 477808 75826 477864
rect 75882 477808 75887 477864
rect 66069 477806 75887 477808
rect 66069 477803 66135 477806
rect 75821 477803 75887 477806
rect 108297 477866 108363 477869
rect 231761 477866 231827 477869
rect 108297 477864 231827 477866
rect 108297 477808 108302 477864
rect 108358 477808 231766 477864
rect 231822 477808 231827 477864
rect 108297 477806 231827 477808
rect 108297 477803 108363 477806
rect 231761 477803 231827 477806
rect 240910 477804 240916 477868
rect 240980 477866 240986 477868
rect 248370 477866 248430 477942
rect 249793 477939 249859 477942
rect 276197 478002 276263 478005
rect 291510 478002 291516 478004
rect 276197 478000 291516 478002
rect 276197 477944 276202 478000
rect 276258 477944 291516 478000
rect 276197 477942 291516 477944
rect 276197 477939 276263 477942
rect 291510 477940 291516 477942
rect 291580 477940 291586 478004
rect 240980 477806 248430 477866
rect 240980 477804 240986 477806
rect 106917 477730 106983 477733
rect 233141 477730 233207 477733
rect 106917 477728 233207 477730
rect 106917 477672 106922 477728
rect 106978 477672 233146 477728
rect 233202 477672 233207 477728
rect 106917 477670 233207 477672
rect 106917 477667 106983 477670
rect 233141 477667 233207 477670
rect 70025 477594 70091 477597
rect 72509 477594 72575 477597
rect 70025 477592 72575 477594
rect 70025 477536 70030 477592
rect 70086 477536 72514 477592
rect 72570 477536 72575 477592
rect 70025 477534 72575 477536
rect 70025 477531 70091 477534
rect 72509 477531 72575 477534
rect 224769 477594 224835 477597
rect 227713 477594 227779 477597
rect 224769 477592 227779 477594
rect 224769 477536 224774 477592
rect 224830 477536 227718 477592
rect 227774 477536 227779 477592
rect 224769 477534 227779 477536
rect 224769 477531 224835 477534
rect 227713 477531 227779 477534
rect 271229 477050 271295 477053
rect 291561 477050 291627 477053
rect 271229 477048 291627 477050
rect 271229 476992 271234 477048
rect 271290 476992 291566 477048
rect 291622 476992 291627 477048
rect 271229 476990 291627 476992
rect 271229 476987 271295 476990
rect 291561 476987 291627 476990
rect 68318 476852 68324 476916
rect 68388 476914 68394 476916
rect 203374 476914 203380 476916
rect 68388 476854 203380 476914
rect 68388 476852 68394 476854
rect 203374 476852 203380 476854
rect 203444 476852 203450 476916
rect 260005 476914 260071 476917
rect 290089 476914 290155 476917
rect 260005 476912 290155 476914
rect 260005 476856 260010 476912
rect 260066 476856 290094 476912
rect 290150 476856 290155 476912
rect 260005 476854 290155 476856
rect 260005 476851 260071 476854
rect 290089 476851 290155 476854
rect 68645 476778 68711 476781
rect 224217 476778 224283 476781
rect 68645 476776 224283 476778
rect 68645 476720 68650 476776
rect 68706 476720 224222 476776
rect 224278 476720 224283 476776
rect 68645 476718 224283 476720
rect 68645 476715 68711 476718
rect 224217 476715 224283 476718
rect 239806 476716 239812 476780
rect 239876 476778 239882 476780
rect 542670 476778 542676 476780
rect 239876 476718 542676 476778
rect 239876 476716 239882 476718
rect 542670 476716 542676 476718
rect 542740 476716 542746 476780
rect 263041 476098 263107 476101
rect 296805 476098 296871 476101
rect 263041 476096 296871 476098
rect 263041 476040 263046 476096
rect 263102 476040 296810 476096
rect 296866 476040 296871 476096
rect 263041 476038 296871 476040
rect 263041 476035 263107 476038
rect 296805 476035 296871 476038
rect 249885 475962 249951 475965
rect 289169 475962 289235 475965
rect 249885 475960 289235 475962
rect 249885 475904 249890 475960
rect 249946 475904 289174 475960
rect 289230 475904 289235 475960
rect 249885 475902 289235 475904
rect 249885 475899 249951 475902
rect 289169 475899 289235 475902
rect 243813 475826 243879 475829
rect 294505 475826 294571 475829
rect 243813 475824 294571 475826
rect -960 475690 480 475780
rect 243813 475768 243818 475824
rect 243874 475768 294510 475824
rect 294566 475768 294571 475824
rect 243813 475766 294571 475768
rect 243813 475763 243879 475766
rect 294505 475763 294571 475766
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 227621 475690 227687 475693
rect 292849 475690 292915 475693
rect 227621 475688 292915 475690
rect 227621 475632 227626 475688
rect 227682 475632 292854 475688
rect 292910 475632 292915 475688
rect 227621 475630 292915 475632
rect 227621 475627 227687 475630
rect 292849 475627 292915 475630
rect 231485 475554 231551 475557
rect 490741 475554 490807 475557
rect 231485 475552 490807 475554
rect 231485 475496 231490 475552
rect 231546 475496 490746 475552
rect 490802 475496 490807 475552
rect 231485 475494 490807 475496
rect 231485 475491 231551 475494
rect 490741 475491 490807 475494
rect 68737 475418 68803 475421
rect 214649 475418 214715 475421
rect 68737 475416 214715 475418
rect 68737 475360 68742 475416
rect 68798 475360 214654 475416
rect 214710 475360 214715 475416
rect 68737 475358 214715 475360
rect 68737 475355 68803 475358
rect 214649 475355 214715 475358
rect 230381 475418 230447 475421
rect 231853 475418 231919 475421
rect 230381 475416 231919 475418
rect 230381 475360 230386 475416
rect 230442 475360 231858 475416
rect 231914 475360 231919 475416
rect 230381 475358 231919 475360
rect 230381 475355 230447 475358
rect 231853 475355 231919 475358
rect 232865 475418 232931 475421
rect 504541 475418 504607 475421
rect 232865 475416 504607 475418
rect 232865 475360 232870 475416
rect 232926 475360 504546 475416
rect 504602 475360 504607 475416
rect 232865 475358 504607 475360
rect 232865 475355 232931 475358
rect 504541 475355 504607 475358
rect 228173 475282 228239 475285
rect 233877 475282 233943 475285
rect 228173 475280 233943 475282
rect 228173 475224 228178 475280
rect 228234 475224 233882 475280
rect 233938 475224 233943 475280
rect 228173 475222 233943 475224
rect 228173 475219 228239 475222
rect 233877 475219 233943 475222
rect 234245 475282 234311 475285
rect 243537 475282 243603 475285
rect 234245 475280 243603 475282
rect 234245 475224 234250 475280
rect 234306 475224 243542 475280
rect 243598 475224 243603 475280
rect 234245 475222 243603 475224
rect 234245 475219 234311 475222
rect 243537 475219 243603 475222
rect 271137 475282 271203 475285
rect 291377 475282 291443 475285
rect 271137 475280 291443 475282
rect 271137 475224 271142 475280
rect 271198 475224 291382 475280
rect 291438 475224 291443 475280
rect 271137 475222 291443 475224
rect 271137 475219 271203 475222
rect 291377 475219 291443 475222
rect 228817 475146 228883 475149
rect 251081 475146 251147 475149
rect 228817 475144 251147 475146
rect 228817 475088 228822 475144
rect 228878 475088 251086 475144
rect 251142 475088 251147 475144
rect 228817 475086 251147 475088
rect 228817 475083 228883 475086
rect 251081 475083 251147 475086
rect 227529 475010 227595 475013
rect 262857 475010 262923 475013
rect 227529 475008 262923 475010
rect 227529 474952 227534 475008
rect 227590 474952 262862 475008
rect 262918 474952 262923 475008
rect 227529 474950 262923 474952
rect 227529 474947 227595 474950
rect 262857 474947 262923 474950
rect 230197 474874 230263 474877
rect 271781 474874 271847 474877
rect 230197 474872 271847 474874
rect 230197 474816 230202 474872
rect 230258 474816 271786 474872
rect 271842 474816 271847 474872
rect 230197 474814 271847 474816
rect 230197 474811 230263 474814
rect 271781 474811 271847 474814
rect 269113 474466 269179 474469
rect 291653 474466 291719 474469
rect 269113 474464 291719 474466
rect 269113 474408 269118 474464
rect 269174 474408 291658 474464
rect 291714 474408 291719 474464
rect 269113 474406 291719 474408
rect 269113 474403 269179 474406
rect 291653 474403 291719 474406
rect 257981 474330 258047 474333
rect 290273 474330 290339 474333
rect 257981 474328 290339 474330
rect 257981 474272 257986 474328
rect 258042 474272 290278 474328
rect 290334 474272 290339 474328
rect 257981 474270 290339 474272
rect 257981 474267 258047 474270
rect 290273 474267 290339 474270
rect 68502 474132 68508 474196
rect 68572 474194 68578 474196
rect 166206 474194 166212 474196
rect 68572 474134 166212 474194
rect 68572 474132 68578 474134
rect 166206 474132 166212 474134
rect 166276 474132 166282 474196
rect 231301 474194 231367 474197
rect 532141 474194 532207 474197
rect 231301 474192 532207 474194
rect 231301 474136 231306 474192
rect 231362 474136 532146 474192
rect 532202 474136 532207 474192
rect 231301 474134 532207 474136
rect 231301 474131 231367 474134
rect 532141 474131 532207 474134
rect 3969 474058 4035 474061
rect 151169 474058 151235 474061
rect 3969 474056 151235 474058
rect 3969 474000 3974 474056
rect 4030 474000 151174 474056
rect 151230 474000 151235 474056
rect 3969 473998 151235 474000
rect 3969 473995 4035 473998
rect 151169 473995 151235 473998
rect 189073 474058 189139 474061
rect 215937 474058 216003 474061
rect 189073 474056 216003 474058
rect 189073 474000 189078 474056
rect 189134 474000 215942 474056
rect 215998 474000 216003 474056
rect 189073 473998 216003 474000
rect 189073 473995 189139 473998
rect 215937 473995 216003 473998
rect 234286 473996 234292 474060
rect 234356 474058 234362 474060
rect 543038 474058 543044 474060
rect 234356 473998 543044 474058
rect 234356 473996 234362 473998
rect 543038 473996 543044 473998
rect 543108 473996 543114 474060
rect 247861 473242 247927 473245
rect 289537 473242 289603 473245
rect 247861 473240 289603 473242
rect 247861 473184 247866 473240
rect 247922 473184 289542 473240
rect 289598 473184 289603 473240
rect 247861 473182 289603 473184
rect 247861 473179 247927 473182
rect 289537 473179 289603 473182
rect 227437 473106 227503 473109
rect 503161 473106 503227 473109
rect 227437 473104 503227 473106
rect 227437 473048 227442 473104
rect 227498 473048 503166 473104
rect 503222 473048 503227 473104
rect 227437 473046 503227 473048
rect 227437 473043 227503 473046
rect 503161 473043 503227 473046
rect 227345 472970 227411 472973
rect 510061 472970 510127 472973
rect 227345 472968 510127 472970
rect 227345 472912 227350 472968
rect 227406 472912 510066 472968
rect 510122 472912 510127 472968
rect 227345 472910 510127 472912
rect 227345 472907 227411 472910
rect 510061 472907 510127 472910
rect 230105 472834 230171 472837
rect 519721 472834 519787 472837
rect 230105 472832 519787 472834
rect 230105 472776 230110 472832
rect 230166 472776 519726 472832
rect 519782 472776 519787 472832
rect 230105 472774 519787 472776
rect 230105 472771 230171 472774
rect 519721 472771 519787 472774
rect 228633 472698 228699 472701
rect 523861 472698 523927 472701
rect 228633 472696 523927 472698
rect 228633 472640 228638 472696
rect 228694 472640 523866 472696
rect 523922 472640 523927 472696
rect 228633 472638 523927 472640
rect 228633 472635 228699 472638
rect 523861 472635 523927 472638
rect 3734 472500 3740 472564
rect 3804 472562 3810 472564
rect 161974 472562 161980 472564
rect 3804 472502 161980 472562
rect 3804 472500 3810 472502
rect 161974 472500 161980 472502
rect 162044 472500 162050 472564
rect 229737 472562 229803 472565
rect 487797 472562 487863 472565
rect 229737 472560 487863 472562
rect 229737 472504 229742 472560
rect 229798 472504 487802 472560
rect 487858 472504 487863 472560
rect 229737 472502 487863 472504
rect 229737 472499 229803 472502
rect 487797 472499 487863 472502
rect 224534 472364 224540 472428
rect 224604 472426 224610 472428
rect 230381 472426 230447 472429
rect 224604 472424 230447 472426
rect 224604 472368 230386 472424
rect 230442 472368 230447 472424
rect 224604 472366 230447 472368
rect 224604 472364 224610 472366
rect 230381 472363 230447 472366
rect 256049 472426 256115 472429
rect 290457 472426 290523 472429
rect 256049 472424 290523 472426
rect 256049 472368 256054 472424
rect 256110 472368 290462 472424
rect 290518 472368 290523 472424
rect 256049 472366 290523 472368
rect 256049 472363 256115 472366
rect 290457 472363 290523 472366
rect 227253 472290 227319 472293
rect 255313 472290 255379 472293
rect 227253 472288 255379 472290
rect 227253 472232 227258 472288
rect 227314 472232 255318 472288
rect 255374 472232 255379 472288
rect 227253 472230 255379 472232
rect 227253 472227 227319 472230
rect 255313 472227 255379 472230
rect 228541 472154 228607 472157
rect 247033 472154 247099 472157
rect 228541 472152 247099 472154
rect 228541 472096 228546 472152
rect 228602 472096 247038 472152
rect 247094 472096 247099 472152
rect 228541 472094 247099 472096
rect 228541 472091 228607 472094
rect 247033 472091 247099 472094
rect 224718 471956 224724 472020
rect 224788 472018 224794 472020
rect 230289 472018 230355 472021
rect 224788 472016 230355 472018
rect 224788 471960 230294 472016
rect 230350 471960 230355 472016
rect 224788 471958 230355 471960
rect 224788 471956 224794 471958
rect 230289 471955 230355 471958
rect 238334 471956 238340 472020
rect 238404 472018 238410 472020
rect 238477 472018 238543 472021
rect 238404 472016 238543 472018
rect 238404 471960 238482 472016
rect 238538 471960 238543 472016
rect 238404 471958 238543 471960
rect 238404 471956 238410 471958
rect 238477 471955 238543 471958
rect 273161 471610 273227 471613
rect 291929 471610 291995 471613
rect 273161 471608 291995 471610
rect 273161 471552 273166 471608
rect 273222 471552 291934 471608
rect 291990 471552 291995 471608
rect 273161 471550 291995 471552
rect 273161 471547 273227 471550
rect 291929 471547 291995 471550
rect 251909 471474 251975 471477
rect 289302 471474 289308 471476
rect 251909 471472 289308 471474
rect 251909 471416 251914 471472
rect 251970 471416 289308 471472
rect 251909 471414 289308 471416
rect 251909 471411 251975 471414
rect 289302 471412 289308 471414
rect 289372 471412 289378 471476
rect 574686 471412 574692 471476
rect 574756 471474 574762 471476
rect 583520 471474 584960 471564
rect 574756 471414 584960 471474
rect 574756 471412 574762 471414
rect 237097 471338 237163 471341
rect 512821 471338 512887 471341
rect 237097 471336 512887 471338
rect 237097 471280 237102 471336
rect 237158 471280 512826 471336
rect 512882 471280 512887 471336
rect 583520 471324 584960 471414
rect 237097 471278 512887 471280
rect 237097 471275 237163 471278
rect 512821 471275 512887 471278
rect 3918 471140 3924 471204
rect 3988 471202 3994 471204
rect 130326 471202 130332 471204
rect 3988 471142 130332 471202
rect 3988 471140 3994 471142
rect 130326 471140 130332 471142
rect 130396 471140 130402 471204
rect 234429 471202 234495 471205
rect 543181 471202 543247 471205
rect 234429 471200 543247 471202
rect 234429 471144 234434 471200
rect 234490 471144 543186 471200
rect 543242 471144 543247 471200
rect 234429 471142 543247 471144
rect 234429 471139 234495 471142
rect 543181 471139 543247 471142
rect 228357 470522 228423 470525
rect 545205 470522 545271 470525
rect 228357 470520 545271 470522
rect 228357 470464 228362 470520
rect 228418 470464 545210 470520
rect 545266 470464 545271 470520
rect 228357 470462 545271 470464
rect 228357 470459 228423 470462
rect 545205 470459 545271 470462
rect 226057 470386 226123 470389
rect 543917 470386 543983 470389
rect 226057 470384 543983 470386
rect 226057 470328 226062 470384
rect 226118 470328 543922 470384
rect 543978 470328 543983 470384
rect 226057 470326 543983 470328
rect 226057 470323 226123 470326
rect 543917 470323 543983 470326
rect 226241 470250 226307 470253
rect 545297 470250 545363 470253
rect 226241 470248 545363 470250
rect 226241 470192 226246 470248
rect 226302 470192 545302 470248
rect 545358 470192 545363 470248
rect 226241 470190 545363 470192
rect 226241 470187 226307 470190
rect 545297 470187 545363 470190
rect 224861 470114 224927 470117
rect 545113 470114 545179 470117
rect 224861 470112 545179 470114
rect 224861 470056 224866 470112
rect 224922 470056 545118 470112
rect 545174 470056 545179 470112
rect 224861 470054 545179 470056
rect 224861 470051 224927 470054
rect 545113 470051 545179 470054
rect 225965 469978 226031 469981
rect 546493 469978 546559 469981
rect 225965 469976 546559 469978
rect 225965 469920 225970 469976
rect 226026 469920 546498 469976
rect 546554 469920 546559 469976
rect 225965 469918 546559 469920
rect 225965 469915 226031 469918
rect 546493 469915 546559 469918
rect 68686 469780 68692 469844
rect 68756 469842 68762 469844
rect 208894 469842 208900 469844
rect 68756 469782 208900 469842
rect 68756 469780 68762 469782
rect 208894 469780 208900 469782
rect 208964 469780 208970 469844
rect 222101 469842 222167 469845
rect 543733 469842 543799 469845
rect 222101 469840 543799 469842
rect 222101 469784 222106 469840
rect 222162 469784 543738 469840
rect 543794 469784 543799 469840
rect 222101 469782 543799 469784
rect 222101 469779 222167 469782
rect 543733 469779 543799 469782
rect 232957 469706 233023 469709
rect 543825 469706 543891 469709
rect 232957 469704 543891 469706
rect 232957 469648 232962 469704
rect 233018 469648 543830 469704
rect 543886 469648 543891 469704
rect 232957 469646 543891 469648
rect 232957 469643 233023 469646
rect 543825 469643 543891 469646
rect 275185 468754 275251 468757
rect 291326 468754 291332 468756
rect 275185 468752 291332 468754
rect 275185 468696 275190 468752
rect 275246 468696 291332 468752
rect 275185 468694 291332 468696
rect 275185 468691 275251 468694
rect 291326 468692 291332 468694
rect 291396 468692 291402 468756
rect 237189 468618 237255 468621
rect 496261 468618 496327 468621
rect 237189 468616 496327 468618
rect 237189 468560 237194 468616
rect 237250 468560 496266 468616
rect 496322 468560 496327 468616
rect 237189 468558 496327 468560
rect 237189 468555 237255 468558
rect 496261 468555 496327 468558
rect 68277 468482 68343 468485
rect 155217 468482 155283 468485
rect 68277 468480 155283 468482
rect 68277 468424 68282 468480
rect 68338 468424 155222 468480
rect 155278 468424 155283 468480
rect 68277 468422 155283 468424
rect 68277 468419 68343 468422
rect 155217 468419 155283 468422
rect 238518 468420 238524 468484
rect 238588 468482 238594 468484
rect 539358 468482 539364 468484
rect 238588 468422 539364 468482
rect 238588 468420 238594 468422
rect 539358 468420 539364 468422
rect 539428 468420 539434 468484
rect 256969 467530 257035 467533
rect 290181 467530 290247 467533
rect 256969 467528 290247 467530
rect 256969 467472 256974 467528
rect 257030 467472 290186 467528
rect 290242 467472 290247 467528
rect 256969 467470 290247 467472
rect 256969 467467 257035 467470
rect 290181 467467 290247 467470
rect 3550 467332 3556 467396
rect 3620 467394 3626 467396
rect 282862 467394 282868 467396
rect 3620 467334 282868 467394
rect 3620 467332 3626 467334
rect 282862 467332 282868 467334
rect 282932 467332 282938 467396
rect 235809 467258 235875 467261
rect 533521 467258 533587 467261
rect 235809 467256 533587 467258
rect 235809 467200 235814 467256
rect 235870 467200 533526 467256
rect 533582 467200 533587 467256
rect 235809 467198 533587 467200
rect 235809 467195 235875 467198
rect 533521 467195 533587 467198
rect 235717 467122 235783 467125
rect 534901 467122 534967 467125
rect 235717 467120 534967 467122
rect 235717 467064 235722 467120
rect 235778 467064 534906 467120
rect 534962 467064 534967 467120
rect 235717 467062 534967 467064
rect 235717 467059 235783 467062
rect 534901 467059 534967 467062
rect 246849 466034 246915 466037
rect 291193 466034 291259 466037
rect 246849 466032 291259 466034
rect 246849 465976 246854 466032
rect 246910 465976 291198 466032
rect 291254 465976 291259 466032
rect 246849 465974 291259 465976
rect 246849 465971 246915 465974
rect 291193 465971 291259 465974
rect 235901 465898 235967 465901
rect 493501 465898 493567 465901
rect 235901 465896 493567 465898
rect 235901 465840 235906 465896
rect 235962 465840 493506 465896
rect 493562 465840 493567 465896
rect 235901 465838 493567 465840
rect 235901 465835 235967 465838
rect 493501 465835 493567 465838
rect 233141 465762 233207 465765
rect 580257 465762 580323 465765
rect 233141 465760 580323 465762
rect 233141 465704 233146 465760
rect 233202 465704 580262 465760
rect 580318 465704 580323 465760
rect 233141 465702 580323 465704
rect 233141 465699 233207 465702
rect 580257 465699 580323 465702
rect 245837 464538 245903 464541
rect 289261 464538 289327 464541
rect 245837 464536 289327 464538
rect 245837 464480 245842 464536
rect 245898 464480 289266 464536
rect 289322 464480 289327 464536
rect 245837 464478 289327 464480
rect 245837 464475 245903 464478
rect 289261 464475 289327 464478
rect 164785 464402 164851 464405
rect 231117 464402 231183 464405
rect 164785 464400 231183 464402
rect 164785 464344 164790 464400
rect 164846 464344 231122 464400
rect 231178 464344 231183 464400
rect 164785 464342 231183 464344
rect 164785 464339 164851 464342
rect 231117 464339 231183 464342
rect 236913 464402 236979 464405
rect 511441 464402 511507 464405
rect 236913 464400 511507 464402
rect 236913 464344 236918 464400
rect 236974 464344 511446 464400
rect 511502 464344 511507 464400
rect 236913 464342 511507 464344
rect 236913 464339 236979 464342
rect 511441 464339 511507 464342
rect 252921 463042 252987 463045
rect 291837 463042 291903 463045
rect 252921 463040 291903 463042
rect 252921 462984 252926 463040
rect 252982 462984 291842 463040
rect 291898 462984 291903 463040
rect 252921 462982 291903 462984
rect 252921 462979 252987 462982
rect 291837 462979 291903 462982
rect 237005 462906 237071 462909
rect 492121 462906 492187 462909
rect 237005 462904 492187 462906
rect 237005 462848 237010 462904
rect 237066 462848 492126 462904
rect 492182 462848 492187 462904
rect 237005 462846 492187 462848
rect 237005 462843 237071 462846
rect 492121 462843 492187 462846
rect -960 462634 480 462724
rect 287094 462634 287100 462636
rect -960 462574 287100 462634
rect -960 462484 480 462574
rect 287094 462572 287100 462574
rect 287164 462572 287170 462636
rect 68134 461484 68140 461548
rect 68204 461546 68210 461548
rect 173014 461546 173020 461548
rect 68204 461486 173020 461546
rect 68204 461484 68210 461486
rect 173014 461484 173020 461486
rect 173084 461484 173090 461548
rect 248873 460322 248939 460325
rect 292021 460322 292087 460325
rect 248873 460320 292087 460322
rect 248873 460264 248878 460320
rect 248934 460264 292026 460320
rect 292082 460264 292087 460320
rect 248873 460262 292087 460264
rect 248873 460259 248939 460262
rect 292021 460259 292087 460262
rect 236821 460186 236887 460189
rect 514201 460186 514267 460189
rect 236821 460184 514267 460186
rect 236821 460128 236826 460184
rect 236882 460128 514206 460184
rect 514262 460128 514267 460184
rect 236821 460126 514267 460128
rect 236821 460123 236887 460126
rect 514201 460123 514267 460126
rect 261017 459098 261083 459101
rect 289813 459098 289879 459101
rect 261017 459096 289879 459098
rect 261017 459040 261022 459096
rect 261078 459040 289818 459096
rect 289874 459040 289879 459096
rect 261017 459038 289879 459040
rect 261017 459035 261083 459038
rect 289813 459035 289879 459038
rect 235441 458962 235507 458965
rect 528001 458962 528067 458965
rect 235441 458960 528067 458962
rect 235441 458904 235446 458960
rect 235502 458904 528006 458960
rect 528062 458904 528067 458960
rect 235441 458902 528067 458904
rect 235441 458899 235507 458902
rect 528001 458899 528067 458902
rect 235758 458764 235764 458828
rect 235828 458826 235834 458828
rect 542905 458826 542971 458829
rect 235828 458824 542971 458826
rect 235828 458768 542910 458824
rect 542966 458768 542971 458824
rect 235828 458766 542971 458768
rect 235828 458764 235834 458766
rect 542905 458763 542971 458766
rect 580349 458146 580415 458149
rect 583520 458146 584960 458236
rect 580349 458144 584960 458146
rect 580349 458088 580354 458144
rect 580410 458088 584960 458144
rect 580349 458086 584960 458088
rect 580349 458083 580415 458086
rect 583520 457996 584960 458086
rect 279233 456242 279299 456245
rect 291142 456242 291148 456244
rect 279233 456240 291148 456242
rect 279233 456184 279238 456240
rect 279294 456184 291148 456240
rect 279233 456182 291148 456184
rect 279233 456179 279299 456182
rect 291142 456180 291148 456182
rect 291212 456180 291218 456244
rect 3366 456044 3372 456108
rect 3436 456106 3442 456108
rect 210366 456106 210372 456108
rect 3436 456046 210372 456106
rect 3436 456044 3442 456046
rect 210366 456044 210372 456046
rect 210436 456044 210442 456108
rect 238150 456044 238156 456108
rect 238220 456106 238226 456108
rect 541014 456106 541020 456108
rect 238220 456046 541020 456106
rect 238220 456044 238226 456046
rect 541014 456044 541020 456046
rect 541084 456044 541090 456108
rect 110137 454746 110203 454749
rect 226977 454746 227043 454749
rect 110137 454744 227043 454746
rect 110137 454688 110142 454744
rect 110198 454688 226982 454744
rect 227038 454688 227043 454744
rect 110137 454686 227043 454688
rect 110137 454683 110203 454686
rect 226977 454683 227043 454686
rect 239489 454746 239555 454749
rect 286225 454746 286291 454749
rect 239489 454744 286291 454746
rect 239489 454688 239494 454744
rect 239550 454688 286230 454744
rect 286286 454688 286291 454744
rect 239489 454686 286291 454688
rect 239489 454683 239555 454686
rect 286225 454683 286291 454686
rect 4061 453386 4127 453389
rect 283005 453386 283071 453389
rect 4061 453384 283071 453386
rect 4061 453328 4066 453384
rect 4122 453328 283010 453384
rect 283066 453328 283071 453384
rect 4061 453326 283071 453328
rect 4061 453323 4127 453326
rect 283005 453323 283071 453326
rect 235073 453250 235139 453253
rect 536281 453250 536347 453253
rect 235073 453248 536347 453250
rect 235073 453192 235078 453248
rect 235134 453192 536286 453248
rect 536342 453192 536347 453248
rect 235073 453190 536347 453192
rect 235073 453187 235139 453190
rect 536281 453187 536347 453190
rect 234153 451890 234219 451893
rect 542813 451890 542879 451893
rect 234153 451888 542879 451890
rect 234153 451832 234158 451888
rect 234214 451832 542818 451888
rect 542874 451832 542879 451888
rect 234153 451830 542879 451832
rect 234153 451827 234219 451830
rect 542813 451827 542879 451830
rect 237281 450802 237347 450805
rect 332501 450802 332567 450805
rect 237281 450800 332567 450802
rect 237281 450744 237286 450800
rect 237342 450744 332506 450800
rect 332562 450744 332567 450800
rect 237281 450742 332567 450744
rect 237281 450739 237347 450742
rect 332501 450739 332567 450742
rect 235165 450666 235231 450669
rect 529381 450666 529447 450669
rect 235165 450664 529447 450666
rect 235165 450608 235170 450664
rect 235226 450608 529386 450664
rect 529442 450608 529447 450664
rect 235165 450606 529447 450608
rect 235165 450603 235231 450606
rect 529381 450603 529447 450606
rect 234102 450468 234108 450532
rect 234172 450530 234178 450532
rect 542854 450530 542860 450532
rect 234172 450470 542860 450530
rect 234172 450468 234178 450470
rect 542854 450468 542860 450470
rect 542924 450468 542930 450532
rect -960 449578 480 449668
rect 227662 449578 227668 449580
rect -960 449518 227668 449578
rect -960 449428 480 449518
rect 227662 449516 227668 449518
rect 227732 449516 227738 449580
rect 237230 449516 237236 449580
rect 237300 449578 237306 449580
rect 397453 449578 397519 449581
rect 237300 449576 397519 449578
rect 237300 449520 397458 449576
rect 397514 449520 397519 449576
rect 237300 449518 397519 449520
rect 237300 449516 237306 449518
rect 397453 449515 397519 449518
rect 239673 449442 239739 449445
rect 521101 449442 521167 449445
rect 239673 449440 521167 449442
rect 239673 449384 239678 449440
rect 239734 449384 521106 449440
rect 521162 449384 521167 449440
rect 239673 449382 521167 449384
rect 239673 449379 239739 449382
rect 521101 449379 521167 449382
rect 237966 449244 237972 449308
rect 238036 449306 238042 449308
rect 539777 449306 539843 449309
rect 238036 449304 539843 449306
rect 238036 449248 539782 449304
rect 539838 449248 539843 449304
rect 238036 449246 539843 449248
rect 238036 449244 238042 449246
rect 539777 449243 539843 449246
rect 233785 449170 233851 449173
rect 542445 449170 542511 449173
rect 233785 449168 542511 449170
rect 233785 449112 233790 449168
rect 233846 449112 542450 449168
rect 542506 449112 542511 449168
rect 233785 449110 542511 449112
rect 233785 449107 233851 449110
rect 542445 449107 542511 449110
rect 234981 448218 235047 448221
rect 494881 448218 494947 448221
rect 234981 448216 494947 448218
rect 234981 448160 234986 448216
rect 235042 448160 494886 448216
rect 494942 448160 494947 448216
rect 234981 448158 494947 448160
rect 234981 448155 235047 448158
rect 494881 448155 494947 448158
rect 236729 448082 236795 448085
rect 500401 448082 500467 448085
rect 236729 448080 500467 448082
rect 236729 448024 236734 448080
rect 236790 448024 500406 448080
rect 500462 448024 500467 448080
rect 236729 448022 500467 448024
rect 236729 448019 236795 448022
rect 500401 448019 500467 448022
rect 239581 447946 239647 447949
rect 518341 447946 518407 447949
rect 239581 447944 518407 447946
rect 239581 447888 239586 447944
rect 239642 447888 518346 447944
rect 518402 447888 518407 447944
rect 239581 447886 518407 447888
rect 239581 447883 239647 447886
rect 518341 447883 518407 447886
rect 236637 447810 236703 447813
rect 515581 447810 515647 447813
rect 236637 447808 515647 447810
rect 236637 447752 236642 447808
rect 236698 447752 515586 447808
rect 515642 447752 515647 447808
rect 236637 447750 515647 447752
rect 236637 447747 236703 447750
rect 515581 447747 515647 447750
rect 239397 446994 239463 446997
rect 280153 446994 280219 446997
rect 239397 446992 280219 446994
rect 239397 446936 239402 446992
rect 239458 446936 280158 446992
rect 280214 446936 280219 446992
rect 239397 446934 280219 446936
rect 239397 446931 239463 446934
rect 280153 446931 280219 446934
rect 235533 446858 235599 446861
rect 497641 446858 497707 446861
rect 235533 446856 497707 446858
rect 235533 446800 235538 446856
rect 235594 446800 497646 446856
rect 497702 446800 497707 446856
rect 235533 446798 497707 446800
rect 235533 446795 235599 446798
rect 497641 446795 497707 446798
rect 238569 446722 238635 446725
rect 539961 446722 540027 446725
rect 238569 446720 540027 446722
rect 238569 446664 238574 446720
rect 238630 446664 539966 446720
rect 540022 446664 540027 446720
rect 238569 446662 540027 446664
rect 238569 446659 238635 446662
rect 539961 446659 540027 446662
rect 235574 446524 235580 446588
rect 235644 446586 235650 446588
rect 537661 446586 537727 446589
rect 235644 446584 537727 446586
rect 235644 446528 537666 446584
rect 537722 446528 537727 446584
rect 235644 446526 537727 446528
rect 235644 446524 235650 446526
rect 537661 446523 537727 446526
rect 68553 446450 68619 446453
rect 199469 446450 199535 446453
rect 68553 446448 199535 446450
rect 68553 446392 68558 446448
rect 68614 446392 199474 446448
rect 199530 446392 199535 446448
rect 68553 446390 199535 446392
rect 68553 446387 68619 446390
rect 199469 446387 199535 446390
rect 233877 446450 233943 446453
rect 542353 446450 542419 446453
rect 233877 446448 542419 446450
rect 233877 446392 233882 446448
rect 233938 446392 542358 446448
rect 542414 446392 542419 446448
rect 233877 446390 542419 446392
rect 233877 446387 233943 446390
rect 542353 446387 542419 446390
rect 239305 445498 239371 445501
rect 274081 445498 274147 445501
rect 239305 445496 274147 445498
rect 239305 445440 239310 445496
rect 239366 445440 274086 445496
rect 274142 445440 274147 445496
rect 239305 445438 274147 445440
rect 239305 445435 239371 445438
rect 274081 445435 274147 445438
rect 235349 445362 235415 445365
rect 501781 445362 501847 445365
rect 235349 445360 501847 445362
rect 235349 445304 235354 445360
rect 235410 445304 501786 445360
rect 501842 445304 501847 445360
rect 235349 445302 501847 445304
rect 235349 445299 235415 445302
rect 501781 445299 501847 445302
rect 236453 445226 236519 445229
rect 522481 445226 522547 445229
rect 236453 445224 522547 445226
rect 236453 445168 236458 445224
rect 236514 445168 522486 445224
rect 522542 445168 522547 445224
rect 236453 445166 522547 445168
rect 236453 445163 236519 445166
rect 522481 445163 522547 445166
rect 238661 445090 238727 445093
rect 540053 445090 540119 445093
rect 238661 445088 540119 445090
rect 238661 445032 238666 445088
rect 238722 445032 540058 445088
rect 540114 445032 540119 445088
rect 238661 445030 540119 445032
rect 238661 445027 238727 445030
rect 540053 445027 540119 445030
rect 233969 444954 234035 444957
rect 542537 444954 542603 444957
rect 233969 444952 542603 444954
rect 233969 444896 233974 444952
rect 234030 444896 542542 444952
rect 542598 444896 542603 444952
rect 233969 444894 542603 444896
rect 233969 444891 234035 444894
rect 542537 444891 542603 444894
rect 583520 444668 584960 444908
rect 57278 444212 57284 444276
rect 57348 444274 57354 444276
rect 240041 444274 240107 444277
rect 57348 444272 240107 444274
rect 57348 444216 240046 444272
rect 240102 444216 240107 444272
rect 57348 444214 240107 444216
rect 57348 444212 57354 444214
rect 240041 444211 240107 444214
rect 59997 444138 60063 444141
rect 226885 444138 226951 444141
rect 59997 444136 226951 444138
rect 59997 444080 60002 444136
rect 60058 444080 226890 444136
rect 226946 444080 226951 444136
rect 59997 444078 226951 444080
rect 59997 444075 60063 444078
rect 226885 444075 226951 444078
rect 227118 444078 231870 444138
rect 59854 443940 59860 444004
rect 59924 444002 59930 444004
rect 227118 444002 227178 444078
rect 59924 443942 227178 444002
rect 231810 444002 231870 444078
rect 235206 444076 235212 444140
rect 235276 444138 235282 444140
rect 235625 444138 235691 444141
rect 235276 444136 235691 444138
rect 235276 444080 235630 444136
rect 235686 444080 235691 444136
rect 235276 444078 235691 444080
rect 235276 444076 235282 444078
rect 235625 444075 235691 444078
rect 239121 444138 239187 444141
rect 268009 444138 268075 444141
rect 239121 444136 268075 444138
rect 239121 444080 239126 444136
rect 239182 444080 268014 444136
rect 268070 444080 268075 444136
rect 239121 444078 268075 444080
rect 239121 444075 239187 444078
rect 268009 444075 268075 444078
rect 287278 444002 287284 444004
rect 231810 443942 287284 444002
rect 59924 443940 59930 443942
rect 287278 443940 287284 443942
rect 287348 443940 287354 444004
rect 226885 443866 226951 443869
rect 237373 443866 237439 443869
rect 226885 443864 237439 443866
rect 226885 443808 226890 443864
rect 226946 443808 237378 443864
rect 237434 443808 237439 443864
rect 226885 443806 237439 443808
rect 226885 443803 226951 443806
rect 237373 443803 237439 443806
rect 237557 443866 237623 443869
rect 499021 443866 499087 443869
rect 237557 443864 499087 443866
rect 237557 443808 237562 443864
rect 237618 443808 499026 443864
rect 499082 443808 499087 443864
rect 237557 443806 499087 443808
rect 237557 443803 237623 443806
rect 499021 443803 499087 443806
rect 236545 443730 236611 443733
rect 516961 443730 517027 443733
rect 236545 443728 517027 443730
rect 236545 443672 236550 443728
rect 236606 443672 516966 443728
rect 517022 443672 517027 443728
rect 236545 443670 517027 443672
rect 236545 443667 236611 443670
rect 516961 443667 517027 443670
rect 235257 443594 235323 443597
rect 237557 443594 237623 443597
rect 235257 443592 237623 443594
rect 235257 443536 235262 443592
rect 235318 443536 237562 443592
rect 237618 443536 237623 443592
rect 235257 443534 237623 443536
rect 235257 443531 235323 443534
rect 237557 443531 237623 443534
rect 238293 443594 238359 443597
rect 539593 443594 539659 443597
rect 238293 443592 539659 443594
rect 238293 443536 238298 443592
rect 238354 443536 539598 443592
rect 539654 443536 539659 443592
rect 238293 443534 539659 443536
rect 238293 443531 238359 443534
rect 539593 443531 539659 443534
rect 238017 443458 238083 443461
rect 300117 443458 300183 443461
rect 238017 443456 300183 443458
rect 238017 443400 238022 443456
rect 238078 443400 300122 443456
rect 300178 443400 300183 443456
rect 238017 443398 300183 443400
rect 238017 443395 238083 443398
rect 300117 443395 300183 443398
rect 218697 443050 218763 443053
rect 283097 443050 283163 443053
rect 218697 443048 283163 443050
rect 218697 442992 218702 443048
rect 218758 442992 283102 443048
rect 283158 442992 283163 443048
rect 218697 442990 283163 442992
rect 218697 442987 218763 442990
rect 283097 442987 283163 442990
rect 270125 442914 270191 442917
rect 271229 442914 271295 442917
rect 270125 442912 271295 442914
rect 270125 442856 270130 442912
rect 270186 442856 271234 442912
rect 271290 442856 271295 442912
rect 270125 442854 271295 442856
rect 270125 442851 270191 442854
rect 271229 442851 271295 442854
rect 272149 442914 272215 442917
rect 288985 442914 289051 442917
rect 272149 442912 289051 442914
rect 272149 442856 272154 442912
rect 272210 442856 288990 442912
rect 289046 442856 289051 442912
rect 272149 442854 289051 442856
rect 272149 442851 272215 442854
rect 288985 442851 289051 442854
rect 289721 442914 289787 442917
rect 292757 442914 292823 442917
rect 289721 442912 292823 442914
rect 289721 442856 289726 442912
rect 289782 442856 292762 442912
rect 292818 442856 292823 442912
rect 289721 442854 292823 442856
rect 289721 442851 289787 442854
rect 292757 442851 292823 442854
rect 228265 442778 228331 442781
rect 254025 442778 254091 442781
rect 228265 442776 254091 442778
rect 228265 442720 228270 442776
rect 228326 442720 254030 442776
rect 254086 442720 254091 442776
rect 228265 442718 254091 442720
rect 228265 442715 228331 442718
rect 254025 442715 254091 442718
rect 265065 442778 265131 442781
rect 295425 442778 295491 442781
rect 265065 442776 295491 442778
rect 265065 442720 265070 442776
rect 265126 442720 295430 442776
rect 295486 442720 295491 442776
rect 265065 442718 295491 442720
rect 265065 442715 265131 442718
rect 295425 442715 295491 442718
rect 239029 442642 239095 442645
rect 261937 442642 262003 442645
rect 239029 442640 262003 442642
rect 239029 442584 239034 442640
rect 239090 442584 261942 442640
rect 261998 442584 262003 442640
rect 239029 442582 262003 442584
rect 239029 442579 239095 442582
rect 261937 442579 262003 442582
rect 266077 442642 266143 442645
rect 296713 442642 296779 442645
rect 266077 442640 296779 442642
rect 266077 442584 266082 442640
rect 266138 442584 296718 442640
rect 296774 442584 296779 442640
rect 266077 442582 296779 442584
rect 266077 442579 266143 442582
rect 296713 442579 296779 442582
rect 48129 442506 48195 442509
rect 240041 442506 240107 442509
rect 48129 442504 240107 442506
rect 48129 442448 48134 442504
rect 48190 442448 240046 442504
rect 240102 442448 240107 442504
rect 48129 442446 240107 442448
rect 48129 442443 48195 442446
rect 240041 442443 240107 442446
rect 250897 442506 250963 442509
rect 254393 442506 254459 442509
rect 293125 442506 293191 442509
rect 250897 442504 254226 442506
rect 250897 442448 250902 442504
rect 250958 442448 254226 442504
rect 250897 442446 254226 442448
rect 250897 442443 250963 442446
rect 224902 442308 224908 442372
rect 224972 442370 224978 442372
rect 253933 442370 253999 442373
rect 224972 442368 253999 442370
rect 224972 442312 253938 442368
rect 253994 442312 253999 442368
rect 224972 442310 253999 442312
rect 224972 442308 224978 442310
rect 253933 442307 253999 442310
rect 226149 442234 226215 442237
rect 251081 442234 251147 442237
rect 226149 442232 251147 442234
rect 226149 442176 226154 442232
rect 226210 442176 251086 442232
rect 251142 442176 251147 442232
rect 226149 442174 251147 442176
rect 254166 442234 254226 442446
rect 254393 442504 293191 442506
rect 254393 442448 254398 442504
rect 254454 442448 293130 442504
rect 293186 442448 293191 442504
rect 254393 442446 293191 442448
rect 254393 442443 254459 442446
rect 293125 442443 293191 442446
rect 254945 442370 255011 442373
rect 294413 442370 294479 442373
rect 254945 442368 294479 442370
rect 254945 442312 254950 442368
rect 255006 442312 294418 442368
rect 294474 442312 294479 442368
rect 254945 442310 294479 442312
rect 254945 442307 255011 442310
rect 294413 442307 294479 442310
rect 290549 442234 290615 442237
rect 254166 442232 290615 442234
rect 254166 442176 290554 442232
rect 290610 442176 290615 442232
rect 254166 442174 290615 442176
rect 226149 442171 226215 442174
rect 251081 442171 251147 442174
rect 290549 442171 290615 442174
rect 223982 442036 223988 442100
rect 224052 442098 224058 442100
rect 229001 442098 229067 442101
rect 224052 442096 229067 442098
rect 224052 442040 229006 442096
rect 229062 442040 229067 442096
rect 224052 442038 229067 442040
rect 224052 442036 224058 442038
rect 229001 442035 229067 442038
rect 229645 442098 229711 442101
rect 264973 442098 265039 442101
rect 229645 442096 265039 442098
rect 229645 442040 229650 442096
rect 229706 442040 264978 442096
rect 265034 442040 265039 442096
rect 229645 442038 265039 442040
rect 229645 442035 229711 442038
rect 264973 442035 265039 442038
rect 274173 442098 274239 442101
rect 289629 442098 289695 442101
rect 274173 442096 289695 442098
rect 274173 442040 274178 442096
rect 274234 442040 289634 442096
rect 289690 442040 289695 442096
rect 274173 442038 289695 442040
rect 274173 442035 274239 442038
rect 289629 442035 289695 442038
rect 218830 441900 218836 441964
rect 218900 441962 218906 441964
rect 270401 441962 270467 441965
rect 218900 441960 270467 441962
rect 218900 441904 270406 441960
rect 270462 441904 270467 441960
rect 218900 441902 270467 441904
rect 218900 441900 218906 441902
rect 270401 441899 270467 441902
rect 289629 441962 289695 441965
rect 293217 441962 293283 441965
rect 289629 441960 293283 441962
rect 289629 441904 289634 441960
rect 289690 441904 293222 441960
rect 293278 441904 293283 441960
rect 289629 441902 293283 441904
rect 289629 441899 289695 441902
rect 293217 441899 293283 441902
rect 218646 441764 218652 441828
rect 218716 441826 218722 441828
rect 273253 441826 273319 441829
rect 218716 441824 273319 441826
rect 218716 441768 273258 441824
rect 273314 441768 273319 441824
rect 218716 441766 273319 441768
rect 218716 441764 218722 441766
rect 273253 441763 273319 441766
rect 221038 441628 221044 441692
rect 221108 441690 221114 441692
rect 229645 441690 229711 441693
rect 233969 441692 234035 441693
rect 233918 441690 233924 441692
rect 221108 441688 229711 441690
rect 221108 441632 229650 441688
rect 229706 441632 229711 441688
rect 221108 441630 229711 441632
rect 233878 441630 233924 441690
rect 233988 441688 234035 441692
rect 234030 441632 234035 441688
rect 221108 441628 221114 441630
rect 229645 441627 229711 441630
rect 233918 441628 233924 441630
rect 233988 441628 234035 441632
rect 233969 441627 234035 441628
rect 228398 441492 228404 441556
rect 228468 441554 228474 441556
rect 281901 441554 281967 441557
rect 228468 441552 281967 441554
rect 228468 441496 281906 441552
rect 281962 441496 281967 441552
rect 228468 441494 281967 441496
rect 228468 441492 228474 441494
rect 281901 441491 281967 441494
rect 226926 441356 226932 441420
rect 226996 441418 227002 441420
rect 282361 441418 282427 441421
rect 226996 441416 282427 441418
rect 226996 441360 282366 441416
rect 282422 441360 282427 441416
rect 226996 441358 282427 441360
rect 226996 441356 227002 441358
rect 282361 441355 282427 441358
rect 112478 441220 112484 441284
rect 112548 441282 112554 441284
rect 280654 441282 280660 441284
rect 112548 441222 280660 441282
rect 112548 441220 112554 441222
rect 280654 441220 280660 441222
rect 280724 441220 280730 441284
rect 230974 441084 230980 441148
rect 231044 441146 231050 441148
rect 231044 441086 279618 441146
rect 231044 441084 231050 441086
rect 219934 440948 219940 441012
rect 220004 441010 220010 441012
rect 220004 440950 229754 441010
rect 220004 440948 220010 440950
rect 222009 440874 222075 440877
rect 229001 440874 229067 440877
rect 222009 440872 229067 440874
rect 222009 440816 222014 440872
rect 222070 440816 229006 440872
rect 229062 440816 229067 440872
rect 222009 440814 229067 440816
rect 229694 440874 229754 440950
rect 230054 440948 230060 441012
rect 230124 441010 230130 441012
rect 230124 440950 279250 441010
rect 230124 440948 230130 440950
rect 229694 440814 279066 440874
rect 222009 440811 222075 440814
rect 229001 440811 229067 440814
rect 112989 440738 113055 440741
rect 229645 440738 229711 440741
rect 112989 440736 229711 440738
rect 112989 440680 112994 440736
rect 113050 440680 229650 440736
rect 229706 440680 229711 440736
rect 112989 440678 229711 440680
rect 112989 440675 113055 440678
rect 229645 440675 229711 440678
rect 112294 440540 112300 440604
rect 112364 440602 112370 440604
rect 230473 440602 230539 440605
rect 112364 440600 230539 440602
rect 112364 440544 230478 440600
rect 230534 440544 230539 440600
rect 112364 440542 230539 440544
rect 112364 440540 112370 440542
rect 230473 440539 230539 440542
rect 112846 440404 112852 440468
rect 112916 440466 112922 440468
rect 278814 440466 278820 440468
rect 112916 440406 278820 440466
rect 112916 440404 112922 440406
rect 278814 440404 278820 440406
rect 278884 440404 278890 440468
rect 279006 440466 279066 440814
rect 279190 440602 279250 440950
rect 279558 440874 279618 441086
rect 282269 440874 282335 440877
rect 279558 440872 282335 440874
rect 279558 440816 282274 440872
rect 282330 440816 282335 440872
rect 279558 440814 282335 440816
rect 282269 440811 282335 440814
rect 281625 440602 281691 440605
rect 279190 440600 281691 440602
rect 279190 440544 281630 440600
rect 281686 440544 281691 440600
rect 279190 440542 281691 440544
rect 281625 440539 281691 440542
rect 281533 440466 281599 440469
rect 279006 440464 281599 440466
rect 279006 440408 281538 440464
rect 281594 440408 281599 440464
rect 279006 440406 281599 440408
rect 281533 440403 281599 440406
rect 226190 440268 226196 440332
rect 226260 440330 226266 440332
rect 227161 440330 227227 440333
rect 226260 440328 227227 440330
rect 226260 440272 227166 440328
rect 227222 440272 227227 440328
rect 226260 440270 227227 440272
rect 226260 440268 226266 440270
rect 227161 440267 227227 440270
rect 227846 440268 227852 440332
rect 227916 440330 227922 440332
rect 228909 440330 228975 440333
rect 227916 440328 228975 440330
rect 227916 440272 228914 440328
rect 228970 440272 228975 440328
rect 227916 440270 228975 440272
rect 227916 440268 227922 440270
rect 228909 440267 228975 440270
rect 230422 440268 230428 440332
rect 230492 440330 230498 440332
rect 231393 440330 231459 440333
rect 230492 440328 231459 440330
rect 230492 440272 231398 440328
rect 231454 440272 231459 440328
rect 230492 440270 231459 440272
rect 230492 440268 230498 440270
rect 231393 440267 231459 440270
rect 231894 440268 231900 440332
rect 231964 440330 231970 440332
rect 232681 440330 232747 440333
rect 231964 440328 232747 440330
rect 231964 440272 232686 440328
rect 232742 440272 232747 440328
rect 231964 440270 232747 440272
rect 231964 440268 231970 440270
rect 232681 440267 232747 440270
rect 222694 440132 222700 440196
rect 222764 440194 222770 440196
rect 222764 440134 224970 440194
rect 222764 440132 222770 440134
rect 224910 440058 224970 440134
rect 227662 440132 227668 440196
rect 227732 440194 227738 440196
rect 228909 440194 228975 440197
rect 227732 440192 228975 440194
rect 227732 440136 228914 440192
rect 228970 440136 228975 440192
rect 227732 440134 228975 440136
rect 227732 440132 227738 440134
rect 228909 440131 228975 440134
rect 234889 440194 234955 440197
rect 282453 440194 282519 440197
rect 234889 440192 282519 440194
rect 234889 440136 234894 440192
rect 234950 440136 282458 440192
rect 282514 440136 282519 440192
rect 234889 440134 282519 440136
rect 234889 440131 234955 440134
rect 282453 440131 282519 440134
rect 229645 440058 229711 440061
rect 281717 440058 281783 440061
rect 224910 440056 229711 440058
rect 224910 440000 229650 440056
rect 229706 440000 229711 440056
rect 224910 439998 229711 440000
rect 229645 439995 229711 439998
rect 229878 440056 281783 440058
rect 229878 440000 281722 440056
rect 281778 440000 281783 440056
rect 229878 439998 281783 440000
rect 228214 439860 228220 439924
rect 228284 439922 228290 439924
rect 229878 439922 229938 439998
rect 281717 439995 281783 439998
rect 228284 439862 229938 439922
rect 230013 439922 230079 439925
rect 281942 439922 281948 439924
rect 230013 439920 281948 439922
rect 230013 439864 230018 439920
rect 230074 439864 281948 439920
rect 230013 439862 281948 439864
rect 228284 439860 228290 439862
rect 230013 439859 230079 439862
rect 281942 439860 281948 439862
rect 282012 439860 282018 439924
rect 224166 439724 224172 439788
rect 224236 439786 224242 439788
rect 281758 439786 281764 439788
rect 224236 439726 281764 439786
rect 224236 439724 224242 439726
rect 281758 439724 281764 439726
rect 281828 439724 281834 439788
rect 227110 439588 227116 439652
rect 227180 439650 227186 439652
rect 229369 439650 229435 439653
rect 227180 439648 229435 439650
rect 227180 439592 229374 439648
rect 229430 439592 229435 439648
rect 227180 439590 229435 439592
rect 227180 439588 227186 439590
rect 229369 439587 229435 439590
rect 229645 439650 229711 439653
rect 282310 439650 282316 439652
rect 229645 439648 282316 439650
rect 229645 439592 229650 439648
rect 229706 439592 282316 439648
rect 229645 439590 282316 439592
rect 229645 439587 229711 439590
rect 282310 439588 282316 439590
rect 282380 439588 282386 439652
rect 178534 439452 178540 439516
rect 178604 439514 178610 439516
rect 178604 439454 279434 439514
rect 178604 439452 178610 439454
rect 221222 439316 221228 439380
rect 221292 439378 221298 439380
rect 229001 439378 229067 439381
rect 221292 439376 229067 439378
rect 221292 439320 229006 439376
rect 229062 439320 229067 439376
rect 221292 439318 229067 439320
rect 221292 439316 221298 439318
rect 229001 439315 229067 439318
rect 231526 439316 231532 439380
rect 231596 439378 231602 439380
rect 234889 439378 234955 439381
rect 231596 439376 234955 439378
rect 231596 439320 234894 439376
rect 234950 439320 234955 439376
rect 231596 439318 234955 439320
rect 231596 439316 231602 439318
rect 234889 439315 234955 439318
rect 227662 439180 227668 439244
rect 227732 439242 227738 439244
rect 228725 439242 228791 439245
rect 227732 439240 228791 439242
rect 227732 439184 228730 439240
rect 228786 439184 228791 439240
rect 227732 439182 228791 439184
rect 227732 439180 227738 439182
rect 228725 439179 228791 439182
rect 113081 439106 113147 439109
rect 229645 439106 229711 439109
rect 113081 439104 229711 439106
rect 113081 439048 113086 439104
rect 113142 439048 229650 439104
rect 229706 439048 229711 439104
rect 113081 439046 229711 439048
rect 113081 439043 113147 439046
rect 229645 439043 229711 439046
rect 229870 439044 229876 439108
rect 229940 439106 229946 439108
rect 231025 439106 231091 439109
rect 229940 439104 231091 439106
rect 229940 439048 231030 439104
rect 231086 439048 231091 439104
rect 229940 439046 231091 439048
rect 229940 439044 229946 439046
rect 231025 439043 231091 439046
rect 239622 439044 239628 439108
rect 239692 439106 239698 439108
rect 239765 439106 239831 439109
rect 239692 439104 239831 439106
rect 239692 439048 239770 439104
rect 239826 439048 239831 439104
rect 239692 439046 239831 439048
rect 239692 439044 239698 439046
rect 239765 439043 239831 439046
rect 279374 438972 279434 439454
rect 112662 438908 112668 438972
rect 112732 438970 112738 438972
rect 112732 438910 279250 438970
rect 112732 438908 112738 438910
rect 279190 438834 279250 438910
rect 279366 438908 279372 438972
rect 279436 438908 279442 438972
rect 280838 438970 280844 438972
rect 279558 438910 280844 438970
rect 279558 438834 279618 438910
rect 280838 438908 280844 438910
rect 280908 438908 280914 438972
rect 279190 438774 279618 438834
rect 278814 438636 278820 438700
rect 278884 438698 278890 438700
rect 278884 438638 279802 438698
rect 278884 438636 278890 438638
rect 231158 438500 231164 438564
rect 231228 438562 231234 438564
rect 279550 438562 279556 438564
rect 231228 438502 279556 438562
rect 231228 438500 231234 438502
rect 279550 438500 279556 438502
rect 279620 438500 279626 438564
rect 279742 438396 279802 438638
rect 279366 437412 279372 437476
rect 279436 437412 279442 437476
rect 279374 437036 279434 437412
rect -960 436508 480 436748
rect 281625 435706 281691 435709
rect 279956 435704 281691 435706
rect 279956 435648 281630 435704
rect 281686 435648 281691 435704
rect 279956 435646 281691 435648
rect 281625 435643 281691 435646
rect 281533 434346 281599 434349
rect 279956 434344 281599 434346
rect 279956 434288 281538 434344
rect 281594 434288 281599 434344
rect 279956 434286 281599 434288
rect 281533 434283 281599 434286
rect 281901 432986 281967 432989
rect 279956 432984 281967 432986
rect 279956 432928 281906 432984
rect 281962 432928 281967 432984
rect 279956 432926 281967 432928
rect 281901 432923 281967 432926
rect 281942 431626 281948 431628
rect 279956 431566 281948 431626
rect 281942 431564 281948 431566
rect 282012 431564 282018 431628
rect 580257 431626 580323 431629
rect 583520 431626 584960 431716
rect 580257 431624 584960 431626
rect 580257 431568 580262 431624
rect 580318 431568 584960 431624
rect 580257 431566 584960 431568
rect 580257 431563 580323 431566
rect 583520 431476 584960 431566
rect 116209 431218 116275 431221
rect 211797 431218 211863 431221
rect 116209 431216 211863 431218
rect 116209 431160 116214 431216
rect 116270 431160 211802 431216
rect 211858 431160 211863 431216
rect 116209 431158 211863 431160
rect 116209 431155 116275 431158
rect 211797 431155 211863 431158
rect 281758 430266 281764 430268
rect 279956 430206 281764 430266
rect 281758 430204 281764 430206
rect 281828 430204 281834 430268
rect 282310 428906 282316 428908
rect 279956 428846 282316 428906
rect 282310 428844 282316 428846
rect 282380 428844 282386 428908
rect 282177 427546 282243 427549
rect 279956 427544 282243 427546
rect 279956 427488 282182 427544
rect 282238 427488 282243 427544
rect 279956 427486 282243 427488
rect 282177 427483 282243 427486
rect 280838 426186 280844 426188
rect 279956 426126 280844 426186
rect 280838 426124 280844 426126
rect 280908 426124 280914 426188
rect 282085 424826 282151 424829
rect 279956 424824 282151 424826
rect 279956 424768 282090 424824
rect 282146 424768 282151 424824
rect 279956 424766 282151 424768
rect 282085 424763 282151 424766
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 280654 423466 280660 423468
rect 279956 423406 280660 423466
rect 280654 423404 280660 423406
rect 280724 423404 280730 423468
rect 281901 422106 281967 422109
rect 279956 422104 281967 422106
rect 279956 422048 281906 422104
rect 281962 422048 281967 422104
rect 279956 422046 281967 422048
rect 281901 422043 281967 422046
rect 281809 420746 281875 420749
rect 279956 420744 281875 420746
rect 279956 420688 281814 420744
rect 281870 420688 281875 420744
rect 279956 420686 281875 420688
rect 281809 420683 281875 420686
rect 281717 419386 281783 419389
rect 279956 419384 281783 419386
rect 279956 419328 281722 419384
rect 281778 419328 281783 419384
rect 279956 419326 281783 419328
rect 281717 419323 281783 419326
rect 500166 418236 500172 418300
rect 500236 418298 500242 418300
rect 583520 418298 584960 418388
rect 500236 418238 584960 418298
rect 500236 418236 500242 418238
rect 583520 418148 584960 418238
rect 281625 418026 281691 418029
rect 279956 418024 281691 418026
rect 279956 417968 281630 418024
rect 281686 417968 281691 418024
rect 279956 417966 281691 417968
rect 281625 417963 281691 417966
rect 280981 416666 281047 416669
rect 279956 416664 281047 416666
rect 279956 416608 280986 416664
rect 281042 416608 281047 416664
rect 279956 416606 281047 416608
rect 280981 416603 281047 416606
rect 281533 415306 281599 415309
rect 279956 415304 281599 415306
rect 279956 415248 281538 415304
rect 281594 415248 281599 415304
rect 279956 415246 281599 415248
rect 281533 415243 281599 415246
rect 280889 413946 280955 413949
rect 279956 413944 280955 413946
rect 279956 413888 280894 413944
rect 280950 413888 280955 413944
rect 279956 413886 280955 413888
rect 280889 413883 280955 413886
rect 280797 412586 280863 412589
rect 279956 412584 280863 412586
rect 279956 412528 280802 412584
rect 280858 412528 280863 412584
rect 279956 412526 280863 412528
rect 280797 412523 280863 412526
rect 283097 411226 283163 411229
rect 279956 411224 283163 411226
rect 279956 411168 283102 411224
rect 283158 411168 283163 411224
rect 279956 411166 283163 411168
rect 283097 411163 283163 411166
rect -960 410546 480 410636
rect 223982 410546 223988 410548
rect -960 410486 223988 410546
rect -960 410396 480 410486
rect 223982 410484 223988 410486
rect 224052 410484 224058 410548
rect 224350 409940 224356 410004
rect 224420 410002 224426 410004
rect 224769 410002 224835 410005
rect 224420 410000 224835 410002
rect 224420 409944 224774 410000
rect 224830 409944 224835 410000
rect 224420 409942 224835 409944
rect 224420 409940 224426 409942
rect 224769 409939 224835 409942
rect 281901 409866 281967 409869
rect 279956 409864 281967 409866
rect 279956 409808 281906 409864
rect 281962 409808 281967 409864
rect 279956 409806 281967 409808
rect 281901 409803 281967 409806
rect 239489 408506 239555 408509
rect 281901 408506 281967 408509
rect 239489 408504 240212 408506
rect 239489 408448 239494 408504
rect 239550 408448 240212 408504
rect 239489 408446 240212 408448
rect 279956 408504 281967 408506
rect 279956 408448 281906 408504
rect 281962 408448 281967 408504
rect 279956 408446 281967 408448
rect 239489 408443 239555 408446
rect 281901 408443 281967 408446
rect 239397 407962 239463 407965
rect 239397 407960 240212 407962
rect 239397 407904 239402 407960
rect 239458 407904 240212 407960
rect 239397 407902 240212 407904
rect 239397 407899 239463 407902
rect 239305 407418 239371 407421
rect 239305 407416 240212 407418
rect 239305 407360 239310 407416
rect 239366 407360 240212 407416
rect 239305 407358 240212 407360
rect 239305 407355 239371 407358
rect 280705 407146 280771 407149
rect 279956 407144 280771 407146
rect 279956 407088 280710 407144
rect 280766 407088 280771 407144
rect 279956 407086 280771 407088
rect 280705 407083 280771 407086
rect 239213 406874 239279 406877
rect 239213 406872 240212 406874
rect 239213 406816 239218 406872
rect 239274 406816 240212 406872
rect 239213 406814 240212 406816
rect 239213 406811 239279 406814
rect 239029 406330 239095 406333
rect 239029 406328 240212 406330
rect 239029 406272 239034 406328
rect 239090 406272 240212 406328
rect 239029 406270 240212 406272
rect 239029 406267 239095 406270
rect 228357 406058 228423 406061
rect 239438 406058 239444 406060
rect 228357 406056 239444 406058
rect 228357 406000 228362 406056
rect 228418 406000 239444 406056
rect 228357 405998 239444 406000
rect 228357 405995 228423 405998
rect 239438 405996 239444 405998
rect 239508 405996 239514 406060
rect 228449 405786 228515 405789
rect 280521 405786 280587 405789
rect 228449 405784 240212 405786
rect 228449 405728 228454 405784
rect 228510 405728 240212 405784
rect 228449 405726 240212 405728
rect 279956 405784 280587 405786
rect 279956 405728 280526 405784
rect 280582 405728 280587 405784
rect 279956 405726 280587 405728
rect 228449 405723 228515 405726
rect 280521 405723 280587 405726
rect 239489 405242 239555 405245
rect 239489 405240 240212 405242
rect 239489 405184 239494 405240
rect 239550 405184 240212 405240
rect 239489 405182 240212 405184
rect 239489 405179 239555 405182
rect 579705 404970 579771 404973
rect 583520 404970 584960 405060
rect 579705 404968 584960 404970
rect 579705 404912 579710 404968
rect 579766 404912 584960 404968
rect 579705 404910 584960 404912
rect 579705 404907 579771 404910
rect 583520 404820 584960 404910
rect 231209 404698 231275 404701
rect 231209 404696 240212 404698
rect 231209 404640 231214 404696
rect 231270 404640 240212 404696
rect 231209 404638 240212 404640
rect 231209 404635 231275 404638
rect 280613 404426 280679 404429
rect 279956 404424 280679 404426
rect 279956 404368 280618 404424
rect 280674 404368 280679 404424
rect 279956 404366 280679 404368
rect 280613 404363 280679 404366
rect 237649 404154 237715 404157
rect 237649 404152 240212 404154
rect 237649 404096 237654 404152
rect 237710 404096 240212 404152
rect 237649 404094 240212 404096
rect 237649 404091 237715 404094
rect 231577 403610 231643 403613
rect 231577 403608 240212 403610
rect 231577 403552 231582 403608
rect 231638 403552 240212 403608
rect 231577 403550 240212 403552
rect 231577 403547 231643 403550
rect 225505 403066 225571 403069
rect 280429 403066 280495 403069
rect 225505 403064 240212 403066
rect 225505 403008 225510 403064
rect 225566 403008 240212 403064
rect 225505 403006 240212 403008
rect 279956 403064 280495 403066
rect 279956 403008 280434 403064
rect 280490 403008 280495 403064
rect 279956 403006 280495 403008
rect 225505 403003 225571 403006
rect 280429 403003 280495 403006
rect 219433 402522 219499 402525
rect 219433 402520 240212 402522
rect 219433 402464 219438 402520
rect 219494 402464 240212 402520
rect 219433 402462 240212 402464
rect 219433 402459 219499 402462
rect 213361 401978 213427 401981
rect 213361 401976 240212 401978
rect 213361 401920 213366 401976
rect 213422 401920 240212 401976
rect 213361 401918 240212 401920
rect 213361 401915 213427 401918
rect 280337 401706 280403 401709
rect 279956 401704 280403 401706
rect 279956 401648 280342 401704
rect 280398 401648 280403 401704
rect 279956 401646 280403 401648
rect 280337 401643 280403 401646
rect 239489 401570 239555 401573
rect 240174 401570 240180 401572
rect 239489 401568 240180 401570
rect 239489 401512 239494 401568
rect 239550 401512 240180 401568
rect 239489 401510 240180 401512
rect 239489 401507 239555 401510
rect 240174 401508 240180 401510
rect 240244 401508 240250 401572
rect 207289 401434 207355 401437
rect 207289 401432 240212 401434
rect 207289 401376 207294 401432
rect 207350 401376 240212 401432
rect 207289 401374 240212 401376
rect 207289 401371 207355 401374
rect 201217 400890 201283 400893
rect 201217 400888 240212 400890
rect 201217 400832 201222 400888
rect 201278 400832 240212 400888
rect 201217 400830 240212 400832
rect 201217 400827 201283 400830
rect 195145 400346 195211 400349
rect 280245 400346 280311 400349
rect 195145 400344 240212 400346
rect 195145 400288 195150 400344
rect 195206 400288 240212 400344
rect 195145 400286 240212 400288
rect 279956 400344 280311 400346
rect 279956 400288 280250 400344
rect 280306 400288 280311 400344
rect 279956 400286 280311 400288
rect 195145 400283 195211 400286
rect 280245 400283 280311 400286
rect 215937 399802 216003 399805
rect 215937 399800 240212 399802
rect 215937 399744 215942 399800
rect 215998 399744 240212 399800
rect 215937 399742 240212 399744
rect 215937 399739 216003 399742
rect 183001 399258 183067 399261
rect 183001 399256 240212 399258
rect 183001 399200 183006 399256
rect 183062 399200 240212 399256
rect 183001 399198 240212 399200
rect 183001 399195 183067 399198
rect 280153 398986 280219 398989
rect 279956 398984 280219 398986
rect 279956 398928 280158 398984
rect 280214 398928 280219 398984
rect 279956 398926 280219 398928
rect 280153 398923 280219 398926
rect 176929 398714 176995 398717
rect 176929 398712 240212 398714
rect 176929 398656 176934 398712
rect 176990 398656 240212 398712
rect 176929 398654 240212 398656
rect 176929 398651 176995 398654
rect 170857 398170 170923 398173
rect 170857 398168 240212 398170
rect 170857 398112 170862 398168
rect 170918 398112 240212 398168
rect 170857 398110 240212 398112
rect 170857 398107 170923 398110
rect 231117 397626 231183 397629
rect 280061 397626 280127 397629
rect 231117 397624 240212 397626
rect -960 397490 480 397580
rect 231117 397568 231122 397624
rect 231178 397568 240212 397624
rect 231117 397566 240212 397568
rect 279956 397624 280127 397626
rect 279956 397568 280066 397624
rect 280122 397568 280127 397624
rect 279956 397566 280127 397568
rect 231117 397563 231183 397566
rect 280061 397563 280127 397566
rect 173198 397490 173204 397492
rect -960 397430 173204 397490
rect -960 397340 480 397430
rect 173198 397428 173204 397430
rect 173268 397428 173274 397492
rect 158713 397082 158779 397085
rect 158713 397080 240212 397082
rect 158713 397024 158718 397080
rect 158774 397024 240212 397080
rect 158713 397022 240212 397024
rect 158713 397019 158779 397022
rect 152641 396538 152707 396541
rect 152641 396536 240212 396538
rect 152641 396480 152646 396536
rect 152702 396480 240212 396536
rect 152641 396478 240212 396480
rect 152641 396475 152707 396478
rect 279550 396204 279556 396268
rect 279620 396204 279626 396268
rect 146569 395994 146635 395997
rect 146569 395992 240212 395994
rect 146569 395936 146574 395992
rect 146630 395936 240212 395992
rect 146569 395934 240212 395936
rect 146569 395931 146635 395934
rect 282821 395722 282887 395725
rect 280110 395720 282887 395722
rect 280110 395664 282826 395720
rect 282882 395664 282887 395720
rect 280110 395662 282887 395664
rect 280110 395586 280170 395662
rect 282821 395659 282887 395662
rect 279926 395526 280170 395586
rect 140497 395450 140563 395453
rect 140497 395448 240212 395450
rect 140497 395392 140502 395448
rect 140558 395392 240212 395448
rect 140497 395390 240212 395392
rect 140497 395387 140563 395390
rect 134425 394906 134491 394909
rect 134425 394904 240212 394906
rect 134425 394848 134430 394904
rect 134486 394848 240212 394904
rect 279926 394876 279986 395526
rect 134425 394846 240212 394848
rect 134425 394843 134491 394846
rect 128353 394362 128419 394365
rect 128353 394360 240212 394362
rect 128353 394304 128358 394360
rect 128414 394304 240212 394360
rect 128353 394302 240212 394304
rect 128353 394299 128419 394302
rect 122281 393818 122347 393821
rect 122281 393816 240212 393818
rect 122281 393760 122286 393816
rect 122342 393760 240212 393816
rect 122281 393758 240212 393760
rect 122281 393755 122347 393758
rect 281809 393546 281875 393549
rect 279956 393544 281875 393546
rect 279956 393488 281814 393544
rect 281870 393488 281875 393544
rect 279956 393486 281875 393488
rect 281809 393483 281875 393486
rect 211797 393274 211863 393277
rect 211797 393272 240212 393274
rect 211797 393216 211802 393272
rect 211858 393216 240212 393272
rect 211797 393214 240212 393216
rect 211797 393211 211863 393214
rect 226977 392730 227043 392733
rect 226977 392728 240212 392730
rect 226977 392672 226982 392728
rect 227038 392672 240212 392728
rect 226977 392670 240212 392672
rect 226977 392667 227043 392670
rect 104065 392186 104131 392189
rect 287462 392186 287468 392188
rect 104065 392184 240212 392186
rect 104065 392128 104070 392184
rect 104126 392128 240212 392184
rect 104065 392126 240212 392128
rect 279956 392126 287468 392186
rect 104065 392123 104131 392126
rect 287462 392124 287468 392126
rect 287532 392124 287538 392188
rect 97993 391642 98059 391645
rect 97993 391640 240212 391642
rect 97993 391584 97998 391640
rect 98054 391584 240212 391640
rect 583520 391628 584960 391868
rect 97993 391582 240212 391584
rect 97993 391579 98059 391582
rect 91921 391098 91987 391101
rect 91921 391096 240212 391098
rect 91921 391040 91926 391096
rect 91982 391040 240212 391096
rect 91921 391038 240212 391040
rect 91921 391035 91987 391038
rect 287646 390826 287652 390828
rect 279956 390766 287652 390826
rect 287646 390764 287652 390766
rect 287716 390764 287722 390828
rect 85849 390554 85915 390557
rect 85849 390552 240212 390554
rect 85849 390496 85854 390552
rect 85910 390496 240212 390552
rect 85849 390494 240212 390496
rect 85849 390491 85915 390494
rect 79777 390010 79843 390013
rect 79777 390008 240212 390010
rect 79777 389952 79782 390008
rect 79838 389952 240212 390008
rect 79777 389950 240212 389952
rect 79777 389947 79843 389950
rect 73705 389466 73771 389469
rect 280153 389466 280219 389469
rect 73705 389464 240212 389466
rect 73705 389408 73710 389464
rect 73766 389408 240212 389464
rect 73705 389406 240212 389408
rect 279956 389464 280219 389466
rect 279956 389408 280158 389464
rect 280214 389408 280219 389464
rect 279956 389406 280219 389408
rect 73705 389403 73771 389406
rect 280153 389403 280219 389406
rect 126329 388922 126395 388925
rect 126329 388920 240212 388922
rect 126329 388864 126334 388920
rect 126390 388864 240212 388920
rect 126329 388862 240212 388864
rect 126329 388859 126395 388862
rect 111057 388378 111123 388381
rect 111057 388376 240212 388378
rect 111057 388320 111062 388376
rect 111118 388320 240212 388376
rect 111057 388318 240212 388320
rect 111057 388315 111123 388318
rect 283097 388106 283163 388109
rect 279956 388104 283163 388106
rect 279956 388048 283102 388104
rect 283158 388048 283163 388104
rect 279956 388046 283163 388048
rect 283097 388043 283163 388046
rect 116577 387834 116643 387837
rect 116577 387832 240212 387834
rect 116577 387776 116582 387832
rect 116638 387776 240212 387832
rect 116577 387774 240212 387776
rect 116577 387771 116643 387774
rect 119429 387290 119495 387293
rect 119429 387288 240212 387290
rect 119429 387232 119434 387288
rect 119490 387232 240212 387288
rect 119429 387230 240212 387232
rect 119429 387227 119495 387230
rect 111241 386746 111307 386749
rect 288893 386746 288959 386749
rect 111241 386744 240212 386746
rect 111241 386688 111246 386744
rect 111302 386688 240212 386744
rect 111241 386686 240212 386688
rect 279956 386744 288959 386746
rect 279956 386688 288898 386744
rect 288954 386688 288959 386744
rect 279956 386686 288959 386688
rect 111241 386683 111307 386686
rect 288893 386683 288959 386686
rect 115197 386202 115263 386205
rect 115197 386200 240212 386202
rect 115197 386144 115202 386200
rect 115258 386144 240212 386200
rect 115197 386142 240212 386144
rect 115197 386139 115263 386142
rect 111425 385658 111491 385661
rect 111425 385656 240212 385658
rect 111425 385600 111430 385656
rect 111486 385600 240212 385656
rect 111425 385598 240212 385600
rect 111425 385595 111491 385598
rect 284477 385386 284543 385389
rect 279956 385384 284543 385386
rect 279956 385328 284482 385384
rect 284538 385328 284543 385384
rect 279956 385326 284543 385328
rect 284477 385323 284543 385326
rect 117957 385114 118023 385117
rect 117957 385112 240212 385114
rect 117957 385056 117962 385112
rect 118018 385056 240212 385112
rect 117957 385054 240212 385056
rect 117957 385051 118023 385054
rect 112621 384570 112687 384573
rect 112621 384568 240212 384570
rect -960 384284 480 384524
rect 112621 384512 112626 384568
rect 112682 384512 240212 384568
rect 112621 384510 240212 384512
rect 112621 384507 112687 384510
rect 237373 384026 237439 384029
rect 280245 384026 280311 384029
rect 237373 384024 240212 384026
rect 237373 383968 237378 384024
rect 237434 383968 240212 384024
rect 237373 383966 240212 383968
rect 279956 384024 280311 384026
rect 279956 383968 280250 384024
rect 280306 383968 280311 384024
rect 279956 383966 280311 383968
rect 237373 383963 237439 383966
rect 280245 383963 280311 383966
rect 237373 383482 237439 383485
rect 237373 383480 240212 383482
rect 237373 383424 237378 383480
rect 237434 383424 240212 383480
rect 237373 383422 240212 383424
rect 237373 383419 237439 383422
rect 237465 382938 237531 382941
rect 237465 382936 240212 382938
rect 237465 382880 237470 382936
rect 237526 382880 240212 382936
rect 237465 382878 240212 382880
rect 237465 382875 237531 382878
rect 281717 382666 281783 382669
rect 279956 382664 281783 382666
rect 279956 382608 281722 382664
rect 281778 382608 281783 382664
rect 279956 382606 281783 382608
rect 281717 382603 281783 382606
rect 237373 382394 237439 382397
rect 237373 382392 240212 382394
rect 237373 382336 237378 382392
rect 237434 382336 240212 382392
rect 237373 382334 240212 382336
rect 237373 382331 237439 382334
rect 237557 381850 237623 381853
rect 237557 381848 240212 381850
rect 237557 381792 237562 381848
rect 237618 381792 240212 381848
rect 237557 381790 240212 381792
rect 237557 381787 237623 381790
rect 237373 381306 237439 381309
rect 281625 381306 281691 381309
rect 237373 381304 240212 381306
rect 237373 381248 237378 381304
rect 237434 381248 240212 381304
rect 237373 381246 240212 381248
rect 279956 381304 281691 381306
rect 279956 381248 281630 381304
rect 281686 381248 281691 381304
rect 279956 381246 281691 381248
rect 237373 381243 237439 381246
rect 281625 381243 281691 381246
rect 237373 380762 237439 380765
rect 237373 380760 240212 380762
rect 237373 380704 237378 380760
rect 237434 380704 240212 380760
rect 237373 380702 240212 380704
rect 237373 380699 237439 380702
rect 114001 380218 114067 380221
rect 114001 380216 240212 380218
rect 114001 380160 114006 380216
rect 114062 380160 240212 380216
rect 114001 380158 240212 380160
rect 114001 380155 114067 380158
rect 281533 379946 281599 379949
rect 279956 379944 281599 379946
rect 279956 379888 281538 379944
rect 281594 379888 281599 379944
rect 279956 379886 281599 379888
rect 281533 379883 281599 379886
rect 113817 379674 113883 379677
rect 113817 379672 240212 379674
rect 113817 379616 113822 379672
rect 113878 379616 240212 379672
rect 113817 379614 240212 379616
rect 113817 379611 113883 379614
rect 111333 379130 111399 379133
rect 111333 379128 240212 379130
rect 111333 379072 111338 379128
rect 111394 379072 240212 379128
rect 111333 379070 240212 379072
rect 111333 379067 111399 379070
rect 120717 378586 120783 378589
rect 280429 378586 280495 378589
rect 120717 378584 240212 378586
rect 120717 378528 120722 378584
rect 120778 378528 240212 378584
rect 120717 378526 240212 378528
rect 279956 378584 280495 378586
rect 279956 378528 280434 378584
rect 280490 378528 280495 378584
rect 279956 378526 280495 378528
rect 120717 378523 120783 378526
rect 280429 378523 280495 378526
rect 580257 378450 580323 378453
rect 583520 378450 584960 378540
rect 580257 378448 584960 378450
rect 580257 378392 580262 378448
rect 580318 378392 584960 378448
rect 580257 378390 584960 378392
rect 580257 378387 580323 378390
rect 583520 378300 584960 378390
rect 237741 378042 237807 378045
rect 237741 378040 240212 378042
rect 237741 377984 237746 378040
rect 237802 377984 240212 378040
rect 237741 377982 240212 377984
rect 237741 377979 237807 377982
rect 237557 377498 237623 377501
rect 237557 377496 240212 377498
rect 237557 377440 237562 377496
rect 237618 377440 240212 377496
rect 237557 377438 240212 377440
rect 237557 377435 237623 377438
rect 284845 377226 284911 377229
rect 279956 377224 284911 377226
rect 279956 377168 284850 377224
rect 284906 377168 284911 377224
rect 279956 377166 284911 377168
rect 284845 377163 284911 377166
rect 237373 376954 237439 376957
rect 237373 376952 240212 376954
rect 237373 376896 237378 376952
rect 237434 376896 240212 376952
rect 237373 376894 240212 376896
rect 237373 376891 237439 376894
rect 237557 376410 237623 376413
rect 237557 376408 240212 376410
rect 237557 376352 237562 376408
rect 237618 376352 240212 376408
rect 237557 376350 240212 376352
rect 237557 376347 237623 376350
rect 237373 375866 237439 375869
rect 284569 375866 284635 375869
rect 237373 375864 240212 375866
rect 237373 375808 237378 375864
rect 237434 375808 240212 375864
rect 237373 375806 240212 375808
rect 279956 375864 284635 375866
rect 279956 375808 284574 375864
rect 284630 375808 284635 375864
rect 279956 375806 284635 375808
rect 237373 375803 237439 375806
rect 284569 375803 284635 375806
rect 237373 375322 237439 375325
rect 237373 375320 240212 375322
rect 237373 375264 237378 375320
rect 237434 375264 240212 375320
rect 237373 375262 240212 375264
rect 237373 375259 237439 375262
rect 140037 374778 140103 374781
rect 140037 374776 240212 374778
rect 140037 374720 140042 374776
rect 140098 374720 240212 374776
rect 140037 374718 240212 374720
rect 140037 374715 140103 374718
rect 284385 374506 284451 374509
rect 279956 374504 284451 374506
rect 279956 374448 284390 374504
rect 284446 374448 284451 374504
rect 279956 374446 284451 374448
rect 284385 374443 284451 374446
rect 237373 374234 237439 374237
rect 237373 374232 240212 374234
rect 237373 374176 237378 374232
rect 237434 374176 240212 374232
rect 237373 374174 240212 374176
rect 237373 374171 237439 374174
rect 122097 373690 122163 373693
rect 122097 373688 240212 373690
rect 122097 373632 122102 373688
rect 122158 373632 240212 373688
rect 122097 373630 240212 373632
rect 122097 373627 122163 373630
rect 123661 373146 123727 373149
rect 280337 373146 280403 373149
rect 123661 373144 240212 373146
rect 123661 373088 123666 373144
rect 123722 373088 240212 373144
rect 123661 373086 240212 373088
rect 279956 373144 280403 373146
rect 279956 373088 280342 373144
rect 280398 373088 280403 373144
rect 279956 373086 280403 373088
rect 123661 373083 123727 373086
rect 280337 373083 280403 373086
rect 127709 372602 127775 372605
rect 127709 372600 240212 372602
rect 127709 372544 127714 372600
rect 127770 372544 240212 372600
rect 127709 372542 240212 372544
rect 127709 372539 127775 372542
rect 130377 372058 130443 372061
rect 130377 372056 240212 372058
rect 130377 372000 130382 372056
rect 130438 372000 240212 372056
rect 130377 371998 240212 372000
rect 130377 371995 130443 371998
rect 284293 371786 284359 371789
rect 279956 371784 284359 371786
rect 279956 371728 284298 371784
rect 284354 371728 284359 371784
rect 279956 371726 284359 371728
rect 284293 371723 284359 371726
rect 237373 371514 237439 371517
rect 237373 371512 240212 371514
rect -960 371378 480 371468
rect 237373 371456 237378 371512
rect 237434 371456 240212 371512
rect 237373 371454 240212 371456
rect 237373 371451 237439 371454
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 237373 370970 237439 370973
rect 237373 370968 240212 370970
rect 237373 370912 237378 370968
rect 237434 370912 240212 370968
rect 237373 370910 240212 370912
rect 237373 370907 237439 370910
rect 134517 370426 134583 370429
rect 284661 370426 284727 370429
rect 134517 370424 240212 370426
rect 134517 370368 134522 370424
rect 134578 370368 240212 370424
rect 134517 370366 240212 370368
rect 279956 370424 284727 370426
rect 279956 370368 284666 370424
rect 284722 370368 284727 370424
rect 279956 370366 284727 370368
rect 134517 370363 134583 370366
rect 284661 370363 284727 370366
rect 231577 369882 231643 369885
rect 231577 369880 240212 369882
rect 231577 369824 231582 369880
rect 231638 369824 240212 369880
rect 231577 369822 240212 369824
rect 231577 369819 231643 369822
rect 232773 369338 232839 369341
rect 232773 369336 240212 369338
rect 232773 369280 232778 369336
rect 232834 369280 240212 369336
rect 232773 369278 240212 369280
rect 232773 369275 232839 369278
rect 282821 369066 282887 369069
rect 279956 369064 282887 369066
rect 279956 369008 282826 369064
rect 282882 369008 282887 369064
rect 279956 369006 282887 369008
rect 282821 369003 282887 369006
rect 235574 368732 235580 368796
rect 235644 368794 235650 368796
rect 235644 368734 240212 368794
rect 235644 368732 235650 368734
rect 235073 368250 235139 368253
rect 235073 368248 240212 368250
rect 235073 368192 235078 368248
rect 235134 368192 240212 368248
rect 235073 368190 240212 368192
rect 235073 368187 235139 368190
rect 50613 367706 50679 367709
rect 231577 367706 231643 367709
rect 50613 367704 231643 367706
rect 50613 367648 50618 367704
rect 50674 367648 231582 367704
rect 231638 367648 231643 367704
rect 50613 367646 231643 367648
rect 50613 367643 50679 367646
rect 231577 367643 231643 367646
rect 235717 367706 235783 367709
rect 280521 367706 280587 367709
rect 235717 367704 240212 367706
rect 235717 367648 235722 367704
rect 235778 367648 240212 367704
rect 235717 367646 240212 367648
rect 279956 367704 280587 367706
rect 279956 367648 280526 367704
rect 280582 367648 280587 367704
rect 279956 367646 280587 367648
rect 235717 367643 235783 367646
rect 280521 367643 280587 367646
rect 235809 367162 235875 367165
rect 235809 367160 240212 367162
rect 235809 367104 235814 367160
rect 235870 367104 240212 367160
rect 235809 367102 240212 367104
rect 235809 367099 235875 367102
rect 231301 366618 231367 366621
rect 231301 366616 240212 366618
rect 231301 366560 231306 366616
rect 231362 366560 240212 366616
rect 231301 366558 240212 366560
rect 231301 366555 231367 366558
rect 283281 366346 283347 366349
rect 279956 366344 283347 366346
rect 279956 366288 283286 366344
rect 283342 366288 283347 366344
rect 279956 366286 283347 366288
rect 283281 366283 283347 366286
rect 238017 366074 238083 366077
rect 238017 366072 240212 366074
rect 238017 366016 238022 366072
rect 238078 366016 240212 366072
rect 238017 366014 240212 366016
rect 238017 366011 238083 366014
rect 235165 365530 235231 365533
rect 235165 365528 240212 365530
rect 235165 365472 235170 365528
rect 235226 365472 240212 365528
rect 235165 365470 240212 365472
rect 235165 365467 235231 365470
rect 580206 365060 580212 365124
rect 580276 365122 580282 365124
rect 583520 365122 584960 365212
rect 580276 365062 584960 365122
rect 580276 365060 580282 365062
rect 8109 364986 8175 364989
rect 231209 364986 231275 364989
rect 8109 364984 231275 364986
rect 8109 364928 8114 364984
rect 8170 364928 231214 364984
rect 231270 364928 231275 364984
rect 8109 364926 231275 364928
rect 8109 364923 8175 364926
rect 231209 364923 231275 364926
rect 235441 364986 235507 364989
rect 281993 364986 282059 364989
rect 235441 364984 240212 364986
rect 235441 364928 235446 364984
rect 235502 364928 240212 364984
rect 235441 364926 240212 364928
rect 279956 364984 282059 364986
rect 279956 364928 281998 364984
rect 282054 364928 282059 364984
rect 583520 364972 584960 365062
rect 279956 364926 282059 364928
rect 235441 364923 235507 364926
rect 281993 364923 282059 364926
rect 228541 364442 228607 364445
rect 228541 364440 240212 364442
rect 228541 364384 228546 364440
rect 228602 364384 240212 364440
rect 228541 364382 240212 364384
rect 228541 364379 228607 364382
rect 227253 363898 227319 363901
rect 227253 363896 240212 363898
rect 227253 363840 227258 363896
rect 227314 363840 240212 363896
rect 227253 363838 240212 363840
rect 227253 363835 227319 363838
rect 283373 363626 283439 363629
rect 279956 363624 283439 363626
rect 279956 363568 283378 363624
rect 283434 363568 283439 363624
rect 279956 363566 283439 363568
rect 283373 363563 283439 363566
rect 228633 363354 228699 363357
rect 228633 363352 240212 363354
rect 228633 363296 228638 363352
rect 228694 363296 240212 363352
rect 228633 363294 240212 363296
rect 228633 363291 228699 363294
rect 236453 362810 236519 362813
rect 236453 362808 240212 362810
rect 236453 362752 236458 362808
rect 236514 362752 240212 362808
rect 236453 362750 240212 362752
rect 236453 362747 236519 362750
rect 239673 362266 239739 362269
rect 280613 362266 280679 362269
rect 239673 362264 240212 362266
rect 239673 362208 239678 362264
rect 239734 362208 240212 362264
rect 239673 362206 240212 362208
rect 279956 362264 280679 362266
rect 279956 362208 280618 362264
rect 280674 362208 280679 362264
rect 279956 362206 280679 362208
rect 239673 362203 239739 362206
rect 280613 362203 280679 362206
rect 230105 361722 230171 361725
rect 230105 361720 240212 361722
rect 230105 361664 230110 361720
rect 230166 361664 240212 361720
rect 230105 361662 240212 361664
rect 230105 361659 230171 361662
rect 239581 361178 239647 361181
rect 239581 361176 240212 361178
rect 239581 361120 239586 361176
rect 239642 361120 240212 361176
rect 239581 361118 240212 361120
rect 239581 361115 239647 361118
rect 281901 360906 281967 360909
rect 279956 360904 281967 360906
rect 279956 360848 281906 360904
rect 281962 360848 281967 360904
rect 279956 360846 281967 360848
rect 281901 360843 281967 360846
rect 236545 360634 236611 360637
rect 236545 360632 240212 360634
rect 236545 360576 236550 360632
rect 236606 360576 240212 360632
rect 236545 360574 240212 360576
rect 236545 360571 236611 360574
rect 236637 360090 236703 360093
rect 236637 360088 240212 360090
rect 236637 360032 236642 360088
rect 236698 360032 240212 360088
rect 236637 360030 240212 360032
rect 236637 360027 236703 360030
rect 236821 359546 236887 359549
rect 282821 359546 282887 359549
rect 236821 359544 240212 359546
rect 236821 359488 236826 359544
rect 236882 359488 240212 359544
rect 236821 359486 240212 359488
rect 279956 359544 282887 359546
rect 279956 359488 282826 359544
rect 282882 359488 282887 359544
rect 279956 359486 282887 359488
rect 236821 359483 236887 359486
rect 282821 359483 282887 359486
rect 237097 359002 237163 359005
rect 237097 359000 240212 359002
rect 237097 358944 237102 359000
rect 237158 358944 240212 359000
rect 237097 358942 240212 358944
rect 237097 358939 237163 358942
rect -960 358458 480 358548
rect 235390 358458 235396 358460
rect -960 358398 235396 358458
rect -960 358308 480 358398
rect 235390 358396 235396 358398
rect 235460 358396 235466 358460
rect 236913 358458 236979 358461
rect 236913 358456 240212 358458
rect 236913 358400 236918 358456
rect 236974 358400 240212 358456
rect 236913 358398 240212 358400
rect 236913 358395 236979 358398
rect 280705 358186 280771 358189
rect 279956 358184 280771 358186
rect 279956 358128 280710 358184
rect 280766 358128 280771 358184
rect 279956 358126 280771 358128
rect 280705 358123 280771 358126
rect 227345 357914 227411 357917
rect 227345 357912 240212 357914
rect 227345 357856 227350 357912
rect 227406 357856 240212 357912
rect 227345 357854 240212 357856
rect 227345 357851 227411 357854
rect 228817 357370 228883 357373
rect 228817 357368 240212 357370
rect 228817 357312 228822 357368
rect 228878 357312 240212 357368
rect 228817 357310 240212 357312
rect 228817 357307 228883 357310
rect 227529 356826 227595 356829
rect 282821 356826 282887 356829
rect 227529 356824 240212 356826
rect 227529 356768 227534 356824
rect 227590 356768 240212 356824
rect 227529 356766 240212 356768
rect 279956 356824 282887 356826
rect 279956 356768 282826 356824
rect 282882 356768 282887 356824
rect 279956 356766 282887 356768
rect 227529 356763 227595 356766
rect 282821 356763 282887 356766
rect 230197 356282 230263 356285
rect 230197 356280 240212 356282
rect 230197 356224 230202 356280
rect 230258 356224 240212 356280
rect 230197 356222 240212 356224
rect 230197 356219 230263 356222
rect 232865 355738 232931 355741
rect 232865 355736 240212 355738
rect 232865 355680 232870 355736
rect 232926 355680 240212 355736
rect 232865 355678 240212 355680
rect 232865 355675 232931 355678
rect 280889 355466 280955 355469
rect 279956 355464 280955 355466
rect 279956 355408 280894 355464
rect 280950 355408 280955 355464
rect 279956 355406 280955 355408
rect 280889 355403 280955 355406
rect 227437 355194 227503 355197
rect 227437 355192 240212 355194
rect 227437 355136 227442 355192
rect 227498 355136 240212 355192
rect 227437 355134 240212 355136
rect 227437 355131 227503 355134
rect 235349 354650 235415 354653
rect 235349 354648 240212 354650
rect 235349 354592 235354 354648
rect 235410 354592 240212 354648
rect 235349 354590 240212 354592
rect 235349 354587 235415 354590
rect 236729 354106 236795 354109
rect 282821 354106 282887 354109
rect 236729 354104 240212 354106
rect 236729 354048 236734 354104
rect 236790 354048 240212 354104
rect 236729 354046 240212 354048
rect 279956 354104 282887 354106
rect 279956 354048 282826 354104
rect 282882 354048 282887 354104
rect 279956 354046 282887 354048
rect 236729 354043 236795 354046
rect 282821 354043 282887 354046
rect 235257 353562 235323 353565
rect 235257 353560 240212 353562
rect 235257 353504 235262 353560
rect 235318 353504 240212 353560
rect 235257 353502 240212 353504
rect 235257 353499 235323 353502
rect 235533 353018 235599 353021
rect 235533 353016 240212 353018
rect 235533 352960 235538 353016
rect 235594 352960 240212 353016
rect 235533 352958 240212 352960
rect 235533 352955 235599 352958
rect 287053 352746 287119 352749
rect 279956 352744 287119 352746
rect 279956 352688 287058 352744
rect 287114 352688 287119 352744
rect 279956 352686 287119 352688
rect 287053 352683 287119 352686
rect 237189 352474 237255 352477
rect 237189 352472 240212 352474
rect 237189 352416 237194 352472
rect 237250 352416 240212 352472
rect 237189 352414 240212 352416
rect 237189 352411 237255 352414
rect 234981 351930 235047 351933
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 234981 351928 240212 351930
rect 234981 351872 234986 351928
rect 235042 351872 240212 351928
rect 234981 351870 240212 351872
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 234981 351867 235047 351870
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 235901 351386 235967 351389
rect 283465 351386 283531 351389
rect 235901 351384 240212 351386
rect 235901 351328 235906 351384
rect 235962 351328 240212 351384
rect 235901 351326 240212 351328
rect 279956 351384 283531 351386
rect 279956 351328 283470 351384
rect 283526 351328 283531 351384
rect 279956 351326 283531 351328
rect 235901 351323 235967 351326
rect 283465 351323 283531 351326
rect 68829 351114 68895 351117
rect 227069 351114 227135 351117
rect 68829 351112 227135 351114
rect 68829 351056 68834 351112
rect 68890 351056 227074 351112
rect 227130 351056 227135 351112
rect 68829 351054 227135 351056
rect 68829 351051 68895 351054
rect 227069 351051 227135 351054
rect 237005 350842 237071 350845
rect 237005 350840 240212 350842
rect 237005 350784 237010 350840
rect 237066 350784 240212 350840
rect 237005 350782 240212 350784
rect 237005 350779 237071 350782
rect 231485 350298 231551 350301
rect 231485 350296 240212 350298
rect 231485 350240 231490 350296
rect 231546 350240 240212 350296
rect 231485 350238 240212 350240
rect 231485 350235 231551 350238
rect 283557 350026 283623 350029
rect 279956 350024 283623 350026
rect 279956 349968 283562 350024
rect 283618 349968 283623 350024
rect 279956 349966 283623 349968
rect 283557 349963 283623 349966
rect 159357 349754 159423 349757
rect 159357 349752 240212 349754
rect 159357 349696 159362 349752
rect 159418 349696 240212 349752
rect 159357 349694 240212 349696
rect 159357 349691 159423 349694
rect 5257 349210 5323 349213
rect 5257 349208 240212 349210
rect 5257 349152 5262 349208
rect 5318 349152 240212 349208
rect 5257 349150 240212 349152
rect 5257 349147 5323 349150
rect 210417 348666 210483 348669
rect 282821 348666 282887 348669
rect 210417 348664 240212 348666
rect 210417 348608 210422 348664
rect 210478 348608 240212 348664
rect 210417 348606 240212 348608
rect 279956 348664 282887 348666
rect 279956 348608 282826 348664
rect 282882 348608 282887 348664
rect 279956 348606 282887 348608
rect 210417 348603 210483 348606
rect 282821 348603 282887 348606
rect 6453 348122 6519 348125
rect 6453 348120 240212 348122
rect 6453 348064 6458 348120
rect 6514 348064 240212 348120
rect 6453 348062 240212 348064
rect 6453 348059 6519 348062
rect 237925 347716 237991 347717
rect 237925 347714 237972 347716
rect 237880 347712 237972 347714
rect 237880 347656 237930 347712
rect 237880 347654 237972 347656
rect 237925 347652 237972 347654
rect 238036 347652 238042 347716
rect 237925 347651 237991 347652
rect 216121 347578 216187 347581
rect 216121 347576 240212 347578
rect 216121 347520 216126 347576
rect 216182 347520 240212 347576
rect 216121 347518 240212 347520
rect 216121 347515 216187 347518
rect 285029 347306 285095 347309
rect 279956 347304 285095 347306
rect 279956 347248 285034 347304
rect 285090 347248 285095 347304
rect 279956 347246 285095 347248
rect 285029 347243 285095 347246
rect 69974 347108 69980 347172
rect 70044 347170 70050 347172
rect 237414 347170 237420 347172
rect 70044 347110 237420 347170
rect 70044 347108 70050 347110
rect 237414 347108 237420 347110
rect 237484 347108 237490 347172
rect 163497 347034 163563 347037
rect 163497 347032 240212 347034
rect 163497 346976 163502 347032
rect 163558 346976 240212 347032
rect 163497 346974 240212 346976
rect 163497 346971 163563 346974
rect 227161 346490 227227 346493
rect 227161 346488 240212 346490
rect 227161 346432 227166 346488
rect 227222 346432 240212 346488
rect 227161 346430 240212 346432
rect 227161 346427 227227 346430
rect 199377 345946 199443 345949
rect 283189 345946 283255 345949
rect 199377 345944 240212 345946
rect 199377 345888 199382 345944
rect 199438 345888 240212 345944
rect 199377 345886 240212 345888
rect 279956 345944 283255 345946
rect 279956 345888 283194 345944
rect 283250 345888 283255 345944
rect 279956 345886 283255 345888
rect 199377 345883 199443 345886
rect 283189 345883 283255 345886
rect -960 345402 480 345492
rect 146937 345402 147003 345405
rect -960 345342 6930 345402
rect -960 345252 480 345342
rect 6870 345266 6930 345342
rect 146937 345400 240212 345402
rect 146937 345344 146942 345400
rect 146998 345344 240212 345400
rect 146937 345342 240212 345344
rect 146937 345339 147003 345342
rect 147070 345266 147076 345268
rect 6870 345206 147076 345266
rect 147070 345204 147076 345206
rect 147140 345204 147146 345268
rect 69606 344932 69612 344996
rect 69676 344994 69682 344996
rect 225597 344994 225663 344997
rect 69676 344992 225663 344994
rect 69676 344936 225602 344992
rect 225658 344936 225663 344992
rect 69676 344934 225663 344936
rect 69676 344932 69682 344934
rect 225597 344931 225663 344934
rect 202137 344858 202203 344861
rect 202137 344856 240212 344858
rect 202137 344800 202142 344856
rect 202198 344800 240212 344856
rect 202137 344798 240212 344800
rect 202137 344795 202203 344798
rect 62982 344660 62988 344724
rect 63052 344722 63058 344724
rect 223062 344722 223068 344724
rect 63052 344662 223068 344722
rect 63052 344660 63058 344662
rect 223062 344660 223068 344662
rect 223132 344660 223138 344724
rect 67449 344586 67515 344589
rect 228449 344586 228515 344589
rect 282821 344586 282887 344589
rect 67449 344584 228515 344586
rect 67449 344528 67454 344584
rect 67510 344528 228454 344584
rect 228510 344528 228515 344584
rect 67449 344526 228515 344528
rect 279956 344584 282887 344586
rect 279956 344528 282826 344584
rect 282882 344528 282887 344584
rect 279956 344526 282887 344528
rect 67449 344523 67515 344526
rect 228449 344523 228515 344526
rect 282821 344523 282887 344526
rect 63166 344388 63172 344452
rect 63236 344450 63242 344452
rect 225413 344450 225479 344453
rect 63236 344448 225479 344450
rect 63236 344392 225418 344448
rect 225474 344392 225479 344448
rect 63236 344390 225479 344392
rect 63236 344388 63242 344390
rect 225413 344387 225479 344390
rect 217317 344314 217383 344317
rect 217317 344312 240212 344314
rect 217317 344256 217322 344312
rect 217378 344256 240212 344312
rect 217317 344254 240212 344256
rect 217317 344251 217383 344254
rect 62021 344178 62087 344181
rect 216673 344178 216739 344181
rect 62021 344176 216739 344178
rect 62021 344120 62026 344176
rect 62082 344120 216678 344176
rect 216734 344120 216739 344176
rect 62021 344118 216739 344120
rect 62021 344115 62087 344118
rect 216673 344115 216739 344118
rect 63350 343980 63356 344044
rect 63420 344042 63426 344044
rect 225781 344042 225847 344045
rect 63420 344040 225847 344042
rect 63420 343984 225786 344040
rect 225842 343984 225847 344040
rect 63420 343982 225847 343984
rect 63420 343980 63426 343982
rect 225781 343979 225847 343982
rect 222837 343770 222903 343773
rect 222837 343768 240212 343770
rect 222837 343712 222842 343768
rect 222898 343712 240212 343768
rect 222837 343710 240212 343712
rect 222837 343707 222903 343710
rect 61745 343634 61811 343637
rect 66161 343634 66227 343637
rect 61745 343632 66227 343634
rect 61745 343576 61750 343632
rect 61806 343576 66166 343632
rect 66222 343576 66227 343632
rect 61745 343574 66227 343576
rect 61745 343571 61811 343574
rect 66161 343571 66227 343574
rect 64689 343498 64755 343501
rect 80329 343498 80395 343501
rect 64689 343496 80395 343498
rect 64689 343440 64694 343496
rect 64750 343440 80334 343496
rect 80390 343440 80395 343496
rect 64689 343438 80395 343440
rect 64689 343435 64755 343438
rect 80329 343435 80395 343438
rect 66069 343362 66135 343365
rect 85573 343362 85639 343365
rect 66069 343360 85639 343362
rect 66069 343304 66074 343360
rect 66130 343304 85578 343360
rect 85634 343304 85639 343360
rect 66069 343302 85639 343304
rect 66069 343299 66135 343302
rect 85573 343299 85639 343302
rect 61929 343226 61995 343229
rect 81985 343226 82051 343229
rect 61929 343224 82051 343226
rect 61929 343168 61934 343224
rect 61990 343168 81990 343224
rect 82046 343168 82051 343224
rect 61929 343166 82051 343168
rect 61929 343163 61995 343166
rect 81985 343163 82051 343166
rect 174537 343226 174603 343229
rect 284753 343226 284819 343229
rect 174537 343224 240212 343226
rect 174537 343168 174542 343224
rect 174598 343168 240212 343224
rect 174537 343166 240212 343168
rect 279956 343224 284819 343226
rect 279956 343168 284758 343224
rect 284814 343168 284819 343224
rect 279956 343166 284819 343168
rect 174537 343163 174603 343166
rect 284753 343163 284819 343166
rect 60641 343090 60707 343093
rect 88609 343090 88675 343093
rect 60641 343088 88675 343090
rect 60641 343032 60646 343088
rect 60702 343032 88614 343088
rect 88670 343032 88675 343088
rect 60641 343030 88675 343032
rect 60641 343027 60707 343030
rect 88609 343027 88675 343030
rect 60549 342954 60615 342957
rect 90265 342954 90331 342957
rect 60549 342952 90331 342954
rect 60549 342896 60554 342952
rect 60610 342896 90270 342952
rect 90326 342896 90331 342952
rect 60549 342894 90331 342896
rect 60549 342891 60615 342894
rect 90265 342891 90331 342894
rect 64781 342818 64847 342821
rect 73705 342818 73771 342821
rect 64781 342816 73771 342818
rect 64781 342760 64786 342816
rect 64842 342760 73710 342816
rect 73766 342760 73771 342816
rect 64781 342758 73771 342760
rect 64781 342755 64847 342758
rect 73705 342755 73771 342758
rect 63125 342682 63191 342685
rect 77293 342682 77359 342685
rect 63125 342680 77359 342682
rect 63125 342624 63130 342680
rect 63186 342624 77298 342680
rect 77354 342624 77359 342680
rect 63125 342622 77359 342624
rect 63125 342619 63191 342622
rect 77293 342619 77359 342622
rect 211797 342682 211863 342685
rect 211797 342680 240212 342682
rect 211797 342624 211802 342680
rect 211858 342624 240212 342680
rect 211797 342622 240212 342624
rect 211797 342619 211863 342622
rect 67449 342140 67515 342141
rect 67398 342138 67404 342140
rect 67358 342078 67404 342138
rect 67468 342136 67515 342140
rect 67510 342080 67515 342136
rect 67398 342076 67404 342078
rect 67468 342076 67515 342080
rect 69790 342076 69796 342140
rect 69860 342138 69866 342140
rect 70301 342138 70367 342141
rect 69860 342136 70367 342138
rect 69860 342080 70306 342136
rect 70362 342080 70367 342136
rect 69860 342078 70367 342080
rect 69860 342076 69866 342078
rect 67449 342075 67515 342076
rect 70301 342075 70367 342078
rect 237557 342138 237623 342141
rect 237557 342136 240212 342138
rect 237557 342080 237562 342136
rect 237618 342080 240212 342136
rect 237557 342078 240212 342080
rect 237557 342075 237623 342078
rect 69422 341940 69428 342004
rect 69492 342002 69498 342004
rect 70209 342002 70275 342005
rect 230933 342002 230999 342005
rect 69492 342000 70275 342002
rect 69492 341944 70214 342000
rect 70270 341944 70275 342000
rect 69492 341942 70275 341944
rect 69492 341940 69498 341942
rect 70209 341939 70275 341942
rect 70350 342000 230999 342002
rect 70350 341944 230938 342000
rect 230994 341944 230999 342000
rect 70350 341942 230999 341944
rect 66110 341804 66116 341868
rect 66180 341866 66186 341868
rect 70350 341866 70410 341942
rect 230933 341939 230999 341942
rect 66180 341806 70410 341866
rect 70485 341866 70551 341869
rect 231301 341866 231367 341869
rect 285121 341866 285187 341869
rect 70485 341864 231367 341866
rect 70485 341808 70490 341864
rect 70546 341808 231306 341864
rect 231362 341808 231367 341864
rect 70485 341806 231367 341808
rect 279956 341864 285187 341866
rect 279956 341808 285126 341864
rect 285182 341808 285187 341864
rect 279956 341806 285187 341808
rect 66180 341804 66186 341806
rect 70485 341803 70551 341806
rect 231301 341803 231367 341806
rect 285121 341803 285187 341806
rect 66846 341668 66852 341732
rect 66916 341730 66922 341732
rect 234654 341730 234660 341732
rect 66916 341670 234660 341730
rect 66916 341668 66922 341670
rect 234654 341668 234660 341670
rect 234724 341668 234730 341732
rect 65742 341532 65748 341596
rect 65812 341594 65818 341596
rect 235022 341594 235028 341596
rect 65812 341534 235028 341594
rect 65812 341532 65818 341534
rect 235022 341532 235028 341534
rect 235092 341532 235098 341596
rect 237373 341594 237439 341597
rect 237373 341592 240212 341594
rect 237373 341536 237378 341592
rect 237434 341536 240212 341592
rect 237373 341534 240212 341536
rect 237373 341531 237439 341534
rect 65926 341396 65932 341460
rect 65996 341458 66002 341460
rect 70485 341458 70551 341461
rect 65996 341456 70551 341458
rect 65996 341400 70490 341456
rect 70546 341400 70551 341456
rect 65996 341398 70551 341400
rect 65996 341396 66002 341398
rect 70485 341395 70551 341398
rect 70669 341458 70735 341461
rect 235574 341458 235580 341460
rect 70669 341456 235580 341458
rect 70669 341400 70674 341456
rect 70730 341400 235580 341456
rect 70669 341398 235580 341400
rect 70669 341395 70735 341398
rect 235574 341396 235580 341398
rect 235644 341396 235650 341460
rect 67030 341260 67036 341324
rect 67100 341322 67106 341324
rect 231117 341322 231183 341325
rect 67100 341320 231183 341322
rect 67100 341264 231122 341320
rect 231178 341264 231183 341320
rect 67100 341262 231183 341264
rect 67100 341260 67106 341262
rect 231117 341259 231183 341262
rect 67214 341124 67220 341188
rect 67284 341186 67290 341188
rect 231485 341186 231551 341189
rect 67284 341184 231551 341186
rect 67284 341128 231490 341184
rect 231546 341128 231551 341184
rect 67284 341126 231551 341128
rect 67284 341124 67290 341126
rect 231485 341123 231551 341126
rect 65558 340988 65564 341052
rect 65628 341050 65634 341052
rect 70669 341050 70735 341053
rect 65628 341048 70735 341050
rect 65628 340992 70674 341048
rect 70730 340992 70735 341048
rect 65628 340990 70735 340992
rect 65628 340988 65634 340990
rect 70669 340987 70735 340990
rect 235206 340988 235212 341052
rect 235276 341050 235282 341052
rect 235809 341050 235875 341053
rect 235276 341048 235875 341050
rect 235276 340992 235814 341048
rect 235870 340992 235875 341048
rect 235276 340990 235875 340992
rect 235276 340988 235282 340990
rect 235809 340987 235875 340990
rect 237373 341050 237439 341053
rect 237373 341048 240212 341050
rect 237373 340992 237378 341048
rect 237434 340992 240212 341048
rect 237373 340990 240212 340992
rect 237373 340987 237439 340990
rect 235758 340852 235764 340916
rect 235828 340914 235834 340916
rect 235901 340914 235967 340917
rect 235828 340912 235967 340914
rect 235828 340856 235906 340912
rect 235962 340856 235967 340912
rect 235828 340854 235967 340856
rect 235828 340852 235834 340854
rect 235901 340851 235967 340854
rect 68921 340778 68987 340781
rect 229737 340778 229803 340781
rect 68921 340776 229803 340778
rect 68921 340720 68926 340776
rect 68982 340720 229742 340776
rect 229798 340720 229803 340776
rect 68921 340718 229803 340720
rect 68921 340715 68987 340718
rect 229737 340715 229803 340718
rect 195237 340506 195303 340509
rect 284937 340506 285003 340509
rect 195237 340504 240212 340506
rect 195237 340448 195242 340504
rect 195298 340448 240212 340504
rect 195237 340446 240212 340448
rect 279956 340504 285003 340506
rect 279956 340448 284942 340504
rect 284998 340448 285003 340504
rect 279956 340446 285003 340448
rect 195237 340443 195303 340446
rect 284937 340443 285003 340446
rect 69565 340234 69631 340237
rect 237833 340234 237899 340237
rect 69565 340232 237899 340234
rect 69565 340176 69570 340232
rect 69626 340176 237838 340232
rect 237894 340176 237899 340232
rect 69565 340174 237899 340176
rect 69565 340171 69631 340174
rect 237833 340171 237899 340174
rect 48221 340098 48287 340101
rect 68921 340098 68987 340101
rect 48221 340096 68987 340098
rect 48221 340040 48226 340096
rect 48282 340040 68926 340096
rect 68982 340040 68987 340096
rect 48221 340038 68987 340040
rect 48221 340035 48287 340038
rect 68921 340035 68987 340038
rect 70117 340098 70183 340101
rect 238017 340098 238083 340101
rect 70117 340096 238083 340098
rect 70117 340040 70122 340096
rect 70178 340040 238022 340096
rect 238078 340040 238083 340096
rect 70117 340038 238083 340040
rect 70117 340035 70183 340038
rect 238017 340035 238083 340038
rect 220077 339962 220143 339965
rect 220077 339960 240212 339962
rect 220077 339904 220082 339960
rect 220138 339904 240212 339960
rect 220077 339902 240212 339904
rect 220077 339899 220143 339902
rect 111742 339356 111748 339420
rect 111812 339418 111818 339420
rect 112989 339418 113055 339421
rect 111812 339416 113055 339418
rect 111812 339360 112994 339416
rect 113050 339360 113055 339416
rect 111812 339358 113055 339360
rect 111812 339356 111818 339358
rect 112989 339355 113055 339358
rect 142797 339418 142863 339421
rect 142797 339416 240212 339418
rect 142797 339360 142802 339416
rect 142858 339360 240212 339416
rect 142797 339358 240212 339360
rect 142797 339355 142863 339358
rect 280838 339146 280844 339148
rect 279956 339086 280844 339146
rect 280838 339084 280844 339086
rect 280908 339084 280914 339148
rect 175917 338874 175983 338877
rect 175917 338872 240212 338874
rect 175917 338816 175922 338872
rect 175978 338816 240212 338872
rect 175917 338814 240212 338816
rect 175917 338811 175983 338814
rect 112846 338602 112852 338604
rect 109940 338542 112852 338602
rect 112846 338540 112852 338542
rect 112916 338540 112922 338604
rect 583520 338452 584960 338692
rect 203517 338330 203583 338333
rect 203517 338328 240212 338330
rect 203517 338272 203522 338328
rect 203578 338272 240212 338328
rect 203517 338270 240212 338272
rect 203517 338267 203583 338270
rect 178677 337786 178743 337789
rect 283649 337786 283715 337789
rect 178677 337784 240212 337786
rect 178677 337728 178682 337784
rect 178738 337728 240212 337784
rect 178677 337726 240212 337728
rect 279956 337784 283715 337786
rect 279956 337728 283654 337784
rect 283710 337728 283715 337784
rect 279956 337726 283715 337728
rect 178677 337723 178743 337726
rect 283649 337723 283715 337726
rect 188337 337242 188403 337245
rect 188337 337240 240212 337242
rect 188337 337184 188342 337240
rect 188398 337184 240212 337240
rect 188337 337182 240212 337184
rect 188337 337179 188403 337182
rect 178534 336970 178540 336972
rect 109940 336910 178540 336970
rect 178534 336908 178540 336910
rect 178604 336908 178610 336972
rect 151077 336698 151143 336701
rect 151077 336696 240212 336698
rect 151077 336640 151082 336696
rect 151138 336640 240212 336696
rect 151077 336638 240212 336640
rect 151077 336635 151143 336638
rect 283741 336426 283807 336429
rect 279956 336424 283807 336426
rect 279956 336368 283746 336424
rect 283802 336368 283807 336424
rect 279956 336366 283807 336368
rect 283741 336363 283807 336366
rect 206277 336154 206343 336157
rect 206277 336152 240212 336154
rect 206277 336096 206282 336152
rect 206338 336096 240212 336152
rect 206277 336094 240212 336096
rect 206277 336091 206343 336094
rect 184197 335610 184263 335613
rect 184197 335608 240212 335610
rect 184197 335552 184202 335608
rect 184258 335552 240212 335608
rect 184197 335550 240212 335552
rect 184197 335547 184263 335550
rect 230054 335338 230060 335340
rect 109940 335278 230060 335338
rect 230054 335276 230060 335278
rect 230124 335276 230130 335340
rect 191097 335066 191163 335069
rect 291193 335066 291259 335069
rect 191097 335064 240212 335066
rect 191097 335008 191102 335064
rect 191158 335008 240212 335064
rect 191097 335006 240212 335008
rect 279956 335064 291259 335066
rect 279956 335008 291198 335064
rect 291254 335008 291259 335064
rect 279956 335006 291259 335008
rect 191097 335003 191163 335006
rect 291193 335003 291259 335006
rect 197997 334522 198063 334525
rect 197997 334520 240212 334522
rect 197997 334464 198002 334520
rect 198058 334464 240212 334520
rect 197997 334462 240212 334464
rect 197997 334459 198063 334462
rect 230289 334116 230355 334117
rect 230238 334114 230244 334116
rect 230198 334054 230244 334114
rect 230308 334112 230355 334116
rect 230350 334056 230355 334112
rect 230238 334052 230244 334054
rect 230308 334052 230355 334056
rect 230289 334051 230355 334052
rect 186957 333978 187023 333981
rect 186957 333976 240212 333978
rect 186957 333920 186962 333976
rect 187018 333920 240212 333976
rect 186957 333918 240212 333920
rect 186957 333915 187023 333918
rect 219934 333706 219940 333708
rect 109940 333646 219940 333706
rect 219934 333644 219940 333646
rect 220004 333644 220010 333708
rect 286133 333706 286199 333709
rect 279956 333704 286199 333706
rect 279956 333648 286138 333704
rect 286194 333648 286199 333704
rect 279956 333646 286199 333648
rect 286133 333643 286199 333646
rect 225689 333434 225755 333437
rect 225689 333432 240212 333434
rect 225689 333376 225694 333432
rect 225750 333376 240212 333432
rect 225689 333374 240212 333376
rect 225689 333371 225755 333374
rect 209037 332890 209103 332893
rect 209037 332888 240212 332890
rect 209037 332832 209042 332888
rect 209098 332832 240212 332888
rect 209037 332830 240212 332832
rect 209037 332827 209103 332830
rect -960 332196 480 332436
rect 224309 332346 224375 332349
rect 288433 332346 288499 332349
rect 224309 332344 240212 332346
rect 224309 332288 224314 332344
rect 224370 332288 240212 332344
rect 224309 332286 240212 332288
rect 279956 332344 288499 332346
rect 279956 332288 288438 332344
rect 288494 332288 288499 332344
rect 279956 332286 288499 332288
rect 224309 332283 224375 332286
rect 288433 332283 288499 332286
rect 228398 332074 228404 332076
rect 109940 332014 228404 332074
rect 228398 332012 228404 332014
rect 228468 332012 228474 332076
rect 229829 331802 229895 331805
rect 229829 331800 240212 331802
rect 229829 331744 229834 331800
rect 229890 331744 240212 331800
rect 229829 331742 240212 331744
rect 229829 331739 229895 331742
rect 228030 331332 228036 331396
rect 228100 331394 228106 331396
rect 228725 331394 228791 331397
rect 228100 331392 228791 331394
rect 228100 331336 228730 331392
rect 228786 331336 228791 331392
rect 228100 331334 228791 331336
rect 228100 331332 228106 331334
rect 228725 331331 228791 331334
rect 119337 331258 119403 331261
rect 119337 331256 240212 331258
rect 119337 331200 119342 331256
rect 119398 331200 240212 331256
rect 119337 331198 240212 331200
rect 119337 331195 119403 331198
rect 286501 330986 286567 330989
rect 279956 330984 286567 330986
rect 279956 330928 286506 330984
rect 286562 330928 286567 330984
rect 279956 330926 286567 330928
rect 286501 330923 286567 330926
rect 226977 330714 227043 330717
rect 226977 330712 240212 330714
rect 226977 330656 226982 330712
rect 227038 330656 240212 330712
rect 226977 330654 240212 330656
rect 226977 330651 227043 330654
rect 227110 330442 227116 330444
rect 109940 330382 227116 330442
rect 227110 330380 227116 330382
rect 227180 330380 227186 330444
rect 214557 330170 214623 330173
rect 214557 330168 240212 330170
rect 214557 330112 214562 330168
rect 214618 330112 240212 330168
rect 214557 330110 240212 330112
rect 214557 330107 214623 330110
rect 229737 329762 229803 329765
rect 229737 329760 240242 329762
rect 229737 329704 229742 329760
rect 229798 329704 240242 329760
rect 229737 329702 240242 329704
rect 229737 329699 229803 329702
rect 240182 329596 240242 329702
rect 285857 329626 285923 329629
rect 279956 329624 285923 329626
rect 279956 329568 285862 329624
rect 285918 329568 285923 329624
rect 279956 329566 285923 329568
rect 285857 329563 285923 329566
rect 231669 329082 231735 329085
rect 231669 329080 240212 329082
rect 231669 329024 231674 329080
rect 231730 329024 240212 329080
rect 231669 329022 240212 329024
rect 231669 329019 231735 329022
rect 299974 329020 299980 329084
rect 300044 329082 300050 329084
rect 580206 329082 580212 329084
rect 300044 329022 580212 329082
rect 300044 329020 300050 329022
rect 580206 329020 580212 329022
rect 580276 329020 580282 329084
rect 224166 328810 224172 328812
rect 109940 328750 224172 328810
rect 224166 328748 224172 328750
rect 224236 328748 224242 328812
rect 225965 328538 226031 328541
rect 225965 328536 240212 328538
rect 225965 328480 225970 328536
rect 226026 328480 240212 328536
rect 225965 328478 240212 328480
rect 225965 328475 226031 328478
rect 286409 328266 286475 328269
rect 279956 328264 286475 328266
rect 279956 328208 286414 328264
rect 286470 328208 286475 328264
rect 279956 328206 286475 328208
rect 286409 328203 286475 328206
rect 222101 327994 222167 327997
rect 222101 327992 240212 327994
rect 222101 327936 222106 327992
rect 222162 327936 240212 327992
rect 222101 327934 240212 327936
rect 222101 327931 222167 327934
rect 224861 327450 224927 327453
rect 224861 327448 240212 327450
rect 224861 327392 224866 327448
rect 224922 327392 240212 327448
rect 224861 327390 240212 327392
rect 224861 327387 224927 327390
rect 222694 327178 222700 327180
rect 109940 327118 222700 327178
rect 222694 327116 222700 327118
rect 222764 327116 222770 327180
rect 232957 326906 233023 326909
rect 286225 326906 286291 326909
rect 232957 326904 240212 326906
rect 232957 326848 232962 326904
rect 233018 326848 240212 326904
rect 232957 326846 240212 326848
rect 279956 326904 286291 326906
rect 279956 326848 286230 326904
rect 286286 326848 286291 326904
rect 279956 326846 286291 326848
rect 232957 326843 233023 326846
rect 286225 326843 286291 326846
rect 239438 326300 239444 326364
rect 239508 326362 239514 326364
rect 239508 326302 240212 326362
rect 239508 326300 239514 326302
rect 237925 325818 237991 325821
rect 237925 325816 240212 325818
rect 237925 325760 237930 325816
rect 237986 325760 240212 325816
rect 237925 325758 240212 325760
rect 237925 325755 237991 325758
rect 231526 325546 231532 325548
rect 109940 325486 231532 325546
rect 231526 325484 231532 325486
rect 231596 325484 231602 325548
rect 286317 325546 286383 325549
rect 279956 325544 286383 325546
rect 279956 325488 286322 325544
rect 286378 325488 286383 325544
rect 279956 325486 286383 325488
rect 286317 325483 286383 325486
rect 226057 325274 226123 325277
rect 226057 325272 240212 325274
rect 226057 325216 226062 325272
rect 226118 325216 240212 325272
rect 226057 325214 240212 325216
rect 226057 325211 226123 325214
rect 580206 325212 580212 325276
rect 580276 325274 580282 325276
rect 583520 325274 584960 325364
rect 580276 325214 584960 325274
rect 580276 325212 580282 325214
rect 583520 325124 584960 325214
rect 48129 325002 48195 325005
rect 48129 325000 50140 325002
rect 48129 324944 48134 325000
rect 48190 324944 50140 325000
rect 48129 324942 50140 324944
rect 48129 324939 48195 324942
rect 235809 324730 235875 324733
rect 235809 324728 240212 324730
rect 235809 324672 235814 324728
rect 235870 324672 240212 324728
rect 235809 324670 240212 324672
rect 235809 324667 235875 324670
rect 230606 324396 230612 324460
rect 230676 324458 230682 324460
rect 231393 324458 231459 324461
rect 230676 324456 231459 324458
rect 230676 324400 231398 324456
rect 231454 324400 231459 324456
rect 230676 324398 231459 324400
rect 230676 324396 230682 324398
rect 231393 324395 231459 324398
rect 238109 324186 238175 324189
rect 285949 324186 286015 324189
rect 238109 324184 240212 324186
rect 238109 324128 238114 324184
rect 238170 324128 240212 324184
rect 238109 324126 240212 324128
rect 279956 324184 286015 324186
rect 279956 324128 285954 324184
rect 286010 324128 286015 324184
rect 279956 324126 286015 324128
rect 238109 324123 238175 324126
rect 285949 324123 286015 324126
rect 112662 323914 112668 323916
rect 109940 323854 112668 323914
rect 112662 323852 112668 323854
rect 112732 323852 112738 323916
rect 238293 323642 238359 323645
rect 238293 323640 240212 323642
rect 238293 323584 238298 323640
rect 238354 323584 240212 323640
rect 238293 323582 240212 323584
rect 238293 323579 238359 323582
rect 239806 323036 239812 323100
rect 239876 323098 239882 323100
rect 239876 323038 240212 323098
rect 239876 323036 239882 323038
rect 111926 322900 111932 322964
rect 111996 322962 112002 322964
rect 113081 322962 113147 322965
rect 111996 322960 113147 322962
rect 111996 322904 113086 322960
rect 113142 322904 113147 322960
rect 111996 322902 113147 322904
rect 111996 322900 112002 322902
rect 113081 322899 113147 322902
rect 286041 322826 286107 322829
rect 279956 322824 286107 322826
rect 279956 322768 286046 322824
rect 286102 322768 286107 322824
rect 279956 322766 286107 322768
rect 286041 322763 286107 322766
rect 234245 322554 234311 322557
rect 234245 322552 240212 322554
rect 234245 322496 234250 322552
rect 234306 322496 240212 322552
rect 234245 322494 240212 322496
rect 234245 322491 234311 322494
rect 226926 322282 226932 322284
rect 109940 322222 226932 322282
rect 226926 322220 226932 322222
rect 226996 322220 227002 322284
rect 238201 322010 238267 322013
rect 238201 322008 240212 322010
rect 238201 321952 238206 322008
rect 238262 321952 240212 322008
rect 238201 321950 240212 321952
rect 238201 321947 238267 321950
rect 234337 321466 234403 321469
rect 285673 321466 285739 321469
rect 234337 321464 240212 321466
rect 234337 321408 234342 321464
rect 234398 321408 240212 321464
rect 234337 321406 240212 321408
rect 279956 321464 285739 321466
rect 279956 321408 285678 321464
rect 285734 321408 285739 321464
rect 279956 321406 285739 321408
rect 234337 321403 234403 321406
rect 285673 321403 285739 321406
rect 231761 320922 231827 320925
rect 237373 320922 237439 320925
rect 231761 320920 237439 320922
rect 231761 320864 231766 320920
rect 231822 320864 237378 320920
rect 237434 320864 237439 320920
rect 231761 320862 237439 320864
rect 231761 320859 231827 320862
rect 237373 320859 237439 320862
rect 238569 320922 238635 320925
rect 238569 320920 240212 320922
rect 238569 320864 238574 320920
rect 238630 320864 240212 320920
rect 238569 320862 240212 320864
rect 238569 320859 238635 320862
rect 112478 320650 112484 320652
rect 109940 320590 112484 320650
rect 112478 320588 112484 320590
rect 112548 320588 112554 320652
rect 234521 320378 234587 320381
rect 234521 320376 240212 320378
rect 234521 320320 234526 320376
rect 234582 320320 240212 320376
rect 234521 320318 240212 320320
rect 234521 320315 234587 320318
rect 285765 320106 285831 320109
rect 279956 320104 285831 320106
rect 279956 320048 285770 320104
rect 285826 320048 285831 320104
rect 279956 320046 285831 320048
rect 285765 320043 285831 320046
rect 238385 319834 238451 319837
rect 238385 319832 240212 319834
rect 238385 319776 238390 319832
rect 238446 319776 240212 319832
rect 238385 319774 240212 319776
rect 238385 319771 238451 319774
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 226241 319290 226307 319293
rect 226241 319288 240212 319290
rect 226241 319232 226246 319288
rect 226302 319232 240212 319288
rect 226241 319230 240212 319232
rect 226241 319227 226307 319230
rect 230974 319018 230980 319020
rect 109940 318958 230980 319018
rect 230974 318956 230980 318958
rect 231044 318956 231050 319020
rect 238661 318746 238727 318749
rect 285622 318746 285628 318748
rect 238661 318744 240212 318746
rect 238661 318688 238666 318744
rect 238722 318688 240212 318744
rect 238661 318686 240212 318688
rect 279956 318686 285628 318746
rect 238661 318683 238727 318686
rect 285622 318684 285628 318686
rect 285692 318684 285698 318748
rect 224350 318140 224356 318204
rect 224420 318202 224426 318204
rect 224420 318142 240212 318202
rect 224420 318140 224426 318142
rect 116393 318066 116459 318069
rect 227161 318066 227227 318069
rect 116393 318064 227227 318066
rect 116393 318008 116398 318064
rect 116454 318008 227166 318064
rect 227222 318008 227227 318064
rect 116393 318006 227227 318008
rect 116393 318003 116459 318006
rect 227161 318003 227227 318006
rect 238477 317658 238543 317661
rect 238477 317656 240212 317658
rect 238477 317600 238482 317656
rect 238538 317600 240212 317656
rect 238477 317598 240212 317600
rect 238477 317595 238543 317598
rect 229870 317386 229876 317388
rect 109940 317326 229876 317386
rect 229870 317324 229876 317326
rect 229940 317324 229946 317388
rect 284334 317386 284340 317388
rect 279956 317326 284340 317386
rect 284334 317324 284340 317326
rect 284404 317324 284410 317388
rect 238334 317052 238340 317116
rect 238404 317114 238410 317116
rect 238404 317054 240212 317114
rect 238404 317052 238410 317054
rect 237373 316978 237439 316981
rect 238334 316978 238340 316980
rect 237373 316976 238340 316978
rect 237373 316920 237378 316976
rect 237434 316920 238340 316976
rect 237373 316918 238340 316920
rect 237373 316915 237439 316918
rect 238334 316916 238340 316918
rect 238404 316916 238410 316980
rect 224534 316508 224540 316572
rect 224604 316570 224610 316572
rect 224604 316510 240212 316570
rect 224604 316508 224610 316510
rect 238150 315964 238156 316028
rect 238220 316026 238226 316028
rect 282913 316026 282979 316029
rect 238220 315966 240212 316026
rect 279956 316024 282979 316026
rect 279956 315968 282918 316024
rect 282974 315968 282979 316024
rect 279956 315966 282979 315968
rect 238220 315964 238226 315966
rect 282913 315963 282979 315966
rect 228214 315754 228220 315756
rect 109940 315694 228220 315754
rect 228214 315692 228220 315694
rect 228284 315692 228290 315756
rect 224718 315420 224724 315484
rect 224788 315482 224794 315484
rect 224788 315422 240212 315482
rect 224788 315420 224794 315422
rect 234061 314938 234127 314941
rect 234061 314936 240212 314938
rect 234061 314880 234066 314936
rect 234122 314880 240212 314936
rect 234061 314878 240212 314880
rect 234061 314875 234127 314878
rect 280654 314666 280660 314668
rect 279956 314606 280660 314666
rect 280654 314604 280660 314606
rect 280724 314604 280730 314668
rect 235901 314394 235967 314397
rect 235901 314392 240212 314394
rect 235901 314336 235906 314392
rect 235962 314336 240212 314392
rect 235901 314334 240212 314336
rect 235901 314331 235967 314334
rect 231894 314122 231900 314124
rect 109940 314062 231900 314122
rect 231894 314060 231900 314062
rect 231964 314060 231970 314124
rect 233877 313850 233943 313853
rect 233877 313848 240212 313850
rect 233877 313792 233882 313848
rect 233938 313792 240212 313848
rect 233877 313790 240212 313792
rect 233877 313787 233943 313790
rect 232078 313244 232084 313308
rect 232148 313306 232154 313308
rect 233049 313306 233115 313309
rect 232148 313304 233115 313306
rect 232148 313248 233054 313304
rect 233110 313248 233115 313304
rect 232148 313246 233115 313248
rect 232148 313244 232154 313246
rect 233049 313243 233115 313246
rect 234429 313306 234495 313309
rect 282269 313306 282335 313309
rect 234429 313304 240212 313306
rect 234429 313248 234434 313304
rect 234490 313248 240212 313304
rect 234429 313246 240212 313248
rect 279956 313304 282335 313306
rect 279956 313248 282274 313304
rect 282330 313248 282335 313304
rect 279956 313246 282335 313248
rect 234429 313243 234495 313246
rect 282269 313243 282335 313246
rect 233969 312762 234035 312765
rect 233969 312760 240212 312762
rect 233969 312704 233974 312760
rect 234030 312704 240212 312760
rect 233969 312702 240212 312704
rect 233969 312699 234035 312702
rect 111742 312490 111748 312492
rect 109940 312430 111748 312490
rect 111742 312428 111748 312430
rect 111812 312428 111818 312492
rect 234153 312218 234219 312221
rect 234153 312216 240212 312218
rect 234153 312160 234158 312216
rect 234214 312160 240212 312216
rect 234153 312158 240212 312160
rect 234153 312155 234219 312158
rect 281441 312082 281507 312085
rect 279926 312080 281507 312082
rect 279926 312024 281446 312080
rect 281502 312024 281507 312080
rect 279926 312022 281507 312024
rect 279926 311916 279986 312022
rect 281441 312019 281507 312022
rect 544326 312020 544332 312084
rect 544396 312082 544402 312084
rect 583520 312082 584960 312172
rect 544396 312022 584960 312082
rect 544396 312020 544402 312022
rect 280797 311946 280863 311949
rect 281533 311946 281599 311949
rect 280797 311944 281599 311946
rect 280797 311888 280802 311944
rect 280858 311888 281538 311944
rect 281594 311888 281599 311944
rect 583520 311932 584960 312022
rect 280797 311886 281599 311888
rect 280797 311883 280863 311886
rect 281533 311883 281599 311886
rect 234102 311612 234108 311676
rect 234172 311674 234178 311676
rect 234172 311614 240212 311674
rect 234172 311612 234178 311614
rect 234286 311068 234292 311132
rect 234356 311130 234362 311132
rect 234356 311070 240212 311130
rect 234356 311068 234362 311070
rect 230422 310858 230428 310860
rect 109940 310798 230428 310858
rect 230422 310796 230428 310798
rect 230492 310796 230498 310860
rect 234470 310524 234476 310588
rect 234540 310586 234546 310588
rect 282361 310586 282427 310589
rect 234540 310526 240212 310586
rect 279956 310584 282427 310586
rect 279956 310528 282366 310584
rect 282422 310528 282427 310584
rect 279956 310526 282427 310528
rect 234540 310524 234546 310526
rect 282361 310523 282427 310526
rect 238518 309980 238524 310044
rect 238588 310042 238594 310044
rect 238588 309982 240212 310042
rect 238588 309980 238594 309982
rect 233918 309436 233924 309500
rect 233988 309498 233994 309500
rect 233988 309438 240212 309498
rect 233988 309436 233994 309438
rect 112294 309226 112300 309228
rect 109940 309166 112300 309226
rect 112294 309164 112300 309166
rect 112364 309164 112370 309228
rect 282177 309226 282243 309229
rect 279956 309224 282243 309226
rect 279956 309168 282182 309224
rect 282238 309168 282243 309224
rect 279956 309166 282243 309168
rect 282177 309163 282243 309166
rect 222694 308892 222700 308956
rect 222764 308954 222770 308956
rect 222764 308894 240212 308954
rect 222764 308892 222770 308894
rect 224166 308348 224172 308412
rect 224236 308410 224242 308412
rect 224236 308350 240212 308410
rect 224236 308348 224242 308350
rect 230974 307804 230980 307868
rect 231044 307866 231050 307868
rect 284518 307866 284524 307868
rect 231044 307806 240212 307866
rect 279956 307806 284524 307866
rect 231044 307804 231050 307806
rect 284518 307804 284524 307806
rect 284588 307804 284594 307868
rect 234654 307668 234660 307732
rect 234724 307730 234730 307732
rect 235901 307730 235967 307733
rect 234724 307728 235967 307730
rect 234724 307672 235906 307728
rect 235962 307672 235967 307728
rect 234724 307670 235967 307672
rect 234724 307668 234730 307670
rect 235901 307667 235967 307670
rect 111926 307594 111932 307596
rect 109940 307534 111932 307594
rect 111926 307532 111932 307534
rect 111996 307532 112002 307596
rect 235206 307260 235212 307324
rect 235276 307322 235282 307324
rect 235276 307262 240212 307322
rect 235276 307260 235282 307262
rect 228214 306716 228220 306780
rect 228284 306778 228290 306780
rect 228284 306718 240212 306778
rect 228284 306716 228290 306718
rect 282545 306506 282611 306509
rect 279956 306504 282611 306506
rect 279956 306448 282550 306504
rect 282606 306448 282611 306504
rect 279956 306446 282611 306448
rect 282545 306443 282611 306446
rect -960 306234 480 306324
rect 48630 306234 48636 306236
rect -960 306174 48636 306234
rect -960 306084 480 306174
rect 48630 306172 48636 306174
rect 48700 306172 48706 306236
rect 231342 306172 231348 306236
rect 231412 306234 231418 306236
rect 231412 306174 240212 306234
rect 231412 306172 231418 306174
rect 218697 305962 218763 305965
rect 109940 305960 218763 305962
rect 109940 305904 218702 305960
rect 218758 305904 218763 305960
rect 109940 305902 218763 305904
rect 218697 305899 218763 305902
rect 122046 305628 122052 305692
rect 122116 305690 122122 305692
rect 122116 305630 240212 305690
rect 122116 305628 122122 305630
rect 147070 305084 147076 305148
rect 147140 305146 147146 305148
rect 281809 305146 281875 305149
rect 147140 305086 240212 305146
rect 279956 305144 281875 305146
rect 279956 305088 281814 305144
rect 281870 305088 281875 305144
rect 279956 305086 281875 305088
rect 147140 305084 147146 305086
rect 281809 305083 281875 305086
rect 173198 304540 173204 304604
rect 173268 304602 173274 304604
rect 173268 304542 240212 304602
rect 173268 304540 173274 304542
rect 218830 304330 218836 304332
rect 109940 304270 218836 304330
rect 218830 304268 218836 304270
rect 218900 304268 218906 304332
rect 228909 304058 228975 304061
rect 228909 304056 240212 304058
rect 228909 304000 228914 304056
rect 228970 304000 240212 304056
rect 228909 303998 240212 304000
rect 228909 303995 228975 303998
rect 279366 303724 279372 303788
rect 279436 303724 279442 303788
rect 130326 303452 130332 303516
rect 130396 303514 130402 303516
rect 130396 303454 240212 303514
rect 130396 303452 130402 303454
rect 161974 302908 161980 302972
rect 162044 302970 162050 302972
rect 162044 302910 240212 302970
rect 162044 302908 162050 302910
rect 218646 302698 218652 302700
rect 109940 302638 218652 302698
rect 218646 302636 218652 302638
rect 218716 302636 218722 302700
rect 210366 302364 210372 302428
rect 210436 302426 210442 302428
rect 281758 302426 281764 302428
rect 210436 302366 240212 302426
rect 279956 302366 281764 302426
rect 210436 302364 210442 302366
rect 281758 302364 281764 302366
rect 281828 302364 281834 302428
rect 151169 301882 151235 301885
rect 151169 301880 240212 301882
rect 151169 301824 151174 301880
rect 151230 301824 240212 301880
rect 151169 301822 240212 301824
rect 151169 301819 151235 301822
rect 231209 301338 231275 301341
rect 231209 301336 240212 301338
rect 231209 301280 231214 301336
rect 231270 301280 240212 301336
rect 231209 301278 240212 301280
rect 231209 301275 231275 301278
rect 221038 301066 221044 301068
rect 109940 301006 221044 301066
rect 221038 301004 221044 301006
rect 221108 301004 221114 301068
rect 284702 301066 284708 301068
rect 279956 301006 284708 301066
rect 284702 301004 284708 301006
rect 284772 301004 284778 301068
rect 237373 300794 237439 300797
rect 237373 300792 240212 300794
rect 237373 300736 237378 300792
rect 237434 300736 240212 300792
rect 237373 300734 240212 300736
rect 237373 300731 237439 300734
rect 239765 300250 239831 300253
rect 239765 300248 240212 300250
rect 239765 300192 239770 300248
rect 239826 300192 240212 300248
rect 239765 300190 240212 300192
rect 239765 300187 239831 300190
rect 239857 299706 239923 299709
rect 282126 299706 282132 299708
rect 239857 299704 240212 299706
rect 239857 299648 239862 299704
rect 239918 299648 240212 299704
rect 239857 299646 240212 299648
rect 279956 299646 282132 299706
rect 239857 299643 239923 299646
rect 282126 299644 282132 299646
rect 282196 299644 282202 299708
rect 222009 299434 222075 299437
rect 109940 299432 222075 299434
rect 109940 299376 222014 299432
rect 222070 299376 222075 299432
rect 109940 299374 222075 299376
rect 222009 299371 222075 299374
rect 280981 299434 281047 299437
rect 281625 299434 281691 299437
rect 280981 299432 281691 299434
rect 280981 299376 280986 299432
rect 281042 299376 281630 299432
rect 281686 299376 281691 299432
rect 280981 299374 281691 299376
rect 280981 299371 281047 299374
rect 281625 299371 281691 299374
rect 227621 299162 227687 299165
rect 227621 299160 240212 299162
rect 227621 299104 227626 299160
rect 227682 299104 240212 299160
rect 227621 299102 240212 299104
rect 227621 299099 227687 299102
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 237281 298618 237347 298621
rect 237281 298616 240212 298618
rect 237281 298560 237286 298616
rect 237342 298560 240212 298616
rect 583520 298604 584960 298694
rect 237281 298558 240212 298560
rect 237281 298555 237347 298558
rect 282085 298346 282151 298349
rect 279956 298344 282151 298346
rect 279956 298288 282090 298344
rect 282146 298288 282151 298344
rect 279956 298286 282151 298288
rect 282085 298283 282151 298286
rect 237230 298012 237236 298076
rect 237300 298074 237306 298076
rect 237300 298014 240212 298074
rect 237300 298012 237306 298014
rect 221222 297802 221228 297804
rect 109940 297742 221228 297802
rect 221222 297740 221228 297742
rect 221292 297740 221298 297804
rect 228173 297530 228239 297533
rect 228173 297528 240212 297530
rect 228173 297472 228178 297528
rect 228234 297472 240212 297528
rect 228173 297470 240212 297472
rect 228173 297467 228239 297470
rect 230381 296986 230447 296989
rect 280061 296986 280127 296989
rect 230381 296984 240212 296986
rect 230381 296928 230386 296984
rect 230442 296928 240212 296984
rect 230381 296926 240212 296928
rect 279956 296984 280127 296986
rect 279956 296928 280066 296984
rect 280122 296928 280127 296984
rect 279956 296926 280127 296928
rect 230381 296923 230447 296926
rect 280061 296923 280127 296926
rect 233141 296442 233207 296445
rect 233141 296440 240212 296442
rect 233141 296384 233146 296440
rect 233202 296384 240212 296440
rect 233141 296382 240212 296384
rect 233141 296379 233207 296382
rect 224902 296170 224908 296172
rect 109940 296110 224908 296170
rect 224902 296108 224908 296110
rect 224972 296108 224978 296172
rect 232078 295836 232084 295900
rect 232148 295898 232154 295900
rect 232148 295838 240212 295898
rect 232148 295836 232154 295838
rect 282821 295626 282887 295629
rect 279956 295624 282887 295626
rect 279956 295568 282826 295624
rect 282882 295568 282887 295624
rect 279956 295566 282887 295568
rect 282821 295563 282887 295566
rect 224902 295292 224908 295356
rect 224972 295354 224978 295356
rect 226149 295354 226215 295357
rect 224972 295352 226215 295354
rect 224972 295296 226154 295352
rect 226210 295296 226215 295352
rect 224972 295294 226215 295296
rect 224972 295292 224978 295294
rect 226149 295291 226215 295294
rect 238334 295292 238340 295356
rect 238404 295354 238410 295356
rect 238404 295294 240212 295354
rect 238404 295292 238410 295294
rect 48221 295082 48287 295085
rect 48221 295080 50140 295082
rect 48221 295024 48226 295080
rect 48282 295024 50140 295080
rect 48221 295022 50140 295024
rect 48221 295019 48287 295022
rect 230238 294748 230244 294812
rect 230308 294810 230314 294812
rect 230308 294750 240212 294810
rect 230308 294748 230314 294750
rect 228030 294538 228036 294540
rect 109940 294478 228036 294538
rect 228030 294476 228036 294478
rect 228100 294476 228106 294540
rect 232262 294204 232268 294268
rect 232332 294266 232338 294268
rect 284886 294266 284892 294268
rect 232332 294206 240212 294266
rect 279956 294206 284892 294266
rect 232332 294204 232338 294206
rect 284886 294204 284892 294206
rect 284956 294204 284962 294268
rect 239622 293660 239628 293724
rect 239692 293722 239698 293724
rect 239692 293662 240212 293722
rect 239692 293660 239698 293662
rect -960 293178 480 293268
rect 3366 293178 3372 293180
rect -960 293118 3372 293178
rect -960 293028 480 293118
rect 3366 293116 3372 293118
rect 3436 293116 3442 293180
rect 238150 293116 238156 293180
rect 238220 293178 238226 293180
rect 238220 293118 240212 293178
rect 238220 293116 238226 293118
rect 227846 292906 227852 292908
rect 109940 292846 227852 292906
rect 227846 292844 227852 292846
rect 227916 292844 227922 292908
rect 281574 292906 281580 292908
rect 279956 292846 281580 292906
rect 281574 292844 281580 292846
rect 281644 292844 281650 292908
rect 238518 292572 238524 292636
rect 238588 292634 238594 292636
rect 238588 292574 240212 292634
rect 238588 292572 238594 292574
rect 238334 292028 238340 292092
rect 238404 292090 238410 292092
rect 238404 292030 240212 292090
rect 238404 292028 238410 292030
rect 239254 291484 239260 291548
rect 239324 291546 239330 291548
rect 281022 291546 281028 291548
rect 239324 291486 240212 291546
rect 279956 291486 281028 291546
rect 239324 291484 239330 291486
rect 281022 291484 281028 291486
rect 281092 291484 281098 291548
rect 227662 291274 227668 291276
rect 109940 291214 227668 291274
rect 227662 291212 227668 291214
rect 227732 291212 227738 291276
rect 239438 290940 239444 291004
rect 239508 291002 239514 291004
rect 239508 290942 240212 291002
rect 239508 290940 239514 290942
rect 239622 290396 239628 290460
rect 239692 290458 239698 290460
rect 239692 290398 240212 290458
rect 239692 290396 239698 290398
rect 283046 290186 283052 290188
rect 279956 290126 283052 290186
rect 283046 290124 283052 290126
rect 283116 290124 283122 290188
rect 239806 289852 239812 289916
rect 239876 289914 239882 289916
rect 239876 289854 240212 289914
rect 239876 289852 239882 289854
rect 230606 289642 230612 289644
rect 109940 289582 230612 289642
rect 230606 289580 230612 289582
rect 230676 289580 230682 289644
rect 239857 289370 239923 289373
rect 239857 289368 240212 289370
rect 239857 289312 239862 289368
rect 239918 289312 240212 289368
rect 239857 289310 240212 289312
rect 239857 289307 239923 289310
rect 239765 288826 239831 288829
rect 287421 288826 287487 288829
rect 239765 288824 240212 288826
rect 239765 288768 239770 288824
rect 239826 288768 240212 288824
rect 239765 288766 240212 288768
rect 279956 288824 287487 288826
rect 279956 288768 287426 288824
rect 287482 288768 287487 288824
rect 279956 288766 287487 288768
rect 239765 288763 239831 288766
rect 287421 288763 287487 288766
rect 214649 288282 214715 288285
rect 214649 288280 240212 288282
rect 214649 288224 214654 288280
rect 214710 288224 240212 288280
rect 214649 288222 240212 288224
rect 214649 288219 214715 288222
rect 231158 288010 231164 288012
rect 109940 287950 231164 288010
rect 231158 287948 231164 287950
rect 231228 287948 231234 288012
rect 224217 287738 224283 287741
rect 224217 287736 240212 287738
rect 224217 287680 224222 287736
rect 224278 287680 240212 287736
rect 224217 287678 240212 287680
rect 224217 287675 224283 287678
rect 288382 287466 288388 287468
rect 279956 287406 288388 287466
rect 288382 287404 288388 287406
rect 288452 287404 288458 287468
rect 237373 287194 237439 287197
rect 237373 287192 240212 287194
rect 237373 287136 237378 287192
rect 237434 287136 240212 287192
rect 237373 287134 240212 287136
rect 237373 287131 237439 287134
rect 237833 286650 237899 286653
rect 237833 286648 240212 286650
rect 237833 286592 237838 286648
rect 237894 286592 240212 286648
rect 237833 286590 240212 286592
rect 237833 286587 237899 286590
rect 224902 286378 224908 286380
rect 109940 286318 224908 286378
rect 224902 286316 224908 286318
rect 224972 286316 224978 286380
rect 237373 286106 237439 286109
rect 283414 286106 283420 286108
rect 237373 286104 240212 286106
rect 237373 286048 237378 286104
rect 237434 286048 240212 286104
rect 237373 286046 240212 286048
rect 279956 286046 283420 286106
rect 237373 286043 237439 286046
rect 283414 286044 283420 286046
rect 283484 286044 283490 286108
rect 237373 285562 237439 285565
rect 237373 285560 240212 285562
rect 237373 285504 237378 285560
rect 237434 285504 240212 285560
rect 237373 285502 240212 285504
rect 237373 285499 237439 285502
rect 583520 285276 584960 285516
rect 123477 285018 123543 285021
rect 123477 285016 240212 285018
rect 123477 284960 123482 285016
rect 123538 284960 240212 285016
rect 123477 284958 240212 284960
rect 123477 284955 123543 284958
rect 226190 284746 226196 284748
rect 109940 284686 226196 284746
rect 226190 284684 226196 284686
rect 226260 284684 226266 284748
rect 283230 284746 283236 284748
rect 279956 284686 283236 284746
rect 283230 284684 283236 284686
rect 283300 284684 283306 284748
rect 238017 284474 238083 284477
rect 238017 284472 240212 284474
rect 238017 284416 238022 284472
rect 238078 284416 240212 284472
rect 238017 284414 240212 284416
rect 238017 284411 238083 284414
rect 225781 283930 225847 283933
rect 225781 283928 240212 283930
rect 225781 283872 225786 283928
rect 225842 283872 240212 283928
rect 225781 283870 240212 283872
rect 225781 283867 225847 283870
rect 225413 283386 225479 283389
rect 287830 283386 287836 283388
rect 225413 283384 240212 283386
rect 225413 283328 225418 283384
rect 225474 283328 240212 283384
rect 225413 283326 240212 283328
rect 279956 283326 287836 283386
rect 225413 283323 225479 283326
rect 287830 283324 287836 283326
rect 287900 283324 287906 283388
rect 237966 283114 237972 283116
rect 109940 283054 237972 283114
rect 237966 283052 237972 283054
rect 238036 283052 238042 283116
rect 237414 282916 237420 282980
rect 237484 282916 237490 282980
rect 287278 282916 287284 282980
rect 287348 282978 287354 282980
rect 287605 282978 287671 282981
rect 287348 282976 287671 282978
rect 287348 282920 287610 282976
rect 287666 282920 287671 282976
rect 287348 282918 287671 282920
rect 287348 282916 287354 282918
rect 237422 282842 237482 282916
rect 287605 282915 287671 282918
rect 237422 282782 240212 282842
rect 237373 282298 237439 282301
rect 237373 282296 240212 282298
rect 237373 282240 237378 282296
rect 237434 282240 240212 282296
rect 237373 282238 240212 282240
rect 237373 282235 237439 282238
rect 287278 282026 287284 282028
rect 279956 281966 287284 282026
rect 287278 281964 287284 281966
rect 287348 281964 287354 282028
rect 287094 281828 287100 281892
rect 287164 281890 287170 281892
rect 287513 281890 287579 281893
rect 287164 281888 287579 281890
rect 287164 281832 287518 281888
rect 287574 281832 287579 281888
rect 287164 281830 287579 281832
rect 287164 281828 287170 281830
rect 287513 281827 287579 281830
rect 228449 281754 228515 281757
rect 228449 281752 240212 281754
rect 228449 281696 228454 281752
rect 228510 281696 240212 281752
rect 228449 281694 240212 281696
rect 228449 281691 228515 281694
rect 237782 281482 237788 281484
rect 109940 281422 237788 281482
rect 237782 281420 237788 281422
rect 237852 281420 237858 281484
rect 238150 281420 238156 281484
rect 238220 281482 238226 281484
rect 238661 281482 238727 281485
rect 238220 281480 238727 281482
rect 238220 281424 238666 281480
rect 238722 281424 238727 281480
rect 238220 281422 238727 281424
rect 238220 281420 238226 281422
rect 238661 281419 238727 281422
rect 237373 281210 237439 281213
rect 237373 281208 240212 281210
rect 237373 281152 237378 281208
rect 237434 281152 240212 281208
rect 237373 281150 240212 281152
rect 237373 281147 237439 281150
rect 237557 280666 237623 280669
rect 282821 280666 282887 280669
rect 237557 280664 240212 280666
rect 237557 280608 237562 280664
rect 237618 280608 240212 280664
rect 237557 280606 240212 280608
rect 279956 280664 282887 280666
rect 279956 280608 282826 280664
rect 282882 280608 282887 280664
rect 279956 280606 282887 280608
rect 237557 280603 237623 280606
rect 282821 280603 282887 280606
rect -960 279972 480 280212
rect 69151 280122 69217 280125
rect 74119 280122 74185 280125
rect 96521 280122 96587 280125
rect 69151 280120 71882 280122
rect 69151 280064 69156 280120
rect 69212 280064 71882 280120
rect 69151 280062 71882 280064
rect 69151 280059 69217 280062
rect 71822 279986 71882 280062
rect 74119 280120 96587 280122
rect 74119 280064 74124 280120
rect 74180 280064 96526 280120
rect 96582 280064 96587 280120
rect 74119 280062 96587 280064
rect 74119 280059 74185 280062
rect 96521 280059 96587 280062
rect 100615 280122 100681 280125
rect 115197 280122 115263 280125
rect 100615 280120 115263 280122
rect 100615 280064 100620 280120
rect 100676 280064 115202 280120
rect 115258 280064 115263 280120
rect 100615 280062 115263 280064
rect 100615 280059 100681 280062
rect 115197 280059 115263 280062
rect 237373 280122 237439 280125
rect 237373 280120 240212 280122
rect 237373 280064 237378 280120
rect 237434 280064 240212 280120
rect 237373 280062 240212 280064
rect 237373 280059 237439 280062
rect 78949 279986 79015 279989
rect 113817 279986 113883 279989
rect 71822 279984 79015 279986
rect 71822 279928 78954 279984
rect 79010 279928 79015 279984
rect 71822 279926 79015 279928
rect 78949 279923 79015 279926
rect 82678 279984 113883 279986
rect 82678 279928 113822 279984
rect 113878 279928 113883 279984
rect 82678 279926 113883 279928
rect 80743 279850 80809 279853
rect 82678 279850 82738 279926
rect 113817 279923 113883 279926
rect 111333 279850 111399 279853
rect 80743 279848 82738 279850
rect 80743 279792 80748 279848
rect 80804 279792 82738 279848
rect 80743 279790 82738 279792
rect 82862 279848 111399 279850
rect 82862 279792 111338 279848
rect 111394 279792 111399 279848
rect 82862 279790 111399 279792
rect 80743 279787 80809 279790
rect 71129 279714 71195 279717
rect 81433 279714 81499 279717
rect 71129 279712 81499 279714
rect 71129 279656 71134 279712
rect 71190 279656 81438 279712
rect 81494 279656 81499 279712
rect 71129 279654 81499 279656
rect 71129 279651 71195 279654
rect 81433 279651 81499 279654
rect 79409 279578 79475 279581
rect 82862 279578 82922 279790
rect 111333 279787 111399 279790
rect 82997 279714 83063 279717
rect 114001 279714 114067 279717
rect 82997 279712 114067 279714
rect 82997 279656 83002 279712
rect 83058 279656 114006 279712
rect 114062 279656 114067 279712
rect 82997 279654 114067 279656
rect 82997 279651 83063 279654
rect 114001 279651 114067 279654
rect 99373 279578 99439 279581
rect 79409 279576 82922 279578
rect 79409 279520 79414 279576
rect 79470 279520 82922 279576
rect 79409 279518 82922 279520
rect 83230 279576 99439 279578
rect 83230 279520 99378 279576
rect 99434 279520 99439 279576
rect 83230 279518 99439 279520
rect 79409 279515 79475 279518
rect 3366 279380 3372 279444
rect 3436 279442 3442 279444
rect 83089 279442 83155 279445
rect 3436 279440 83155 279442
rect 3436 279384 83094 279440
rect 83150 279384 83155 279440
rect 3436 279382 83155 279384
rect 3436 279380 3442 279382
rect 83089 279379 83155 279382
rect 75821 279306 75887 279309
rect 83230 279306 83290 279518
rect 99373 279515 99439 279518
rect 231485 279578 231551 279581
rect 231485 279576 240212 279578
rect 231485 279520 231490 279576
rect 231546 279520 240212 279576
rect 231485 279518 240212 279520
rect 231485 279515 231551 279518
rect 83365 279442 83431 279445
rect 122046 279442 122052 279444
rect 83365 279440 122052 279442
rect 83365 279384 83370 279440
rect 83426 279384 122052 279440
rect 83365 279382 122052 279384
rect 83365 279379 83431 279382
rect 122046 279380 122052 279382
rect 122116 279380 122122 279444
rect 120717 279306 120783 279309
rect 287513 279306 287579 279309
rect 75821 279304 83290 279306
rect 75821 279248 75826 279304
rect 75882 279248 83290 279304
rect 75821 279246 83290 279248
rect 84150 279304 120783 279306
rect 84150 279248 120722 279304
rect 120778 279248 120783 279304
rect 84150 279246 120783 279248
rect 279956 279304 287579 279306
rect 279956 279248 287518 279304
rect 287574 279248 287579 279304
rect 279956 279246 287579 279248
rect 75821 279243 75887 279246
rect 67541 279170 67607 279173
rect 78581 279170 78647 279173
rect 67541 279168 78647 279170
rect 67541 279112 67546 279168
rect 67602 279112 78586 279168
rect 78642 279112 78647 279168
rect 67541 279110 78647 279112
rect 67541 279107 67607 279110
rect 78581 279107 78647 279110
rect 72785 279034 72851 279037
rect 80053 279034 80119 279037
rect 72785 279032 80119 279034
rect 72785 278976 72790 279032
rect 72846 278976 80058 279032
rect 80114 278976 80119 279032
rect 72785 278974 80119 278976
rect 72785 278971 72851 278974
rect 80053 278971 80119 278974
rect 77753 278898 77819 278901
rect 84150 278898 84210 279246
rect 120717 279243 120783 279246
rect 287513 279243 287579 279246
rect 95969 279170 96035 279173
rect 112621 279170 112687 279173
rect 95969 279168 112687 279170
rect 95969 279112 95974 279168
rect 96030 279112 112626 279168
rect 112682 279112 112687 279168
rect 95969 279110 112687 279112
rect 95969 279107 96035 279110
rect 112621 279107 112687 279110
rect 230933 279034 230999 279037
rect 230933 279032 240212 279034
rect 230933 278976 230938 279032
rect 230994 278976 240212 279032
rect 230933 278974 240212 278976
rect 230933 278971 230999 278974
rect 77753 278896 84210 278898
rect 77753 278840 77758 278896
rect 77814 278840 84210 278896
rect 77753 278838 84210 278840
rect 77753 278835 77819 278838
rect 54569 278762 54635 278765
rect 91093 278762 91159 278765
rect 54569 278760 91159 278762
rect 54569 278704 54574 278760
rect 54630 278704 91098 278760
rect 91154 278704 91159 278760
rect 54569 278702 91159 278704
rect 54569 278699 54635 278702
rect 91093 278699 91159 278702
rect 92381 278762 92447 278765
rect 107377 278762 107443 278765
rect 92381 278760 107443 278762
rect 92381 278704 92386 278760
rect 92442 278704 107382 278760
rect 107438 278704 107443 278760
rect 92381 278702 107443 278704
rect 92381 278699 92447 278702
rect 107377 278699 107443 278702
rect 107561 278762 107627 278765
rect 111057 278762 111123 278765
rect 107561 278760 111123 278762
rect 107561 278704 107566 278760
rect 107622 278704 111062 278760
rect 111118 278704 111123 278760
rect 107561 278702 111123 278704
rect 107561 278699 107627 278702
rect 111057 278699 111123 278702
rect 56225 278626 56291 278629
rect 89713 278626 89779 278629
rect 56225 278624 89779 278626
rect 56225 278568 56230 278624
rect 56286 278568 89718 278624
rect 89774 278568 89779 278624
rect 56225 278566 89779 278568
rect 56225 278563 56291 278566
rect 89713 278563 89779 278566
rect 108941 278626 109007 278629
rect 126329 278626 126395 278629
rect 108941 278624 126395 278626
rect 108941 278568 108946 278624
rect 109002 278568 126334 278624
rect 126390 278568 126395 278624
rect 108941 278566 126395 278568
rect 108941 278563 109007 278566
rect 126329 278563 126395 278566
rect 89345 278490 89411 278493
rect 102133 278490 102199 278493
rect 89345 278488 102199 278490
rect 89345 278432 89350 278488
rect 89406 278432 102138 278488
rect 102194 278432 102199 278488
rect 89345 278430 102199 278432
rect 89345 278427 89411 278430
rect 102133 278427 102199 278430
rect 104249 278490 104315 278493
rect 119429 278490 119495 278493
rect 104249 278488 119495 278490
rect 104249 278432 104254 278488
rect 104310 278432 119434 278488
rect 119490 278432 119495 278488
rect 104249 278430 119495 278432
rect 104249 278427 104315 278430
rect 119429 278427 119495 278430
rect 231117 278490 231183 278493
rect 231117 278488 240212 278490
rect 231117 278432 231122 278488
rect 231178 278432 240212 278488
rect 231117 278430 240212 278432
rect 231117 278427 231183 278430
rect 91001 278354 91067 278357
rect 106181 278354 106247 278357
rect 91001 278352 106247 278354
rect 91001 278296 91006 278352
rect 91062 278296 106186 278352
rect 106242 278296 106247 278352
rect 91001 278294 106247 278296
rect 91001 278291 91067 278294
rect 106181 278291 106247 278294
rect 94313 278218 94379 278221
rect 108297 278218 108363 278221
rect 94313 278216 108363 278218
rect 94313 278160 94318 278216
rect 94374 278160 108302 278216
rect 108358 278160 108363 278216
rect 94313 278158 108363 278160
rect 94313 278155 94379 278158
rect 108297 278155 108363 278158
rect 84101 278082 84167 278085
rect 97901 278082 97967 278085
rect 84101 278080 97967 278082
rect 84101 278024 84106 278080
rect 84162 278024 97906 278080
rect 97962 278024 97967 278080
rect 84101 278022 97967 278024
rect 84101 278019 84167 278022
rect 97901 278019 97967 278022
rect 99281 278082 99347 278085
rect 111425 278082 111491 278085
rect 99281 278080 111491 278082
rect 99281 278024 99286 278080
rect 99342 278024 111430 278080
rect 111486 278024 111491 278080
rect 99281 278022 111491 278024
rect 99281 278019 99347 278022
rect 111425 278019 111491 278022
rect 64505 277946 64571 277949
rect 95141 277946 95207 277949
rect 64505 277944 95207 277946
rect 64505 277888 64510 277944
rect 64566 277888 95146 277944
rect 95202 277888 95207 277944
rect 64505 277886 95207 277888
rect 64505 277883 64571 277886
rect 95141 277883 95207 277886
rect 97625 277946 97691 277949
rect 117957 277946 118023 277949
rect 97625 277944 118023 277946
rect 97625 277888 97630 277944
rect 97686 277888 117962 277944
rect 118018 277888 118023 277944
rect 97625 277886 118023 277888
rect 97625 277883 97691 277886
rect 117957 277883 118023 277886
rect 231301 277946 231367 277949
rect 287605 277946 287671 277949
rect 231301 277944 240212 277946
rect 231301 277888 231306 277944
rect 231362 277888 240212 277944
rect 231301 277886 240212 277888
rect 279956 277944 287671 277946
rect 279956 277888 287610 277944
rect 287666 277888 287671 277944
rect 279956 277886 287671 277888
rect 231301 277883 231367 277886
rect 287605 277883 287671 277886
rect 86033 277810 86099 277813
rect 98637 277810 98703 277813
rect 86033 277808 98703 277810
rect 86033 277752 86038 277808
rect 86094 277752 98642 277808
rect 98698 277752 98703 277808
rect 86033 277750 98703 277752
rect 86033 277747 86099 277750
rect 98637 277747 98703 277750
rect 105905 277810 105971 277813
rect 116577 277810 116643 277813
rect 105905 277808 116643 277810
rect 105905 277752 105910 277808
rect 105966 277752 116582 277808
rect 116638 277752 116643 277808
rect 105905 277750 116643 277752
rect 105905 277747 105971 277750
rect 116577 277747 116643 277750
rect 87689 277674 87755 277677
rect 104801 277674 104867 277677
rect 87689 277672 104867 277674
rect 87689 277616 87694 277672
rect 87750 277616 104806 277672
rect 104862 277616 104867 277672
rect 87689 277614 104867 277616
rect 87689 277611 87755 277614
rect 104801 277611 104867 277614
rect 102593 277538 102659 277541
rect 111241 277538 111307 277541
rect 102593 277536 111307 277538
rect 102593 277480 102598 277536
rect 102654 277480 111246 277536
rect 111302 277480 111307 277536
rect 102593 277478 111307 277480
rect 102593 277475 102659 277478
rect 111241 277475 111307 277478
rect 52913 277402 52979 277405
rect 134517 277402 134583 277405
rect 52913 277400 134583 277402
rect 52913 277344 52918 277400
rect 52974 277344 134522 277400
rect 134578 277344 134583 277400
rect 52913 277342 134583 277344
rect 52913 277339 52979 277342
rect 134517 277339 134583 277342
rect 235901 277402 235967 277405
rect 235901 277400 240212 277402
rect 235901 277344 235906 277400
rect 235962 277344 240212 277400
rect 235901 277342 240212 277344
rect 235901 277339 235967 277342
rect 66161 277266 66227 277269
rect 140037 277266 140103 277269
rect 66161 277264 140103 277266
rect 66161 277208 66166 277264
rect 66222 277208 140042 277264
rect 140098 277208 140103 277264
rect 66161 277206 140103 277208
rect 66161 277203 66227 277206
rect 140037 277203 140103 277206
rect 57697 277130 57763 277133
rect 130377 277130 130443 277133
rect 57697 277128 130443 277130
rect 57697 277072 57702 277128
rect 57758 277072 130382 277128
rect 130438 277072 130443 277128
rect 57697 277070 130443 277072
rect 57697 277067 57763 277070
rect 130377 277067 130443 277070
rect 59261 276994 59327 276997
rect 127709 276994 127775 276997
rect 59261 276992 127775 276994
rect 59261 276936 59266 276992
rect 59322 276936 127714 276992
rect 127770 276936 127775 276992
rect 59261 276934 127775 276936
rect 59261 276931 59327 276934
rect 127709 276931 127775 276934
rect 61193 276858 61259 276861
rect 123661 276858 123727 276861
rect 61193 276856 123727 276858
rect 61193 276800 61198 276856
rect 61254 276800 123666 276856
rect 123722 276800 123727 276856
rect 61193 276798 123727 276800
rect 61193 276795 61259 276798
rect 123661 276795 123727 276798
rect 235022 276796 235028 276860
rect 235092 276858 235098 276860
rect 235092 276798 240212 276858
rect 235092 276796 235098 276798
rect 62849 276722 62915 276725
rect 122097 276722 122163 276725
rect 62849 276720 122163 276722
rect 62849 276664 62854 276720
rect 62910 276664 122102 276720
rect 122158 276664 122163 276720
rect 62849 276662 122163 276664
rect 62849 276659 62915 276662
rect 122097 276659 122163 276662
rect 282862 276586 282868 276588
rect 279956 276526 282868 276586
rect 282862 276524 282868 276526
rect 282932 276524 282938 276588
rect 227069 276314 227135 276317
rect 227069 276312 240212 276314
rect 227069 276256 227074 276312
rect 227130 276256 240212 276312
rect 227069 276254 240212 276256
rect 227069 276251 227135 276254
rect 155217 275770 155283 275773
rect 155217 275768 240212 275770
rect 155217 275712 155222 275768
rect 155278 275712 240212 275768
rect 155217 275710 240212 275712
rect 155217 275707 155283 275710
rect 199469 275226 199535 275229
rect 283005 275226 283071 275229
rect 199469 275224 240212 275226
rect 199469 275168 199474 275224
rect 199530 275168 240212 275224
rect 199469 275166 240212 275168
rect 279956 275224 283071 275226
rect 279956 275168 283010 275224
rect 283066 275168 283071 275224
rect 279956 275166 283071 275168
rect 199469 275163 199535 275166
rect 283005 275163 283071 275166
rect 173014 274620 173020 274684
rect 173084 274682 173090 274684
rect 173084 274622 240212 274682
rect 173084 274620 173090 274622
rect 282126 274620 282132 274684
rect 282196 274682 282202 274684
rect 283833 274682 283899 274685
rect 282196 274680 283899 274682
rect 282196 274624 283838 274680
rect 283894 274624 283899 274680
rect 282196 274622 283899 274624
rect 282196 274620 282202 274622
rect 283833 274619 283899 274622
rect 208894 274076 208900 274140
rect 208964 274138 208970 274140
rect 208964 274078 240212 274138
rect 208964 274076 208970 274078
rect 282821 273866 282887 273869
rect 279956 273864 282887 273866
rect 279956 273808 282826 273864
rect 282882 273808 282887 273864
rect 279956 273806 282887 273808
rect 282821 273803 282887 273806
rect 166206 273532 166212 273596
rect 166276 273594 166282 273596
rect 166276 273534 240212 273594
rect 166276 273532 166282 273534
rect 223062 272988 223068 273052
rect 223132 273050 223138 273052
rect 223132 272990 240212 273050
rect 223132 272988 223138 272990
rect 98637 272642 98703 272645
rect 222837 272642 222903 272645
rect 98637 272640 222903 272642
rect 98637 272584 98642 272640
rect 98698 272584 222842 272640
rect 222898 272584 222903 272640
rect 98637 272582 222903 272584
rect 98637 272579 98703 272582
rect 222837 272579 222903 272582
rect 203374 272444 203380 272508
rect 203444 272506 203450 272508
rect 282821 272506 282887 272509
rect 203444 272446 240212 272506
rect 279956 272504 282887 272506
rect 279956 272448 282826 272504
rect 282882 272448 282887 272504
rect 279956 272446 282887 272448
rect 203444 272444 203450 272446
rect 282821 272443 282887 272446
rect 580390 272172 580396 272236
rect 580460 272234 580466 272236
rect 583520 272234 584960 272324
rect 580460 272174 584960 272234
rect 580460 272172 580466 272174
rect 583520 272084 584960 272174
rect 225597 271962 225663 271965
rect 225597 271960 240212 271962
rect 225597 271904 225602 271960
rect 225658 271904 240212 271960
rect 225597 271902 240212 271904
rect 225597 271899 225663 271902
rect 235574 271356 235580 271420
rect 235644 271418 235650 271420
rect 235644 271358 240212 271418
rect 235644 271356 235650 271358
rect 295333 271146 295399 271149
rect 279956 271144 295399 271146
rect 279956 271088 295338 271144
rect 295394 271088 295399 271144
rect 279956 271086 295399 271088
rect 295333 271083 295399 271086
rect 18229 269786 18295 269789
rect 229829 269786 229895 269789
rect 292573 269786 292639 269789
rect 18229 269784 229895 269786
rect 18229 269728 18234 269784
rect 18290 269728 229834 269784
rect 229890 269728 229895 269784
rect 18229 269726 229895 269728
rect 279956 269784 292639 269786
rect 279956 269728 292578 269784
rect 292634 269728 292639 269784
rect 279956 269726 292639 269728
rect 18229 269723 18295 269726
rect 229829 269723 229895 269726
rect 292573 269723 292639 269726
rect 23013 268426 23079 268429
rect 224309 268426 224375 268429
rect 294045 268426 294111 268429
rect 23013 268424 224375 268426
rect 23013 268368 23018 268424
rect 23074 268368 224314 268424
rect 224370 268368 224375 268424
rect 23013 268366 224375 268368
rect 279956 268424 294111 268426
rect 279956 268368 294050 268424
rect 294106 268368 294111 268424
rect 279956 268366 294111 268368
rect 23013 268363 23079 268366
rect 224309 268363 224375 268366
rect 294045 268363 294111 268366
rect -960 267202 480 267292
rect 3417 267202 3483 267205
rect -960 267200 3483 267202
rect -960 267144 3422 267200
rect 3478 267144 3483 267200
rect -960 267142 3483 267144
rect -960 267052 480 267142
rect 3417 267139 3483 267142
rect 293953 267066 294019 267069
rect 279956 267064 294019 267066
rect 279956 267008 293958 267064
rect 294014 267008 294019 267064
rect 279956 267006 294019 267008
rect 293953 267003 294019 267006
rect 302877 265706 302943 265709
rect 279956 265704 302943 265706
rect 279956 265648 302882 265704
rect 302938 265648 302943 265704
rect 279956 265646 302943 265648
rect 302877 265643 302943 265646
rect 123477 265570 123543 265573
rect 216121 265570 216187 265573
rect 123477 265568 216187 265570
rect 123477 265512 123482 265568
rect 123538 265512 216126 265568
rect 216182 265512 216187 265568
rect 123477 265510 216187 265512
rect 123477 265507 123543 265510
rect 216121 265507 216187 265510
rect 298737 264346 298803 264349
rect 279956 264344 298803 264346
rect 279956 264288 298742 264344
rect 298798 264288 298803 264344
rect 279956 264286 298803 264288
rect 298737 264283 298803 264286
rect 31293 264210 31359 264213
rect 225689 264210 225755 264213
rect 31293 264208 225755 264210
rect 31293 264152 31298 264208
rect 31354 264152 225694 264208
rect 225750 264152 225755 264208
rect 31293 264150 225755 264152
rect 31293 264147 31359 264150
rect 225689 264147 225755 264150
rect 295977 262986 296043 262989
rect 279956 262984 296043 262986
rect 279956 262928 295982 262984
rect 296038 262928 296043 262984
rect 279956 262926 296043 262928
rect 295977 262923 296043 262926
rect 353937 261626 354003 261629
rect 279956 261624 354003 261626
rect 279956 261568 353942 261624
rect 353998 261568 354003 261624
rect 279956 261566 354003 261568
rect 353937 261563 354003 261566
rect 355174 260266 355180 260268
rect 279956 260206 355180 260266
rect 355174 260204 355180 260206
rect 355244 260204 355250 260268
rect 306966 258906 306972 258908
rect 279956 258846 306972 258906
rect 306966 258844 306972 258846
rect 307036 258844 307042 258908
rect 320766 258844 320772 258908
rect 320836 258906 320842 258908
rect 583520 258906 584960 258996
rect 320836 258846 584960 258906
rect 320836 258844 320842 258846
rect 583520 258756 584960 258846
rect 313774 257546 313780 257548
rect 279956 257486 313780 257546
rect 313774 257484 313780 257486
rect 313844 257484 313850 257548
rect 309726 256186 309732 256188
rect 279956 256126 309732 256186
rect 309726 256124 309732 256126
rect 309796 256124 309802 256188
rect 574686 254826 574692 254828
rect 279956 254766 574692 254826
rect 574686 254764 574692 254766
rect 574756 254764 574762 254828
rect -960 254146 480 254236
rect 3366 254146 3372 254148
rect -960 254086 3372 254146
rect -960 253996 480 254086
rect 3366 254084 3372 254086
rect 3436 254084 3442 254148
rect 500166 253466 500172 253468
rect 279956 253406 500172 253466
rect 500166 253404 500172 253406
rect 500236 253404 500242 253468
rect 299974 252106 299980 252108
rect 279956 252046 299980 252106
rect 299974 252044 299980 252046
rect 300044 252044 300050 252108
rect 544326 250746 544332 250748
rect 279956 250686 544332 250746
rect 544326 250684 544332 250686
rect 544396 250684 544402 250748
rect 320766 249386 320772 249388
rect 279956 249326 320772 249386
rect 320766 249324 320772 249326
rect 320836 249324 320842 249388
rect 355174 248026 355180 248028
rect 279956 247966 355180 248026
rect 355174 247964 355180 247966
rect 355244 247964 355250 248028
rect 353886 246666 353892 246668
rect 279956 246606 353892 246666
rect 353886 246604 353892 246606
rect 353956 246604 353962 246668
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 346894 245306 346900 245308
rect 279956 245246 346900 245306
rect 346894 245244 346900 245246
rect 346964 245244 346970 245308
rect 34789 244898 34855 244901
rect 186957 244898 187023 244901
rect 34789 244896 187023 244898
rect 34789 244840 34794 244896
rect 34850 244840 186962 244896
rect 187018 244840 187023 244896
rect 34789 244838 187023 244840
rect 34789 244835 34855 244838
rect 186957 244835 187023 244838
rect 500166 243946 500172 243948
rect 279956 243886 500172 243946
rect 500166 243884 500172 243886
rect 500236 243884 500242 243948
rect 105721 243538 105787 243541
rect 202137 243538 202203 243541
rect 105721 243536 202203 243538
rect 105721 243480 105726 243536
rect 105782 243480 202142 243536
rect 202198 243480 202203 243536
rect 105721 243478 202203 243480
rect 105721 243475 105787 243478
rect 202137 243475 202203 243478
rect 559414 242586 559420 242588
rect 279956 242526 559420 242586
rect 559414 242524 559420 242526
rect 559484 242524 559490 242588
rect 231342 242178 231348 242180
rect 6870 242118 231348 242178
rect 6870 241634 6930 242118
rect 231342 242116 231348 242118
rect 231412 242116 231418 242180
rect 279550 241844 279556 241908
rect 279620 241906 279626 241908
rect 280061 241906 280127 241909
rect 279620 241904 280127 241906
rect 279620 241848 280066 241904
rect 280122 241848 280127 241904
rect 279620 241846 280127 241848
rect 279620 241844 279626 241846
rect 280061 241843 280127 241846
rect 280061 241770 280127 241773
rect 282361 241770 282427 241773
rect 280061 241768 282427 241770
rect 280061 241712 280066 241768
rect 280122 241712 282366 241768
rect 282422 241712 282427 241768
rect 280061 241710 282427 241712
rect 280061 241707 280127 241710
rect 282361 241707 282427 241710
rect 3374 241574 6930 241634
rect -960 241090 480 241180
rect 3374 241090 3434 241574
rect 287094 241436 287100 241500
rect 287164 241498 287170 241500
rect 287421 241498 287487 241501
rect 287164 241496 287487 241498
rect 287164 241440 287426 241496
rect 287482 241440 287487 241496
rect 287164 241438 287487 241440
rect 287164 241436 287170 241438
rect 287421 241435 287487 241438
rect 457294 241226 457300 241228
rect 279956 241166 457300 241226
rect 457294 241164 457300 241166
rect 457364 241164 457370 241228
rect -960 241030 3434 241090
rect -960 240940 480 241030
rect 282269 240954 282335 240957
rect 287646 240954 287652 240956
rect 282269 240952 287652 240954
rect 282269 240896 282274 240952
rect 282330 240896 287652 240952
rect 282269 240894 287652 240896
rect 282269 240891 282335 240894
rect 287646 240892 287652 240894
rect 287716 240892 287722 240956
rect 3366 240620 3372 240684
rect 3436 240682 3442 240684
rect 283230 240682 283236 240684
rect 3436 240622 283236 240682
rect 3436 240620 3442 240622
rect 283230 240620 283236 240622
rect 283300 240620 283306 240684
rect 235390 240484 235396 240548
rect 235460 240546 235466 240548
rect 287278 240546 287284 240548
rect 235460 240486 287284 240546
rect 235460 240484 235466 240486
rect 287278 240484 287284 240486
rect 287348 240484 287354 240548
rect 237782 240348 237788 240412
rect 237852 240410 237858 240412
rect 282269 240410 282335 240413
rect 237852 240408 282335 240410
rect 237852 240352 282274 240408
rect 282330 240352 282335 240408
rect 237852 240350 282335 240352
rect 237852 240348 237858 240350
rect 282269 240347 282335 240350
rect 238661 240274 238727 240277
rect 580257 240274 580323 240277
rect 238661 240272 580323 240274
rect 238661 240216 238666 240272
rect 238722 240216 580262 240272
rect 580318 240216 580323 240272
rect 238661 240214 580323 240216
rect 238661 240211 238727 240214
rect 580257 240211 580323 240214
rect 284477 240138 284543 240141
rect 284702 240138 284708 240140
rect 284477 240136 284708 240138
rect 284477 240080 284482 240136
rect 284538 240080 284708 240136
rect 284477 240078 284708 240080
rect 284477 240075 284543 240078
rect 284702 240076 284708 240078
rect 284772 240076 284778 240140
rect 238518 239940 238524 240004
rect 238588 240002 238594 240004
rect 580206 240002 580212 240004
rect 238588 239942 580212 240002
rect 238588 239940 238594 239942
rect 580206 239940 580212 239942
rect 580276 239940 580282 240004
rect 48630 239804 48636 239868
rect 48700 239866 48706 239868
rect 287830 239866 287836 239868
rect 48700 239806 287836 239866
rect 48700 239804 48706 239806
rect 287830 239804 287836 239806
rect 287900 239804 287906 239868
rect 237966 239668 237972 239732
rect 238036 239730 238042 239732
rect 287462 239730 287468 239732
rect 238036 239670 287468 239730
rect 238036 239668 238042 239670
rect 287462 239668 287468 239670
rect 287532 239668 287538 239732
rect 101397 239594 101463 239597
rect 186313 239594 186379 239597
rect 101397 239592 186379 239594
rect 101397 239536 101402 239592
rect 101458 239536 186318 239592
rect 186374 239536 186379 239592
rect 101397 239534 186379 239536
rect 101397 239531 101463 239534
rect 186313 239531 186379 239534
rect 237005 239594 237071 239597
rect 280429 239594 280495 239597
rect 237005 239592 280495 239594
rect 237005 239536 237010 239592
rect 237066 239536 280434 239592
rect 280490 239536 280495 239592
rect 237005 239534 280495 239536
rect 237005 239531 237071 239534
rect 280429 239531 280495 239534
rect 176653 239458 176719 239461
rect 237373 239458 237439 239461
rect 176653 239456 237439 239458
rect 176653 239400 176658 239456
rect 176714 239400 237378 239456
rect 237434 239400 237439 239456
rect 176653 239398 237439 239400
rect 176653 239395 176719 239398
rect 237373 239395 237439 239398
rect 258257 239458 258323 239461
rect 288893 239458 288959 239461
rect 258257 239456 288959 239458
rect 258257 239400 258262 239456
rect 258318 239400 288898 239456
rect 288954 239400 288959 239456
rect 258257 239398 288959 239400
rect 258257 239395 258323 239398
rect 288893 239395 288959 239398
rect 148317 239322 148383 239325
rect 212441 239322 212507 239325
rect 148317 239320 212507 239322
rect 148317 239264 148322 239320
rect 148378 239264 212446 239320
rect 212502 239264 212507 239320
rect 148317 239262 212507 239264
rect 148317 239259 148383 239262
rect 212441 239259 212507 239262
rect 212717 239322 212783 239325
rect 264973 239322 265039 239325
rect 212717 239320 265039 239322
rect 212717 239264 212722 239320
rect 212778 239264 264978 239320
rect 265034 239264 265039 239320
rect 212717 239262 265039 239264
rect 212717 239259 212783 239262
rect 264973 239259 265039 239262
rect 173157 239186 173223 239189
rect 237465 239186 237531 239189
rect 173157 239184 237531 239186
rect 173157 239128 173162 239184
rect 173218 239128 237470 239184
rect 237526 239128 237531 239184
rect 173157 239126 237531 239128
rect 173157 239123 173223 239126
rect 237465 239123 237531 239126
rect 265341 239186 265407 239189
rect 280153 239186 280219 239189
rect 265341 239184 280219 239186
rect 265341 239128 265346 239184
rect 265402 239128 280158 239184
rect 280214 239128 280219 239184
rect 265341 239126 280219 239128
rect 265341 239123 265407 239126
rect 280153 239123 280219 239126
rect 158897 239050 158963 239053
rect 235993 239050 236059 239053
rect 158897 239048 236059 239050
rect 158897 238992 158902 239048
rect 158958 238992 235998 239048
rect 236054 238992 236059 239048
rect 158897 238990 236059 238992
rect 158897 238987 158963 238990
rect 235993 238987 236059 238990
rect 238334 238988 238340 239052
rect 238404 239050 238410 239052
rect 580390 239050 580396 239052
rect 238404 238990 580396 239050
rect 238404 238988 238410 238990
rect 580390 238988 580396 238990
rect 580460 238988 580466 239052
rect 180241 238914 180307 238917
rect 237557 238914 237623 238917
rect 180241 238912 237623 238914
rect 180241 238856 180246 238912
rect 180302 238856 237562 238912
rect 237618 238856 237623 238912
rect 180241 238854 237623 238856
rect 180241 238851 180307 238854
rect 237557 238851 237623 238854
rect 35985 238778 36051 238781
rect 179413 238778 179479 238781
rect 35985 238776 179479 238778
rect 35985 238720 35990 238776
rect 36046 238720 179418 238776
rect 179474 238720 179479 238776
rect 35985 238718 179479 238720
rect 35985 238715 36051 238718
rect 179413 238715 179479 238718
rect 187325 238778 187391 238781
rect 259269 238778 259335 238781
rect 187325 238776 259335 238778
rect 187325 238720 187330 238776
rect 187386 238720 259274 238776
rect 259330 238720 259335 238776
rect 187325 238718 259335 238720
rect 187325 238715 187391 238718
rect 259269 238715 259335 238718
rect 44265 238642 44331 238645
rect 252185 238642 252251 238645
rect 44265 238640 252251 238642
rect 44265 238584 44270 238640
rect 44326 238584 252190 238640
rect 252246 238584 252251 238640
rect 44265 238582 252251 238584
rect 44265 238579 44331 238582
rect 252185 238579 252251 238582
rect 40677 238506 40743 238509
rect 250989 238506 251055 238509
rect 40677 238504 251055 238506
rect 40677 238448 40682 238504
rect 40738 238448 250994 238504
rect 251050 238448 251055 238504
rect 40677 238446 251055 238448
rect 40677 238443 40743 238446
rect 250989 238443 251055 238446
rect 37181 238370 37247 238373
rect 249793 238370 249859 238373
rect 37181 238368 249859 238370
rect 37181 238312 37186 238368
rect 37242 238312 249798 238368
rect 249854 238312 249859 238368
rect 37181 238310 249859 238312
rect 37181 238307 37247 238310
rect 249793 238307 249859 238310
rect 261753 238370 261819 238373
rect 283097 238370 283163 238373
rect 261753 238368 283163 238370
rect 261753 238312 261758 238368
rect 261814 238312 283102 238368
rect 283158 238312 283163 238368
rect 261753 238310 283163 238312
rect 261753 238307 261819 238310
rect 283097 238307 283163 238310
rect 33593 238234 33659 238237
rect 248597 238234 248663 238237
rect 33593 238232 248663 238234
rect 33593 238176 33598 238232
rect 33654 238176 248602 238232
rect 248658 238176 248663 238232
rect 33593 238174 248663 238176
rect 33593 238171 33659 238174
rect 248597 238171 248663 238174
rect 251173 238234 251239 238237
rect 280245 238234 280311 238237
rect 251173 238232 280311 238234
rect 251173 238176 251178 238232
rect 251234 238176 280250 238232
rect 280306 238176 280311 238232
rect 251173 238174 280311 238176
rect 251173 238171 251239 238174
rect 280245 238171 280311 238174
rect 30097 238098 30163 238101
rect 247401 238098 247467 238101
rect 30097 238096 247467 238098
rect 30097 238040 30102 238096
rect 30158 238040 247406 238096
rect 247462 238040 247467 238096
rect 30097 238038 247467 238040
rect 30097 238035 30163 238038
rect 247401 238035 247467 238038
rect 254669 238098 254735 238101
rect 284845 238098 284911 238101
rect 254669 238096 284911 238098
rect 254669 238040 254674 238096
rect 254730 238040 284850 238096
rect 284906 238040 284911 238096
rect 254669 238038 284911 238040
rect 254669 238035 254735 238038
rect 284845 238035 284911 238038
rect 26509 237962 26575 237965
rect 246205 237962 246271 237965
rect 26509 237960 246271 237962
rect 26509 237904 26514 237960
rect 26570 237904 246210 237960
rect 246266 237904 246271 237960
rect 26509 237902 246271 237904
rect 26509 237899 26575 237902
rect 246205 237899 246271 237902
rect 247585 237962 247651 237965
rect 281717 237962 281783 237965
rect 247585 237960 281783 237962
rect 247585 237904 247590 237960
rect 247646 237904 281722 237960
rect 281778 237904 281783 237960
rect 247585 237902 281783 237904
rect 247585 237899 247651 237902
rect 281717 237899 281783 237902
rect 122281 237826 122347 237829
rect 278497 237826 278563 237829
rect 122281 237824 278563 237826
rect 122281 237768 122286 237824
rect 122342 237768 278502 237824
rect 278558 237768 278563 237824
rect 122281 237766 278563 237768
rect 122281 237763 122347 237766
rect 278497 237763 278563 237766
rect 17033 237554 17099 237557
rect 44173 237554 44239 237557
rect 17033 237552 44239 237554
rect 17033 237496 17038 237552
rect 17094 237496 44178 237552
rect 44234 237496 44239 237552
rect 17033 237494 44239 237496
rect 17033 237491 17099 237494
rect 44173 237491 44239 237494
rect 21817 237418 21883 237421
rect 121453 237418 121519 237421
rect 21817 237416 121519 237418
rect 21817 237360 21822 237416
rect 21878 237360 121458 237416
rect 121514 237360 121519 237416
rect 21817 237358 121519 237360
rect 21817 237355 21883 237358
rect 121453 237355 121519 237358
rect 233417 237146 233483 237149
rect 285121 237146 285187 237149
rect 233417 237144 285187 237146
rect 233417 237088 233422 237144
rect 233478 237088 285126 237144
rect 285182 237088 285187 237144
rect 233417 237086 285187 237088
rect 233417 237083 233483 237086
rect 285121 237083 285187 237086
rect 201493 237010 201559 237013
rect 281993 237010 282059 237013
rect 201493 237008 282059 237010
rect 201493 236952 201498 237008
rect 201554 236952 281998 237008
rect 282054 236952 282059 237008
rect 201493 236950 282059 236952
rect 201493 236947 201559 236950
rect 281993 236947 282059 236950
rect 162485 236874 162551 236877
rect 283557 236874 283623 236877
rect 162485 236872 283623 236874
rect 162485 236816 162490 236872
rect 162546 236816 283562 236872
rect 283618 236816 283623 236872
rect 162485 236814 283623 236816
rect 162485 236811 162551 236814
rect 283557 236811 283623 236814
rect 114001 236738 114067 236741
rect 286501 236738 286567 236741
rect 114001 236736 286567 236738
rect 114001 236680 114006 236736
rect 114062 236680 286506 236736
rect 286562 236680 286567 236736
rect 114001 236678 286567 236680
rect 114001 236675 114067 236678
rect 286501 236675 286567 236678
rect 239765 236602 239831 236605
rect 580257 236602 580323 236605
rect 239765 236600 580323 236602
rect 239765 236544 239770 236600
rect 239826 236544 580262 236600
rect 580318 236544 580323 236600
rect 239765 236542 580323 236544
rect 239765 236539 239831 236542
rect 580257 236539 580323 236542
rect 183737 235650 183803 235653
rect 280705 235650 280771 235653
rect 183737 235648 280771 235650
rect 183737 235592 183742 235648
rect 183798 235592 280710 235648
rect 280766 235592 280771 235648
rect 183737 235590 280771 235592
rect 183737 235587 183803 235590
rect 280705 235587 280771 235590
rect 141233 235514 141299 235517
rect 285213 235514 285279 235517
rect 141233 235512 285279 235514
rect 141233 235456 141238 235512
rect 141294 235456 285218 235512
rect 285274 235456 285279 235512
rect 141233 235454 285279 235456
rect 141233 235451 141299 235454
rect 285213 235451 285279 235454
rect 14733 235378 14799 235381
rect 284886 235378 284892 235380
rect 14733 235376 284892 235378
rect 14733 235320 14738 235376
rect 14794 235320 284892 235376
rect 14733 235318 284892 235320
rect 14733 235315 14799 235318
rect 284886 235316 284892 235318
rect 284956 235316 284962 235380
rect 239857 235242 239923 235245
rect 580349 235242 580415 235245
rect 239857 235240 580415 235242
rect 239857 235184 239862 235240
rect 239918 235184 580354 235240
rect 580410 235184 580415 235240
rect 239857 235182 580415 235184
rect 239857 235179 239923 235182
rect 580349 235179 580415 235182
rect 197905 234154 197971 234157
rect 283373 234154 283439 234157
rect 197905 234152 283439 234154
rect 197905 234096 197910 234152
rect 197966 234096 283378 234152
rect 283434 234096 283439 234152
rect 197905 234094 283439 234096
rect 197905 234091 197971 234094
rect 283373 234091 283439 234094
rect 106917 234018 106983 234021
rect 286409 234018 286475 234021
rect 106917 234016 286475 234018
rect 106917 233960 106922 234016
rect 106978 233960 286414 234016
rect 286470 233960 286475 234016
rect 106917 233958 286475 233960
rect 106917 233955 106983 233958
rect 286409 233955 286475 233958
rect 39573 233882 39639 233885
rect 281758 233882 281764 233884
rect 39573 233880 281764 233882
rect 39573 233824 39578 233880
rect 39634 233824 281764 233880
rect 39573 233822 281764 233824
rect 39573 233819 39639 233822
rect 281758 233820 281764 233822
rect 281828 233820 281834 233884
rect 208577 232794 208643 232797
rect 280521 232794 280587 232797
rect 208577 232792 280587 232794
rect 208577 232736 208582 232792
rect 208638 232736 280526 232792
rect 280582 232736 280587 232792
rect 208577 232734 280587 232736
rect 208577 232731 208643 232734
rect 280521 232731 280587 232734
rect 126973 232658 127039 232661
rect 283741 232658 283807 232661
rect 126973 232656 283807 232658
rect 126973 232600 126978 232656
rect 127034 232600 283746 232656
rect 283802 232600 283807 232656
rect 126973 232598 283807 232600
rect 126973 232595 127039 232598
rect 283741 232595 283807 232598
rect 121085 232522 121151 232525
rect 286133 232522 286199 232525
rect 121085 232520 286199 232522
rect 121085 232464 121090 232520
rect 121146 232464 286138 232520
rect 286194 232464 286199 232520
rect 121085 232462 286199 232464
rect 121085 232459 121151 232462
rect 286133 232459 286199 232462
rect 239254 232324 239260 232388
rect 239324 232386 239330 232388
rect 583520 232386 584960 232476
rect 239324 232326 584960 232386
rect 239324 232324 239330 232326
rect 583520 232236 584960 232326
rect 194409 231298 194475 231301
rect 280613 231298 280679 231301
rect 194409 231296 280679 231298
rect 194409 231240 194414 231296
rect 194470 231240 280618 231296
rect 280674 231240 280679 231296
rect 194409 231238 280679 231240
rect 194409 231235 194475 231238
rect 280613 231235 280679 231238
rect 155401 231162 155467 231165
rect 285029 231162 285095 231165
rect 155401 231160 285095 231162
rect 155401 231104 155406 231160
rect 155462 231104 285034 231160
rect 285090 231104 285095 231160
rect 155401 231102 285095 231104
rect 155401 231099 155467 231102
rect 285029 231099 285095 231102
rect 222745 230074 222811 230077
rect 280337 230074 280403 230077
rect 222745 230072 280403 230074
rect 222745 230016 222750 230072
rect 222806 230016 280342 230072
rect 280398 230016 280403 230072
rect 222745 230014 280403 230016
rect 222745 230011 222811 230014
rect 280337 230011 280403 230014
rect 190821 229938 190887 229941
rect 281901 229938 281967 229941
rect 190821 229936 281967 229938
rect 190821 229880 190826 229936
rect 190882 229880 281906 229936
rect 281962 229880 281967 229936
rect 190821 229878 281967 229880
rect 190821 229875 190887 229878
rect 281901 229875 281967 229878
rect 99833 229802 99899 229805
rect 286317 229802 286383 229805
rect 99833 229800 286383 229802
rect 99833 229744 99838 229800
rect 99894 229744 286322 229800
rect 286378 229744 286383 229800
rect 99833 229742 286383 229744
rect 99833 229739 99899 229742
rect 286317 229739 286383 229742
rect 229829 228578 229895 228581
rect 284569 228578 284635 228581
rect 229829 228576 284635 228578
rect 229829 228520 229834 228576
rect 229890 228520 284574 228576
rect 284630 228520 284635 228576
rect 229829 228518 284635 228520
rect 229829 228515 229895 228518
rect 284569 228515 284635 228518
rect 166073 228442 166139 228445
rect 283465 228442 283531 228445
rect 166073 228440 283531 228442
rect 166073 228384 166078 228440
rect 166134 228384 283470 228440
rect 283526 228384 283531 228440
rect 166073 228382 283531 228384
rect 166073 228379 166139 228382
rect 283465 228379 283531 228382
rect 43069 228306 43135 228309
rect 279366 228306 279372 228308
rect 43069 228304 279372 228306
rect 43069 228248 43074 228304
rect 43130 228248 279372 228304
rect 43069 228246 279372 228248
rect 43069 228243 43135 228246
rect 279366 228244 279372 228246
rect 279436 228244 279442 228308
rect -960 227884 480 228124
rect 103329 226946 103395 226949
rect 286225 226946 286291 226949
rect 103329 226944 286291 226946
rect 103329 226888 103334 226944
rect 103390 226888 286230 226944
rect 286286 226888 286291 226944
rect 103329 226886 286291 226888
rect 103329 226883 103395 226886
rect 286225 226883 286291 226886
rect 130561 225722 130627 225725
rect 283649 225722 283715 225725
rect 130561 225720 283715 225722
rect 130561 225664 130566 225720
rect 130622 225664 283654 225720
rect 283710 225664 283715 225720
rect 130561 225662 283715 225664
rect 130561 225659 130627 225662
rect 283649 225659 283715 225662
rect 24209 225586 24275 225589
rect 279550 225586 279556 225588
rect 24209 225584 279556 225586
rect 24209 225528 24214 225584
rect 24270 225528 279556 225584
rect 24209 225526 279556 225528
rect 24209 225523 24275 225526
rect 279550 225524 279556 225526
rect 279620 225524 279626 225588
rect 215661 224362 215727 224365
rect 284661 224362 284727 224365
rect 215661 224360 284727 224362
rect 215661 224304 215666 224360
rect 215722 224304 284666 224360
rect 284722 224304 284727 224360
rect 215661 224302 284727 224304
rect 215661 224299 215727 224302
rect 284661 224299 284727 224302
rect 87965 224226 88031 224229
rect 215937 224226 216003 224229
rect 87965 224224 216003 224226
rect 87965 224168 87970 224224
rect 88026 224168 215942 224224
rect 215998 224168 216003 224224
rect 87965 224166 216003 224168
rect 87965 224163 88031 224166
rect 215937 224163 216003 224166
rect 205081 223002 205147 223005
rect 283281 223002 283347 223005
rect 205081 223000 283347 223002
rect 205081 222944 205086 223000
rect 205142 222944 283286 223000
rect 283342 222944 283347 223000
rect 205081 222942 283347 222944
rect 205081 222939 205147 222942
rect 283281 222939 283347 222942
rect 110505 222866 110571 222869
rect 285857 222866 285923 222869
rect 110505 222864 285923 222866
rect 110505 222808 110510 222864
rect 110566 222808 285862 222864
rect 285918 222808 285923 222864
rect 110505 222806 285923 222808
rect 110505 222803 110571 222806
rect 285857 222803 285923 222806
rect 226333 221642 226399 221645
rect 284385 221642 284451 221645
rect 226333 221640 284451 221642
rect 226333 221584 226338 221640
rect 226394 221584 284390 221640
rect 284446 221584 284451 221640
rect 226333 221582 284451 221584
rect 226333 221579 226399 221582
rect 284385 221579 284451 221582
rect 96245 221506 96311 221509
rect 285949 221506 286015 221509
rect 96245 221504 286015 221506
rect 96245 221448 96250 221504
rect 96306 221448 285954 221504
rect 286010 221448 286015 221504
rect 96245 221446 286015 221448
rect 96245 221443 96311 221446
rect 285949 221443 286015 221446
rect 134149 220282 134215 220285
rect 280838 220282 280844 220284
rect 134149 220280 280844 220282
rect 134149 220224 134154 220280
rect 134210 220224 280844 220280
rect 134149 220222 280844 220224
rect 134149 220219 134215 220222
rect 280838 220220 280844 220222
rect 280908 220220 280914 220284
rect 92749 220146 92815 220149
rect 286041 220146 286107 220149
rect 92749 220144 286107 220146
rect 92749 220088 92754 220144
rect 92810 220088 286046 220144
rect 286102 220088 286107 220144
rect 92749 220086 286107 220088
rect 92749 220083 92815 220086
rect 286041 220083 286107 220086
rect 355174 218996 355180 219060
rect 355244 219058 355250 219060
rect 583520 219058 584960 219148
rect 355244 218998 584960 219058
rect 355244 218996 355250 218998
rect 583520 218908 584960 218998
rect 25497 218650 25563 218653
rect 281574 218650 281580 218652
rect 25497 218648 281580 218650
rect 25497 218592 25502 218648
rect 25558 218592 281580 218648
rect 25497 218590 281580 218592
rect 25497 218587 25563 218590
rect 281574 218588 281580 218590
rect 281644 218588 281650 218652
rect 3550 217228 3556 217292
rect 3620 217290 3626 217292
rect 283046 217290 283052 217292
rect 3620 217230 283052 217290
rect 3620 217228 3626 217230
rect 283046 217228 283052 217230
rect 283116 217228 283122 217292
rect 3734 215868 3740 215932
rect 3804 215930 3810 215932
rect 283414 215930 283420 215932
rect 3804 215870 283420 215930
rect 3804 215868 3810 215870
rect 283414 215868 283420 215870
rect 283484 215868 283490 215932
rect -960 214978 480 215068
rect 3417 214978 3483 214981
rect -960 214976 3483 214978
rect -960 214920 3422 214976
rect 3478 214920 3483 214976
rect -960 214918 3483 214920
rect -960 214828 480 214918
rect 3417 214915 3483 214918
rect 91737 214570 91803 214573
rect 282177 214570 282243 214573
rect 91737 214568 282243 214570
rect 91737 214512 91742 214568
rect 91798 214512 282182 214568
rect 282238 214512 282243 214568
rect 91737 214510 282243 214512
rect 91737 214507 91803 214510
rect 282177 214507 282243 214510
rect 90357 213210 90423 213213
rect 267733 213210 267799 213213
rect 90357 213208 267799 213210
rect 90357 213152 90362 213208
rect 90418 213152 267738 213208
rect 267794 213152 267799 213208
rect 90357 213150 267799 213152
rect 90357 213147 90423 213150
rect 267733 213147 267799 213150
rect 93945 211850 94011 211853
rect 268929 211850 268995 211853
rect 93945 211848 268995 211850
rect 93945 211792 93950 211848
rect 94006 211792 268934 211848
rect 268990 211792 268995 211848
rect 93945 211790 268995 211792
rect 93945 211787 94011 211790
rect 268929 211787 268995 211790
rect 97441 210354 97507 210357
rect 270125 210354 270191 210357
rect 97441 210352 270191 210354
rect 97441 210296 97446 210352
rect 97502 210296 270130 210352
rect 270186 210296 270191 210352
rect 97441 210294 270191 210296
rect 97441 210291 97507 210294
rect 270125 210291 270191 210294
rect 104525 208994 104591 208997
rect 272517 208994 272583 208997
rect 104525 208992 272583 208994
rect 104525 208936 104530 208992
rect 104586 208936 272522 208992
rect 272578 208936 272583 208992
rect 104525 208934 272583 208936
rect 104525 208931 104591 208934
rect 272517 208931 272583 208934
rect 115197 207634 115263 207637
rect 275277 207634 275343 207637
rect 115197 207632 275343 207634
rect 115197 207576 115202 207632
rect 115258 207576 275282 207632
rect 275338 207576 275343 207632
rect 115197 207574 275343 207576
rect 115197 207571 115263 207574
rect 275277 207571 275343 207574
rect 126237 206274 126303 206277
rect 277301 206274 277367 206277
rect 126237 206272 277367 206274
rect 126237 206216 126242 206272
rect 126298 206216 277306 206272
rect 277362 206216 277367 206272
rect 126237 206214 277367 206216
rect 126237 206211 126303 206214
rect 277301 206211 277367 206214
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect 85665 204914 85731 204917
rect 285765 204914 285831 204917
rect 85665 204912 285831 204914
rect 85665 204856 85670 204912
rect 85726 204856 285770 204912
rect 285826 204856 285831 204912
rect 85665 204854 285831 204856
rect 85665 204851 85731 204854
rect 285765 204851 285831 204854
rect 219249 203690 219315 203693
rect 284293 203690 284359 203693
rect 219249 203688 284359 203690
rect 219249 203632 219254 203688
rect 219310 203632 284298 203688
rect 284354 203632 284359 203688
rect 219249 203630 284359 203632
rect 219249 203627 219315 203630
rect 284293 203627 284359 203630
rect 32397 203554 32463 203557
rect 282085 203554 282151 203557
rect 32397 203552 282151 203554
rect 32397 203496 32402 203552
rect 32458 203496 282090 203552
rect 282146 203496 282151 203552
rect 32397 203494 282151 203496
rect 32397 203491 32463 203494
rect 282085 203491 282151 203494
rect 3366 202132 3372 202196
rect 3436 202194 3442 202196
rect 281022 202194 281028 202196
rect 3436 202134 281028 202194
rect 3436 202132 3442 202134
rect 281022 202132 281028 202134
rect 281092 202132 281098 202196
rect -960 201922 480 202012
rect 3734 201922 3740 201924
rect -960 201862 3740 201922
rect -960 201772 480 201862
rect 3734 201860 3740 201862
rect 3804 201860 3810 201924
rect 137645 200698 137711 200701
rect 284937 200698 285003 200701
rect 137645 200696 285003 200698
rect 137645 200640 137650 200696
rect 137706 200640 284942 200696
rect 284998 200640 285003 200696
rect 137645 200638 285003 200640
rect 137645 200635 137711 200638
rect 284937 200635 285003 200638
rect 144729 197978 144795 197981
rect 284753 197978 284819 197981
rect 144729 197976 284819 197978
rect 144729 197920 144734 197976
rect 144790 197920 284758 197976
rect 284814 197920 284819 197976
rect 144729 197918 284819 197920
rect 144729 197915 144795 197918
rect 284753 197915 284819 197918
rect 151813 196618 151879 196621
rect 283189 196618 283255 196621
rect 151813 196616 283255 196618
rect 151813 196560 151818 196616
rect 151874 196560 283194 196616
rect 283250 196560 283255 196616
rect 151813 196558 283255 196560
rect 151813 196555 151879 196558
rect 283189 196555 283255 196558
rect 239438 192476 239444 192540
rect 239508 192538 239514 192540
rect 583520 192538 584960 192628
rect 239508 192478 584960 192538
rect 239508 192476 239514 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 228214 188866 228220 188868
rect -960 188806 228220 188866
rect -960 188716 480 188806
rect 228214 188804 228220 188806
rect 228284 188804 228290 188868
rect 353886 179148 353892 179212
rect 353956 179210 353962 179212
rect 583520 179210 584960 179300
rect 353956 179150 584960 179210
rect 353956 179148 353962 179150
rect 583520 179060 584960 179150
rect 108113 178666 108179 178669
rect 273713 178666 273779 178669
rect 108113 178664 273779 178666
rect 108113 178608 108118 178664
rect 108174 178608 273718 178664
rect 273774 178608 273779 178664
rect 108113 178606 273779 178608
rect 108113 178603 108179 178606
rect 273713 178603 273779 178606
rect 101029 177306 101095 177309
rect 271321 177306 271387 177309
rect 101029 177304 271387 177306
rect 101029 177248 101034 177304
rect 101090 177248 271326 177304
rect 271382 177248 271387 177304
rect 101029 177246 271387 177248
rect 101029 177243 101095 177246
rect 271321 177243 271387 177246
rect -960 175796 480 176036
rect 46657 174586 46723 174589
rect 281809 174586 281875 174589
rect 46657 174584 281875 174586
rect 46657 174528 46662 174584
rect 46718 174528 281814 174584
rect 281870 174528 281875 174584
rect 46657 174526 281875 174528
rect 46657 174523 46723 174526
rect 281809 174523 281875 174526
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 3417 162890 3483 162893
rect -960 162888 3483 162890
rect -960 162832 3422 162888
rect 3478 162832 3483 162888
rect -960 162830 3483 162832
rect -960 162740 480 162830
rect 3417 162827 3483 162830
rect 239622 152628 239628 152692
rect 239692 152690 239698 152692
rect 583520 152690 584960 152780
rect 239692 152630 584960 152690
rect 239692 152628 239698 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 288382 149834 288388 149836
rect -960 149774 288388 149834
rect -960 149684 480 149774
rect 288382 149772 288388 149774
rect 288452 149772 288458 149836
rect 346894 139300 346900 139364
rect 346964 139362 346970 139364
rect 583520 139362 584960 139452
rect 346964 139302 584960 139362
rect 346964 139300 346970 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 235206 136778 235212 136780
rect -960 136718 235212 136778
rect -960 136628 480 136718
rect 235206 136716 235212 136718
rect 235276 136716 235282 136780
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 239806 112780 239812 112844
rect 239876 112842 239882 112844
rect 583520 112842 584960 112932
rect 239876 112782 584960 112842
rect 239876 112780 239882 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 45461 106858 45527 106861
rect 184197 106858 184263 106861
rect 45461 106856 184263 106858
rect 45461 106800 45466 106856
rect 45522 106800 184202 106856
rect 184258 106800 184263 106856
rect 45461 106798 184263 106800
rect 45461 106795 45527 106798
rect 184197 106795 184263 106798
rect 41873 105498 41939 105501
rect 191097 105498 191163 105501
rect 41873 105496 191163 105498
rect 41873 105440 41878 105496
rect 41934 105440 191102 105496
rect 191158 105440 191163 105496
rect 41873 105438 191163 105440
rect 41873 105435 41939 105438
rect 191097 105435 191163 105438
rect 38377 104138 38443 104141
rect 197997 104138 198063 104141
rect 38377 104136 198063 104138
rect 38377 104080 38382 104136
rect 38438 104080 198002 104136
rect 198058 104080 198063 104136
rect 38377 104078 198063 104080
rect 38377 104075 38443 104078
rect 197997 104075 198063 104078
rect 27705 102778 27771 102781
rect 209037 102778 209103 102781
rect 27705 102776 209103 102778
rect 27705 102720 27710 102776
rect 27766 102720 209042 102776
rect 209098 102720 209103 102776
rect 27705 102718 209103 102720
rect 27705 102715 27771 102718
rect 209037 102715 209103 102718
rect 112805 101418 112871 101421
rect 199377 101418 199443 101421
rect 112805 101416 199443 101418
rect 112805 101360 112810 101416
rect 112866 101360 199382 101416
rect 199438 101360 199443 101416
rect 112805 101358 199443 101360
rect 112805 101355 112871 101358
rect 199377 101355 199443 101358
rect 102225 100058 102291 100061
rect 217317 100058 217383 100061
rect 102225 100056 217383 100058
rect 102225 100000 102230 100056
rect 102286 100000 217322 100056
rect 217378 100000 217383 100056
rect 102225 99998 217383 100000
rect 102225 99995 102291 99998
rect 217317 99995 217383 99998
rect 500166 99452 500172 99516
rect 500236 99514 500242 99516
rect 583520 99514 584960 99604
rect 500236 99454 584960 99514
rect 500236 99452 500242 99454
rect 583520 99364 584960 99454
rect 95141 98698 95207 98701
rect 174537 98698 174603 98701
rect 95141 98696 174603 98698
rect 95141 98640 95146 98696
rect 95202 98640 174542 98696
rect 174598 98640 174603 98696
rect 95141 98638 174603 98640
rect 95141 98635 95207 98638
rect 174537 98635 174603 98638
rect -960 97610 480 97700
rect 287094 97610 287100 97612
rect -960 97550 287100 97610
rect -960 97460 480 97550
rect 287094 97548 287100 97550
rect 287164 97548 287170 97612
rect 91553 97202 91619 97205
rect 211797 97202 211863 97205
rect 91553 97200 211863 97202
rect 91553 97144 91558 97200
rect 91614 97144 211802 97200
rect 211858 97144 211863 97200
rect 91553 97142 211863 97144
rect 91553 97139 91619 97142
rect 211797 97139 211863 97142
rect 8753 95842 8819 95845
rect 226977 95842 227043 95845
rect 8753 95840 227043 95842
rect 8753 95784 8758 95840
rect 8814 95784 226982 95840
rect 227038 95784 227043 95840
rect 8753 95782 227043 95784
rect 8753 95779 8819 95782
rect 226977 95779 227043 95782
rect 4061 94482 4127 94485
rect 210417 94482 210483 94485
rect 4061 94480 210483 94482
rect 4061 94424 4066 94480
rect 4122 94424 210422 94480
rect 210478 94424 210483 94480
rect 4061 94422 210483 94424
rect 4061 94419 4127 94422
rect 210417 94419 210483 94422
rect 111609 93122 111675 93125
rect 274909 93122 274975 93125
rect 111609 93120 274975 93122
rect 111609 93064 111614 93120
rect 111670 93064 274914 93120
rect 274970 93064 274975 93120
rect 111609 93062 274975 93064
rect 111609 93059 111675 93062
rect 274909 93059 274975 93062
rect 86861 91762 86927 91765
rect 266537 91762 266603 91765
rect 86861 91760 266603 91762
rect 86861 91704 86866 91760
rect 86922 91704 266542 91760
rect 266598 91704 266603 91760
rect 86861 91702 266603 91704
rect 86861 91699 86927 91702
rect 266537 91699 266603 91702
rect 87597 90402 87663 90405
rect 214557 90402 214623 90405
rect 87597 90400 214623 90402
rect 87597 90344 87602 90400
rect 87658 90344 214562 90400
rect 214618 90344 214623 90400
rect 87597 90342 214623 90344
rect 87597 90339 87663 90342
rect 214557 90339 214623 90342
rect 89161 89042 89227 89045
rect 285673 89042 285739 89045
rect 89161 89040 285739 89042
rect 89161 88984 89166 89040
rect 89222 88984 285678 89040
rect 285734 88984 285739 89040
rect 89161 88982 285739 88984
rect 89161 88979 89227 88982
rect 285673 88979 285739 88982
rect 52913 87818 52979 87821
rect 86217 87818 86283 87821
rect 52913 87816 86283 87818
rect 52913 87760 52918 87816
rect 52974 87760 86222 87816
rect 86278 87760 86283 87816
rect 52913 87758 86283 87760
rect 52913 87755 52979 87758
rect 86217 87755 86283 87758
rect 63861 87682 63927 87685
rect 87873 87682 87939 87685
rect 63861 87680 87939 87682
rect 63861 87624 63866 87680
rect 63922 87624 87878 87680
rect 87934 87624 87939 87680
rect 63861 87622 87939 87624
rect 63861 87619 63927 87622
rect 87873 87619 87939 87622
rect 59261 87546 59327 87549
rect 84929 87546 84995 87549
rect 59261 87544 84995 87546
rect 59261 87488 59266 87544
rect 59322 87488 84934 87544
rect 84990 87488 84995 87544
rect 59261 87486 84995 87488
rect 59261 87483 59327 87486
rect 84929 87483 84995 87486
rect 62021 87410 62087 87413
rect 90633 87410 90699 87413
rect 62021 87408 90699 87410
rect 62021 87352 62026 87408
rect 62082 87352 90638 87408
rect 90694 87352 90699 87408
rect 62021 87350 90699 87352
rect 62021 87347 62087 87350
rect 90633 87347 90699 87350
rect 57605 87274 57671 87277
rect 86401 87274 86467 87277
rect 57605 87272 86467 87274
rect 57605 87216 57610 87272
rect 57666 87216 86406 87272
rect 86462 87216 86467 87272
rect 57605 87214 86467 87216
rect 57605 87211 57671 87214
rect 86401 87211 86467 87214
rect 54661 87138 54727 87141
rect 87689 87138 87755 87141
rect 54661 87136 87755 87138
rect 54661 87080 54666 87136
rect 54722 87080 87694 87136
rect 87750 87080 87755 87136
rect 54661 87078 87755 87080
rect 54661 87075 54727 87078
rect 87689 87075 87755 87078
rect 65609 87002 65675 87005
rect 90449 87002 90515 87005
rect 65609 87000 90515 87002
rect 65609 86944 65614 87000
rect 65670 86944 90454 87000
rect 90510 86944 90515 87000
rect 65609 86942 90515 86944
rect 65609 86939 65675 86942
rect 90449 86939 90515 86942
rect 3182 86260 3188 86324
rect 3252 86322 3258 86324
rect 230974 86322 230980 86324
rect 3252 86262 230980 86322
rect 3252 86260 3258 86262
rect 230974 86260 230980 86262
rect 231044 86260 231050 86324
rect 56501 86186 56567 86189
rect 311433 86186 311499 86189
rect 56501 86184 311499 86186
rect 56501 86128 56506 86184
rect 56562 86128 311438 86184
rect 311494 86128 311499 86184
rect 56501 86126 311499 86128
rect 56501 86123 56567 86126
rect 311433 86123 311499 86126
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 68645 86050 68711 86053
rect 275277 86050 275343 86053
rect 68645 86048 275343 86050
rect 68645 85992 68650 86048
rect 68706 85992 275282 86048
rect 275338 85992 275343 86048
rect 583520 86036 584960 86126
rect 68645 85990 275343 85992
rect 68645 85987 68711 85990
rect 275277 85987 275343 85990
rect 50981 85914 51047 85917
rect 271137 85914 271203 85917
rect 50981 85912 271203 85914
rect 50981 85856 50986 85912
rect 51042 85856 271142 85912
rect 271198 85856 271203 85912
rect 50981 85854 271203 85856
rect 50981 85851 51047 85854
rect 271137 85851 271203 85854
rect 60641 85778 60707 85781
rect 322105 85778 322171 85781
rect 60641 85776 322171 85778
rect 60641 85720 60646 85776
rect 60702 85720 322110 85776
rect 322166 85720 322171 85776
rect 60641 85718 322171 85720
rect 60641 85715 60707 85718
rect 322105 85715 322171 85718
rect 66989 85642 67055 85645
rect 336273 85642 336339 85645
rect 66989 85640 336339 85642
rect 66989 85584 66994 85640
rect 67050 85584 336278 85640
rect 336334 85584 336339 85640
rect 66989 85582 336339 85584
rect 66989 85579 67055 85582
rect 336273 85579 336339 85582
rect 82307 84962 82373 84965
rect 368197 84962 368263 84965
rect 82307 84960 368263 84962
rect 82307 84904 82312 84960
rect 82368 84904 368202 84960
rect 368258 84904 368263 84960
rect 82307 84902 368263 84904
rect 82307 84899 82373 84902
rect 368197 84899 368263 84902
rect 77615 84826 77681 84829
rect 357525 84826 357591 84829
rect 77615 84824 357591 84826
rect -960 84690 480 84780
rect 77615 84768 77620 84824
rect 77676 84768 357530 84824
rect 357586 84768 357591 84824
rect 77615 84766 357591 84768
rect 77615 84763 77681 84766
rect 357525 84763 357591 84766
rect 3182 84690 3188 84692
rect -960 84630 3188 84690
rect -960 84540 480 84630
rect 3182 84628 3188 84630
rect 3252 84628 3258 84692
rect 71359 84690 71425 84693
rect 343357 84690 343423 84693
rect 71359 84688 343423 84690
rect 71359 84632 71364 84688
rect 71420 84632 343362 84688
rect 343418 84632 343423 84688
rect 71359 84630 343423 84632
rect 71359 84627 71425 84630
rect 343357 84627 343423 84630
rect 79179 84554 79245 84557
rect 361113 84554 361179 84557
rect 79179 84552 361179 84554
rect 79179 84496 79184 84552
rect 79240 84496 361118 84552
rect 361174 84496 361179 84552
rect 79179 84494 361179 84496
rect 79179 84491 79245 84494
rect 361113 84491 361179 84494
rect 84285 83466 84351 83469
rect 284937 83466 285003 83469
rect 84285 83464 285003 83466
rect 84285 83408 84290 83464
rect 84346 83408 284942 83464
rect 284998 83408 285003 83464
rect 84285 83406 285003 83408
rect 84285 83403 84351 83406
rect 284937 83403 285003 83406
rect 435357 83058 435423 83061
rect 84916 83056 435423 83058
rect 84916 83000 435362 83056
rect 435418 83000 435423 83056
rect 84916 82998 435423 83000
rect 435357 82995 435423 82998
rect 48037 81698 48103 81701
rect 432597 81698 432663 81701
rect 48037 81696 50140 81698
rect 48037 81640 48042 81696
rect 48098 81640 50140 81696
rect 48037 81638 50140 81640
rect 84916 81696 432663 81698
rect 84916 81640 432602 81696
rect 432658 81640 432663 81696
rect 84916 81638 432663 81640
rect 48037 81635 48103 81638
rect 432597 81635 432663 81638
rect 84929 80746 84995 80749
rect 318517 80746 318583 80749
rect 84929 80744 318583 80746
rect 84929 80688 84934 80744
rect 84990 80688 318522 80744
rect 318578 80688 318583 80744
rect 84929 80686 318583 80688
rect 84929 80683 84995 80686
rect 318517 80683 318583 80686
rect 48129 80338 48195 80341
rect 428549 80338 428615 80341
rect 48129 80336 50140 80338
rect 48129 80280 48134 80336
rect 48190 80280 50140 80336
rect 48129 80278 50140 80280
rect 84916 80336 428615 80338
rect 84916 80280 428554 80336
rect 428610 80280 428615 80336
rect 84916 80278 428615 80280
rect 48129 80275 48195 80278
rect 428549 80275 428615 80278
rect 49325 78978 49391 78981
rect 250437 78978 250503 78981
rect 49325 78976 50140 78978
rect 49325 78920 49330 78976
rect 49386 78920 50140 78976
rect 49325 78918 50140 78920
rect 84916 78976 250503 78978
rect 84916 78920 250442 78976
rect 250498 78920 250503 78976
rect 84916 78918 250503 78920
rect 49325 78915 49391 78918
rect 250437 78915 250503 78918
rect 49601 77618 49667 77621
rect 421557 77618 421623 77621
rect 49601 77616 50140 77618
rect 49601 77560 49606 77616
rect 49662 77560 50140 77616
rect 49601 77558 50140 77560
rect 84916 77616 421623 77618
rect 84916 77560 421562 77616
rect 421618 77560 421623 77616
rect 84916 77558 421623 77560
rect 49601 77555 49667 77558
rect 421557 77555 421623 77558
rect 417417 76258 417483 76261
rect 84916 76256 417483 76258
rect 50294 75989 50354 76228
rect 84916 76200 417422 76256
rect 417478 76200 417483 76256
rect 84916 76198 417483 76200
rect 417417 76195 417483 76198
rect 50245 75984 50354 75989
rect 50245 75928 50250 75984
rect 50306 75928 50354 75984
rect 50245 75926 50354 75928
rect 50245 75923 50311 75926
rect 49509 74898 49575 74901
rect 414657 74898 414723 74901
rect 49509 74896 50140 74898
rect 49509 74840 49514 74896
rect 49570 74840 50140 74896
rect 49509 74838 50140 74840
rect 84916 74896 414723 74898
rect 84916 74840 414662 74896
rect 414718 74840 414723 74896
rect 84916 74838 414723 74840
rect 49509 74835 49575 74838
rect 414657 74835 414723 74838
rect 450537 73538 450603 73541
rect 84916 73536 450603 73538
rect 50478 73269 50538 73508
rect 84916 73480 450542 73536
rect 450598 73480 450603 73536
rect 84916 73478 450603 73480
rect 450537 73475 450603 73478
rect 50429 73264 50538 73269
rect 50429 73208 50434 73264
rect 50490 73208 50538 73264
rect 50429 73206 50538 73208
rect 50429 73203 50495 73206
rect 580349 72994 580415 72997
rect 583520 72994 584960 73084
rect 580349 72992 584960 72994
rect 580349 72936 580354 72992
rect 580410 72936 584960 72992
rect 580349 72934 584960 72936
rect 580349 72931 580415 72934
rect 583520 72844 584960 72934
rect 49417 72178 49483 72181
rect 447777 72178 447843 72181
rect 49417 72176 50140 72178
rect 49417 72120 49422 72176
rect 49478 72120 50140 72176
rect 49417 72118 50140 72120
rect 84916 72176 447843 72178
rect 84916 72120 447782 72176
rect 447838 72120 447843 72176
rect 84916 72118 447843 72120
rect 49417 72115 49483 72118
rect 447777 72115 447843 72118
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 443637 70818 443703 70821
rect 84916 70816 443703 70818
rect 50110 70413 50170 70788
rect 84916 70760 443642 70816
rect 443698 70760 443703 70816
rect 84916 70758 443703 70760
rect 443637 70755 443703 70758
rect 50110 70408 50219 70413
rect 50110 70352 50158 70408
rect 50214 70352 50219 70408
rect 50110 70350 50219 70352
rect 50153 70347 50219 70350
rect 90633 69594 90699 69597
rect 325601 69594 325667 69597
rect 90633 69592 325667 69594
rect 90633 69536 90638 69592
rect 90694 69536 325606 69592
rect 325662 69536 325667 69592
rect 90633 69534 325667 69536
rect 90633 69531 90699 69534
rect 325601 69531 325667 69534
rect 49233 69458 49299 69461
rect 246297 69458 246363 69461
rect 49233 69456 50140 69458
rect 49233 69400 49238 69456
rect 49294 69400 50140 69456
rect 49233 69398 50140 69400
rect 84916 69456 246363 69458
rect 84916 69400 246302 69456
rect 246358 69400 246363 69456
rect 84916 69398 246363 69400
rect 49233 69395 49299 69398
rect 246297 69395 246363 69398
rect 49049 68098 49115 68101
rect 431217 68098 431283 68101
rect 49049 68096 50140 68098
rect 49049 68040 49054 68096
rect 49110 68040 50140 68096
rect 49049 68038 50140 68040
rect 84916 68096 431283 68098
rect 84916 68040 431222 68096
rect 431278 68040 431283 68096
rect 84916 68038 431283 68040
rect 49049 68035 49115 68038
rect 431217 68035 431283 68038
rect 436737 66738 436803 66741
rect 84916 66736 436803 66738
rect 50294 66333 50354 66708
rect 84916 66680 436742 66736
rect 436798 66680 436803 66736
rect 84916 66678 436803 66680
rect 436737 66675 436803 66678
rect 50294 66328 50403 66333
rect 50294 66272 50342 66328
rect 50398 66272 50403 66328
rect 50294 66270 50403 66272
rect 50337 66267 50403 66270
rect 429837 65378 429903 65381
rect 84916 65376 429903 65378
rect 50478 65106 50538 65348
rect 84916 65320 429842 65376
rect 429898 65320 429903 65376
rect 84916 65318 429903 65320
rect 429837 65315 429903 65318
rect 50613 65106 50679 65109
rect 50478 65104 50679 65106
rect 50478 65048 50618 65104
rect 50674 65048 50679 65104
rect 50478 65046 50679 65048
rect 50613 65043 50679 65046
rect 47577 64018 47643 64021
rect 406377 64018 406443 64021
rect 47577 64016 50140 64018
rect 47577 63960 47582 64016
rect 47638 63960 50140 64016
rect 47577 63958 50140 63960
rect 84916 64016 406443 64018
rect 84916 63960 406382 64016
rect 406438 63960 406443 64016
rect 84916 63958 406443 63960
rect 47577 63955 47643 63958
rect 406377 63955 406443 63958
rect 47945 62658 48011 62661
rect 425697 62658 425763 62661
rect 47945 62656 50140 62658
rect 47945 62600 47950 62656
rect 48006 62600 50140 62656
rect 47945 62598 50140 62600
rect 84916 62656 425763 62658
rect 84916 62600 425702 62656
rect 425758 62600 425763 62656
rect 84916 62598 425763 62600
rect 47945 62595 48011 62598
rect 425697 62595 425763 62598
rect 47853 61298 47919 61301
rect 422937 61298 423003 61301
rect 47853 61296 50140 61298
rect 47853 61240 47858 61296
rect 47914 61240 50140 61296
rect 47853 61238 50140 61240
rect 84916 61296 423003 61298
rect 84916 61240 422942 61296
rect 422998 61240 423003 61296
rect 84916 61238 423003 61240
rect 47853 61235 47919 61238
rect 422937 61235 423003 61238
rect 47761 59938 47827 59941
rect 418797 59938 418863 59941
rect 47761 59936 50140 59938
rect 47761 59880 47766 59936
rect 47822 59880 50140 59936
rect 47761 59878 50140 59880
rect 84916 59936 418863 59938
rect 84916 59880 418802 59936
rect 418858 59880 418863 59936
rect 84916 59878 418863 59880
rect 47761 59875 47827 59878
rect 418797 59875 418863 59878
rect 559414 59604 559420 59668
rect 559484 59666 559490 59668
rect 583520 59666 584960 59756
rect 559484 59606 584960 59666
rect 559484 59604 559490 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3550 58578 3556 58580
rect -960 58518 3556 58578
rect -960 58428 480 58518
rect 3550 58516 3556 58518
rect 3620 58516 3626 58580
rect 47669 58578 47735 58581
rect 411897 58578 411963 58581
rect 47669 58576 50140 58578
rect 47669 58520 47674 58576
rect 47730 58520 50140 58576
rect 47669 58518 50140 58520
rect 84916 58576 411963 58578
rect 84916 58520 411902 58576
rect 411958 58520 411963 58576
rect 84916 58518 411963 58520
rect 47669 58515 47735 58518
rect 411897 58515 411963 58518
rect 47485 57218 47551 57221
rect 353937 57218 354003 57221
rect 47485 57216 50140 57218
rect 47485 57160 47490 57216
rect 47546 57160 50140 57216
rect 47485 57158 50140 57160
rect 84916 57216 354003 57218
rect 84916 57160 353942 57216
rect 353998 57160 354003 57216
rect 84916 57158 354003 57160
rect 47485 57155 47551 57158
rect 353937 57155 354003 57158
rect 351177 55858 351243 55861
rect 84916 55856 351243 55858
rect 50478 55589 50538 55828
rect 84916 55800 351182 55856
rect 351238 55800 351243 55856
rect 84916 55798 351243 55800
rect 351177 55795 351243 55798
rect 50478 55584 50587 55589
rect 50478 55528 50526 55584
rect 50582 55528 50587 55584
rect 50478 55526 50587 55528
rect 50521 55523 50587 55526
rect 87873 54634 87939 54637
rect 329189 54634 329255 54637
rect 87873 54632 329255 54634
rect 87873 54576 87878 54632
rect 87934 54576 329194 54632
rect 329250 54576 329255 54632
rect 87873 54574 329255 54576
rect 87873 54571 87939 54574
rect 329189 54571 329255 54574
rect 49141 54498 49207 54501
rect 273897 54498 273963 54501
rect 49141 54496 50140 54498
rect 49141 54440 49146 54496
rect 49202 54440 50140 54496
rect 49141 54438 50140 54440
rect 84916 54496 273963 54498
rect 84916 54440 273902 54496
rect 273958 54440 273963 54496
rect 84916 54438 273963 54440
rect 49141 54435 49207 54438
rect 273897 54435 273963 54438
rect 84653 53274 84719 53277
rect 213177 53274 213243 53277
rect 84653 53272 213243 53274
rect 84653 53216 84658 53272
rect 84714 53216 213182 53272
rect 213238 53216 213243 53272
rect 84653 53214 213243 53216
rect 84653 53211 84719 53214
rect 213177 53211 213243 53214
rect 86401 53138 86467 53141
rect 315021 53138 315087 53141
rect 86401 53136 315087 53138
rect 50110 52597 50170 53108
rect 86401 53080 86406 53136
rect 86462 53080 315026 53136
rect 315082 53080 315087 53136
rect 86401 53078 315087 53080
rect 86401 53075 86467 53078
rect 315021 53075 315087 53078
rect 50061 52592 50170 52597
rect 50061 52536 50066 52592
rect 50122 52536 50170 52592
rect 50061 52534 50170 52536
rect 84886 52594 84946 53040
rect 86953 52594 87019 52597
rect 87597 52594 87663 52597
rect 84886 52592 87663 52594
rect 84886 52536 86958 52592
rect 87014 52536 87602 52592
rect 87658 52536 87663 52592
rect 84886 52534 87663 52536
rect 50061 52531 50127 52534
rect 86953 52531 87019 52534
rect 87597 52531 87663 52534
rect 565 51778 631 51781
rect 86217 51778 86283 51781
rect 304349 51778 304415 51781
rect 565 51776 45570 51778
rect 565 51720 570 51776
rect 626 51720 45570 51776
rect 86217 51776 304415 51778
rect 565 51718 45570 51720
rect 565 51715 631 51718
rect 45510 51506 45570 51718
rect 48221 51506 48287 51509
rect 45510 51504 64890 51506
rect 45510 51448 48226 51504
rect 48282 51448 64890 51504
rect 45510 51446 64890 51448
rect 48221 51443 48287 51446
rect 64830 51370 64890 51446
rect 84334 51370 84394 51748
rect 86217 51720 86222 51776
rect 86278 51720 304354 51776
rect 304410 51720 304415 51776
rect 86217 51718 304415 51720
rect 86217 51715 86283 51718
rect 304349 51715 304415 51718
rect 64830 51310 84394 51370
rect 83273 50554 83339 50557
rect 265249 50554 265315 50557
rect 83273 50552 265315 50554
rect 83273 50496 83278 50552
rect 83334 50496 265254 50552
rect 265310 50496 265315 50552
rect 83273 50494 265315 50496
rect 83273 50491 83339 50494
rect 265249 50491 265315 50494
rect 250437 50418 250503 50421
rect 467465 50418 467531 50421
rect 250437 50416 467531 50418
rect 250437 50360 250442 50416
rect 250498 50360 467470 50416
rect 467526 50360 467531 50416
rect 250437 50358 467531 50360
rect 250437 50355 250503 50358
rect 467465 50355 467531 50358
rect 87689 50282 87755 50285
rect 307937 50282 308003 50285
rect 87689 50280 308003 50282
rect 87689 50224 87694 50280
rect 87750 50224 307942 50280
rect 307998 50224 308003 50280
rect 87689 50222 308003 50224
rect 87689 50219 87755 50222
rect 307937 50219 308003 50222
rect 48129 49058 48195 49061
rect 268837 49058 268903 49061
rect 48129 49056 268903 49058
rect 48129 49000 48134 49056
rect 48190 49000 268842 49056
rect 268898 49000 268903 49056
rect 48129 48998 268903 49000
rect 48129 48995 48195 48998
rect 268837 48995 268903 48998
rect 49049 48922 49115 48925
rect 520733 48922 520799 48925
rect 49049 48920 520799 48922
rect 49049 48864 49054 48920
rect 49110 48864 520738 48920
rect 520794 48864 520799 48920
rect 49049 48862 520799 48864
rect 49049 48859 49115 48862
rect 520733 48859 520799 48862
rect 82721 47970 82787 47973
rect 83457 47970 83523 47973
rect 82721 47968 83523 47970
rect 82721 47912 82726 47968
rect 82782 47912 83462 47968
rect 83518 47912 83523 47968
rect 82721 47910 83523 47912
rect 82721 47907 82787 47910
rect 83457 47907 83523 47910
rect 50981 47834 51047 47837
rect 439497 47834 439563 47837
rect 50981 47832 439563 47834
rect 50981 47776 50986 47832
rect 51042 47776 439502 47832
rect 439558 47776 439563 47832
rect 50981 47774 439563 47776
rect 50981 47771 51047 47774
rect 439497 47771 439563 47774
rect 52361 47698 52427 47701
rect 442257 47698 442323 47701
rect 52361 47696 442323 47698
rect 52361 47640 52366 47696
rect 52422 47640 442262 47696
rect 442318 47640 442323 47696
rect 52361 47638 442323 47640
rect 52361 47635 52427 47638
rect 442257 47635 442323 47638
rect 53741 47562 53807 47565
rect 446397 47562 446463 47565
rect 53741 47560 446463 47562
rect 53741 47504 53746 47560
rect 53802 47504 446402 47560
rect 446458 47504 446463 47560
rect 53741 47502 446463 47504
rect 53741 47499 53807 47502
rect 446397 47499 446463 47502
rect 74441 47018 74507 47021
rect 75177 47018 75243 47021
rect 74441 47016 75243 47018
rect 74441 46960 74446 47016
rect 74502 46960 75182 47016
rect 75238 46960 75243 47016
rect 74441 46958 75243 46960
rect 74441 46955 74507 46958
rect 75177 46955 75243 46958
rect 50613 46338 50679 46341
rect 293677 46338 293743 46341
rect 50613 46336 293743 46338
rect 50613 46280 50618 46336
rect 50674 46280 293682 46336
rect 293738 46280 293743 46336
rect 50613 46278 293743 46280
rect 50613 46275 50679 46278
rect 293677 46275 293743 46278
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 56501 46202 56567 46205
rect 481725 46202 481791 46205
rect 56501 46200 481791 46202
rect 56501 46144 56506 46200
rect 56562 46144 481730 46200
rect 481786 46144 481791 46200
rect 583520 46188 584960 46278
rect 56501 46142 481791 46144
rect 56501 46139 56567 46142
rect 481725 46139 481791 46142
rect -960 45522 480 45612
rect 224166 45522 224172 45524
rect -960 45462 224172 45522
rect -960 45372 480 45462
rect 224166 45460 224172 45462
rect 224236 45460 224242 45524
rect 49325 44842 49391 44845
rect 549069 44842 549135 44845
rect 49325 44840 549135 44842
rect 49325 44784 49330 44840
rect 49386 44784 549074 44840
rect 549130 44784 549135 44840
rect 49325 44782 549135 44784
rect 49325 44779 49391 44782
rect 549069 44779 549135 44782
rect 50061 43618 50127 43621
rect 297265 43618 297331 43621
rect 50061 43616 297331 43618
rect 50061 43560 50066 43616
rect 50122 43560 297270 43616
rect 297326 43560 297331 43616
rect 50061 43558 297331 43560
rect 50061 43555 50127 43558
rect 297265 43555 297331 43558
rect 64689 43482 64755 43485
rect 502977 43482 503043 43485
rect 64689 43480 503043 43482
rect 64689 43424 64694 43480
rect 64750 43424 502982 43480
rect 503038 43424 503043 43480
rect 64689 43422 503043 43424
rect 64689 43419 64755 43422
rect 502977 43419 503043 43422
rect 48037 42258 48103 42261
rect 300761 42258 300827 42261
rect 48037 42256 300827 42258
rect 48037 42200 48042 42256
rect 48098 42200 300766 42256
rect 300822 42200 300827 42256
rect 48037 42198 300827 42200
rect 48037 42195 48103 42198
rect 300761 42195 300827 42198
rect 67449 42122 67515 42125
rect 508497 42122 508563 42125
rect 67449 42120 508563 42122
rect 67449 42064 67454 42120
rect 67510 42064 508502 42120
rect 508558 42064 508563 42120
rect 67449 42062 508563 42064
rect 67449 42059 67515 42062
rect 508497 42059 508563 42062
rect 7557 40898 7623 40901
rect 86953 40898 87019 40901
rect 7557 40896 87019 40898
rect 7557 40840 7562 40896
rect 7618 40840 86958 40896
rect 87014 40840 87019 40896
rect 7557 40838 87019 40840
rect 7557 40835 7623 40838
rect 86953 40835 87019 40838
rect 81249 40762 81315 40765
rect 400121 40762 400187 40765
rect 81249 40760 400187 40762
rect 81249 40704 81254 40760
rect 81310 40704 400126 40760
rect 400182 40704 400187 40760
rect 81249 40702 400187 40704
rect 81249 40699 81315 40702
rect 400121 40699 400187 40702
rect 68829 40626 68895 40629
rect 512637 40626 512703 40629
rect 68829 40624 512703 40626
rect 68829 40568 68834 40624
rect 68890 40568 512642 40624
rect 512698 40568 512703 40624
rect 68829 40566 512703 40568
rect 68829 40563 68895 40566
rect 512637 40563 512703 40566
rect 84009 39402 84075 39405
rect 407205 39402 407271 39405
rect 84009 39400 407271 39402
rect 84009 39344 84014 39400
rect 84070 39344 407210 39400
rect 407266 39344 407271 39400
rect 84009 39342 407271 39344
rect 84009 39339 84075 39342
rect 407205 39339 407271 39342
rect 49233 39266 49299 39269
rect 524229 39266 524295 39269
rect 49233 39264 524295 39266
rect 49233 39208 49238 39264
rect 49294 39208 524234 39264
rect 524290 39208 524295 39264
rect 49233 39206 524295 39208
rect 49233 39203 49299 39206
rect 524229 39203 524295 39206
rect 51349 38042 51415 38045
rect 254577 38042 254643 38045
rect 51349 38040 254643 38042
rect 51349 37984 51354 38040
rect 51410 37984 254582 38040
rect 254638 37984 254643 38040
rect 51349 37982 254643 37984
rect 51349 37979 51415 37982
rect 254577 37979 254643 37982
rect 49417 37906 49483 37909
rect 531313 37906 531379 37909
rect 49417 37904 531379 37906
rect 49417 37848 49422 37904
rect 49478 37848 531318 37904
rect 531374 37848 531379 37904
rect 49417 37846 531379 37848
rect 49417 37843 49483 37846
rect 531313 37843 531379 37846
rect 77385 36818 77451 36821
rect 195237 36818 195303 36821
rect 77385 36816 195303 36818
rect 77385 36760 77390 36816
rect 77446 36760 195242 36816
rect 195298 36760 195303 36816
rect 77385 36758 195303 36760
rect 77385 36755 77451 36758
rect 195237 36755 195303 36758
rect 51717 36682 51783 36685
rect 282545 36682 282611 36685
rect 51717 36680 282611 36682
rect 51717 36624 51722 36680
rect 51778 36624 282550 36680
rect 282606 36624 282611 36680
rect 51717 36622 282611 36624
rect 51717 36619 51783 36622
rect 282545 36619 282611 36622
rect 50429 36546 50495 36549
rect 534901 36546 534967 36549
rect 50429 36544 534967 36546
rect 50429 36488 50434 36544
rect 50490 36488 534906 36544
rect 534962 36488 534967 36544
rect 50429 36486 534967 36488
rect 50429 36483 50495 36486
rect 534901 36483 534967 36486
rect 73797 35322 73863 35325
rect 220077 35322 220143 35325
rect 73797 35320 220143 35322
rect 73797 35264 73802 35320
rect 73858 35264 220082 35320
rect 220138 35264 220143 35320
rect 73797 35262 220143 35264
rect 73797 35259 73863 35262
rect 220077 35259 220143 35262
rect 49509 35186 49575 35189
rect 538397 35186 538463 35189
rect 49509 35184 538463 35186
rect 49509 35128 49514 35184
rect 49570 35128 538402 35184
rect 538458 35128 538463 35184
rect 49509 35126 538463 35128
rect 49509 35123 49575 35126
rect 538397 35123 538463 35126
rect 70301 34098 70367 34101
rect 142797 34098 142863 34101
rect 70301 34096 142863 34098
rect 70301 34040 70306 34096
rect 70362 34040 142802 34096
rect 142858 34040 142863 34096
rect 70301 34038 142863 34040
rect 70301 34035 70367 34038
rect 142797 34035 142863 34038
rect 80881 33962 80947 33965
rect 228357 33962 228423 33965
rect 80881 33960 228423 33962
rect 80881 33904 80886 33960
rect 80942 33904 228362 33960
rect 228418 33904 228423 33960
rect 80881 33902 228423 33904
rect 80881 33899 80947 33902
rect 228357 33899 228423 33902
rect 50245 33826 50311 33829
rect 541985 33826 542051 33829
rect 50245 33824 542051 33826
rect 50245 33768 50250 33824
rect 50306 33768 541990 33824
rect 542046 33768 542051 33824
rect 50245 33766 542051 33768
rect 50245 33763 50311 33766
rect 541985 33763 542051 33766
rect 580257 33146 580323 33149
rect 583520 33146 584960 33236
rect 580257 33144 584960 33146
rect 580257 33088 580262 33144
rect 580318 33088 584960 33144
rect 580257 33086 584960 33088
rect 580257 33083 580323 33086
rect 583520 32996 584960 33086
rect 66713 32738 66779 32741
rect 175917 32738 175983 32741
rect 66713 32736 175983 32738
rect 66713 32680 66718 32736
rect 66774 32680 175922 32736
rect 175978 32680 175983 32736
rect 66713 32678 175983 32680
rect 66713 32675 66779 32678
rect 175917 32675 175983 32678
rect 71497 32602 71563 32605
rect 280654 32602 280660 32604
rect 71497 32600 280660 32602
rect -960 32466 480 32556
rect 71497 32544 71502 32600
rect 71558 32544 280660 32600
rect 71497 32542 280660 32544
rect 71497 32539 71563 32542
rect 280654 32540 280660 32542
rect 280724 32540 280730 32604
rect 3417 32466 3483 32469
rect -960 32464 3483 32466
rect -960 32408 3422 32464
rect 3478 32408 3483 32464
rect -960 32406 3483 32408
rect -960 32316 480 32406
rect 3417 32403 3483 32406
rect 49601 32466 49667 32469
rect 545481 32466 545547 32469
rect 49601 32464 545547 32466
rect 49601 32408 49606 32464
rect 49662 32408 545486 32464
rect 545542 32408 545547 32464
rect 49601 32406 545547 32408
rect 49601 32403 49667 32406
rect 545481 32403 545547 32406
rect 63217 31106 63283 31109
rect 203517 31106 203583 31109
rect 63217 31104 203583 31106
rect 63217 31048 63222 31104
rect 63278 31048 203522 31104
rect 203578 31048 203583 31104
rect 63217 31046 203583 31048
rect 63217 31043 63283 31046
rect 203517 31043 203583 31046
rect 49141 30970 49207 30973
rect 552657 30970 552723 30973
rect 49141 30968 552723 30970
rect 49141 30912 49146 30968
rect 49202 30912 552662 30968
rect 552718 30912 552723 30968
rect 49141 30910 552723 30912
rect 49141 30907 49207 30910
rect 552657 30907 552723 30910
rect 56041 29882 56107 29885
rect 188337 29882 188403 29885
rect 56041 29880 188403 29882
rect 56041 29824 56046 29880
rect 56102 29824 188342 29880
rect 188398 29824 188403 29880
rect 56041 29822 188403 29824
rect 56041 29819 56107 29822
rect 188337 29819 188403 29822
rect 82077 29746 82143 29749
rect 285622 29746 285628 29748
rect 82077 29744 285628 29746
rect 82077 29688 82082 29744
rect 82138 29688 285628 29744
rect 82077 29686 285628 29688
rect 82077 29683 82143 29686
rect 285622 29684 285628 29686
rect 285692 29684 285698 29748
rect 50521 29610 50587 29613
rect 556153 29610 556219 29613
rect 50521 29608 556219 29610
rect 50521 29552 50526 29608
rect 50582 29552 556158 29608
rect 556214 29552 556219 29608
rect 50521 29550 556219 29552
rect 50521 29547 50587 29550
rect 556153 29547 556219 29550
rect 59629 28522 59695 28525
rect 178677 28522 178743 28525
rect 59629 28520 178743 28522
rect 59629 28464 59634 28520
rect 59690 28464 178682 28520
rect 178738 28464 178743 28520
rect 59629 28462 178743 28464
rect 59629 28459 59695 28462
rect 178677 28459 178743 28462
rect 74993 28386 75059 28389
rect 282913 28386 282979 28389
rect 74993 28384 282979 28386
rect 74993 28328 74998 28384
rect 75054 28328 282918 28384
rect 282974 28328 282979 28384
rect 74993 28326 282979 28328
rect 74993 28323 75059 28326
rect 282913 28323 282979 28326
rect 47669 28250 47735 28253
rect 562317 28250 562383 28253
rect 47669 28248 562383 28250
rect 47669 28192 47674 28248
rect 47730 28192 562322 28248
rect 562378 28192 562383 28248
rect 47669 28190 562383 28192
rect 47669 28187 47735 28190
rect 562317 28187 562383 28190
rect 52545 27162 52611 27165
rect 151077 27162 151143 27165
rect 52545 27160 151143 27162
rect 52545 27104 52550 27160
rect 52606 27104 151082 27160
rect 151138 27104 151143 27160
rect 52545 27102 151143 27104
rect 52545 27099 52611 27102
rect 151077 27099 151143 27102
rect 53741 27026 53807 27029
rect 284518 27026 284524 27028
rect 53741 27024 284524 27026
rect 53741 26968 53746 27024
rect 53802 26968 284524 27024
rect 53741 26966 284524 26968
rect 53741 26963 53807 26966
rect 284518 26964 284524 26966
rect 284588 26964 284594 27028
rect 47761 26890 47827 26893
rect 566825 26890 566891 26893
rect 47761 26888 566891 26890
rect 47761 26832 47766 26888
rect 47822 26832 566830 26888
rect 566886 26832 566891 26888
rect 47761 26830 566891 26832
rect 47761 26827 47827 26830
rect 566825 26827 566891 26830
rect 79685 25666 79751 25669
rect 264145 25666 264211 25669
rect 79685 25664 264211 25666
rect 79685 25608 79690 25664
rect 79746 25608 264150 25664
rect 264206 25608 264211 25664
rect 79685 25606 264211 25608
rect 79685 25603 79751 25606
rect 264145 25603 264211 25606
rect 50337 25530 50403 25533
rect 517145 25530 517211 25533
rect 50337 25528 517211 25530
rect 50337 25472 50342 25528
rect 50398 25472 517150 25528
rect 517206 25472 517211 25528
rect 50337 25470 517211 25472
rect 50337 25467 50403 25470
rect 517145 25467 517211 25470
rect 65517 24306 65583 24309
rect 259361 24306 259427 24309
rect 65517 24304 259427 24306
rect 65517 24248 65522 24304
rect 65578 24248 259366 24304
rect 259422 24248 259427 24304
rect 65517 24246 259427 24248
rect 65517 24243 65583 24246
rect 259361 24243 259427 24246
rect 47853 24170 47919 24173
rect 570321 24170 570387 24173
rect 47853 24168 570387 24170
rect 47853 24112 47858 24168
rect 47914 24112 570326 24168
rect 570382 24112 570387 24168
rect 47853 24110 570387 24112
rect 47853 24107 47919 24110
rect 570321 24107 570387 24110
rect 83457 22810 83523 22813
rect 403617 22810 403683 22813
rect 83457 22808 403683 22810
rect 83457 22752 83462 22808
rect 83518 22752 403622 22808
rect 403678 22752 403683 22808
rect 83457 22750 403683 22752
rect 83457 22747 83523 22750
rect 403617 22747 403683 22750
rect 47945 22674 48011 22677
rect 573909 22674 573975 22677
rect 47945 22672 573975 22674
rect 47945 22616 47950 22672
rect 48006 22616 573914 22672
rect 573970 22616 573975 22672
rect 47945 22614 573975 22616
rect 47945 22611 48011 22614
rect 573909 22611 573975 22614
rect 70209 21450 70275 21453
rect 278037 21450 278103 21453
rect 70209 21448 278103 21450
rect 70209 21392 70214 21448
rect 70270 21392 278042 21448
rect 278098 21392 278103 21448
rect 70209 21390 278103 21392
rect 70209 21387 70275 21390
rect 278037 21387 278103 21390
rect 72969 21314 73035 21317
rect 378869 21314 378935 21317
rect 72969 21312 378935 21314
rect 72969 21256 72974 21312
rect 73030 21256 378874 21312
rect 378930 21256 378935 21312
rect 72969 21254 378935 21256
rect 72969 21251 73035 21254
rect 378869 21251 378935 21254
rect 69105 20090 69171 20093
rect 260557 20090 260623 20093
rect 69105 20088 260623 20090
rect 69105 20032 69110 20088
rect 69166 20032 260562 20088
rect 260618 20032 260623 20088
rect 69105 20030 260623 20032
rect 69105 20027 69171 20030
rect 260557 20027 260623 20030
rect 47577 19954 47643 19957
rect 576117 19954 576183 19957
rect 47577 19952 576183 19954
rect 47577 19896 47582 19952
rect 47638 19896 576122 19952
rect 576178 19896 576183 19952
rect 47577 19894 576183 19896
rect 47577 19891 47643 19894
rect 576117 19891 576183 19894
rect 457294 19756 457300 19820
rect 457364 19818 457370 19820
rect 583520 19818 584960 19908
rect 457364 19758 584960 19818
rect 457364 19756 457370 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3366 19410 3372 19412
rect -960 19350 3372 19410
rect -960 19260 480 19350
rect 3366 19348 3372 19350
rect 3436 19348 3442 19412
rect 2865 18866 2931 18869
rect 159357 18866 159423 18869
rect 2865 18864 159423 18866
rect 2865 18808 2870 18864
rect 2926 18808 159362 18864
rect 159418 18808 159423 18864
rect 2865 18806 159423 18808
rect 2865 18803 2931 18806
rect 159357 18803 159423 18806
rect 64321 18730 64387 18733
rect 281533 18730 281599 18733
rect 64321 18728 281599 18730
rect 64321 18672 64326 18728
rect 64382 18672 281538 18728
rect 281594 18672 281599 18728
rect 64321 18670 281599 18672
rect 64321 18667 64387 18670
rect 281533 18667 281599 18670
rect 47485 18594 47551 18597
rect 559741 18594 559807 18597
rect 47485 18592 559807 18594
rect 47485 18536 47490 18592
rect 47546 18536 559746 18592
rect 559802 18536 559807 18592
rect 47485 18534 559807 18536
rect 47485 18531 47551 18534
rect 559741 18531 559807 18534
rect 79869 17370 79935 17373
rect 396533 17370 396599 17373
rect 79869 17368 396599 17370
rect 79869 17312 79874 17368
rect 79930 17312 396538 17368
rect 396594 17312 396599 17368
rect 79869 17310 396599 17312
rect 79869 17307 79935 17310
rect 396533 17307 396599 17310
rect 50153 17234 50219 17237
rect 527817 17234 527883 17237
rect 50153 17232 527883 17234
rect 50153 17176 50158 17232
rect 50214 17176 527822 17232
rect 527878 17176 527883 17232
rect 50153 17174 527883 17176
rect 50153 17171 50219 17174
rect 527817 17171 527883 17174
rect 79317 16010 79383 16013
rect 393037 16010 393103 16013
rect 79317 16008 393103 16010
rect 79317 15952 79322 16008
rect 79378 15952 393042 16008
rect 393098 15952 393103 16008
rect 79317 15950 393103 15952
rect 79317 15947 79383 15950
rect 393037 15947 393103 15950
rect 66069 15874 66135 15877
rect 506473 15874 506539 15877
rect 66069 15872 506539 15874
rect 66069 15816 66074 15872
rect 66130 15816 506478 15872
rect 506534 15816 506539 15872
rect 66069 15814 506539 15816
rect 66069 15811 66135 15814
rect 506473 15811 506539 15814
rect 77109 14650 77175 14653
rect 389449 14650 389515 14653
rect 77109 14648 389515 14650
rect 77109 14592 77114 14648
rect 77170 14592 389454 14648
rect 389510 14592 389515 14648
rect 77109 14590 389515 14592
rect 77109 14587 77175 14590
rect 389449 14587 389515 14590
rect 63309 14514 63375 14517
rect 499389 14514 499455 14517
rect 63309 14512 499455 14514
rect 63309 14456 63314 14512
rect 63370 14456 499394 14512
rect 499450 14456 499455 14512
rect 63309 14454 499455 14456
rect 63309 14451 63375 14454
rect 499389 14451 499455 14454
rect 76557 13154 76623 13157
rect 385953 13154 386019 13157
rect 76557 13152 386019 13154
rect 76557 13096 76562 13152
rect 76618 13096 385958 13152
rect 386014 13096 386019 13152
rect 76557 13094 386019 13096
rect 76557 13091 76623 13094
rect 385953 13091 386019 13094
rect 61929 13018 61995 13021
rect 495893 13018 495959 13021
rect 61929 13016 495959 13018
rect 61929 12960 61934 13016
rect 61990 12960 495898 13016
rect 495954 12960 495959 13016
rect 61929 12958 495959 12960
rect 61929 12955 61995 12958
rect 495893 12955 495959 12958
rect 75177 11794 75243 11797
rect 382365 11794 382431 11797
rect 75177 11792 382431 11794
rect 75177 11736 75182 11792
rect 75238 11736 382370 11792
rect 382426 11736 382431 11792
rect 75177 11734 382431 11736
rect 75177 11731 75243 11734
rect 382365 11731 382431 11734
rect 60549 11658 60615 11661
rect 492305 11658 492371 11661
rect 60549 11656 492371 11658
rect 60549 11600 60554 11656
rect 60610 11600 492310 11656
rect 492366 11600 492371 11656
rect 60549 11598 492371 11600
rect 60549 11595 60615 11598
rect 492305 11595 492371 11598
rect 71589 10434 71655 10437
rect 375281 10434 375347 10437
rect 71589 10432 375347 10434
rect 71589 10376 71594 10432
rect 71650 10376 375286 10432
rect 375342 10376 375347 10432
rect 71589 10374 375347 10376
rect 71589 10371 71655 10374
rect 375281 10371 375347 10374
rect 59169 10298 59235 10301
rect 488809 10298 488875 10301
rect 59169 10296 488875 10298
rect 59169 10240 59174 10296
rect 59230 10240 488814 10296
rect 488870 10240 488875 10296
rect 59169 10238 488875 10240
rect 59169 10235 59235 10238
rect 488809 10235 488875 10238
rect 90449 9074 90515 9077
rect 332685 9074 332751 9077
rect 90449 9072 332751 9074
rect 90449 9016 90454 9072
rect 90510 9016 332690 9072
rect 332746 9016 332751 9072
rect 90449 9014 332751 9016
rect 90449 9011 90515 9014
rect 332685 9011 332751 9014
rect 58617 8938 58683 8941
rect 485221 8938 485287 8941
rect 58617 8936 485287 8938
rect 58617 8880 58622 8936
rect 58678 8880 485226 8936
rect 485282 8880 485287 8936
rect 58617 8878 485287 8880
rect 58617 8875 58683 8878
rect 485221 8875 485287 8878
rect 48957 7850 49023 7853
rect 206277 7850 206343 7853
rect 48957 7848 206343 7850
rect 48957 7792 48962 7848
rect 49018 7792 206282 7848
rect 206338 7792 206343 7848
rect 48957 7790 206343 7792
rect 48957 7787 49023 7790
rect 206277 7787 206343 7790
rect 78581 7714 78647 7717
rect 284334 7714 284340 7716
rect 78581 7712 284340 7714
rect 78581 7656 78586 7712
rect 78642 7656 284340 7712
rect 78581 7654 284340 7656
rect 78581 7651 78647 7654
rect 284334 7652 284340 7654
rect 284404 7652 284410 7716
rect 406377 7714 406443 7717
rect 432045 7714 432111 7717
rect 406377 7712 432111 7714
rect 406377 7656 406382 7712
rect 406438 7656 432050 7712
rect 432106 7656 432111 7712
rect 406377 7654 432111 7656
rect 406377 7651 406443 7654
rect 432045 7651 432111 7654
rect 222694 7578 222700 7580
rect 6870 7518 222700 7578
rect 6870 7034 6930 7518
rect 222694 7516 222700 7518
rect 222764 7516 222770 7580
rect 353937 7578 354003 7581
rect 414289 7578 414355 7581
rect 353937 7576 414355 7578
rect 353937 7520 353942 7576
rect 353998 7520 414294 7576
rect 414350 7520 414355 7576
rect 353937 7518 414355 7520
rect 353937 7515 354003 7518
rect 414289 7515 414355 7518
rect 431217 7578 431283 7581
rect 442625 7578 442691 7581
rect 431217 7576 442691 7578
rect 431217 7520 431222 7576
rect 431278 7520 442630 7576
rect 442686 7520 442691 7576
rect 431217 7518 442691 7520
rect 431217 7515 431283 7518
rect 442625 7515 442691 7518
rect 4110 6974 6930 7034
rect -960 6490 480 6580
rect 4110 6490 4170 6974
rect 72601 6898 72667 6901
rect 261661 6898 261727 6901
rect 72601 6896 261727 6898
rect 72601 6840 72606 6896
rect 72662 6840 261666 6896
rect 261722 6840 261727 6896
rect 72601 6838 261727 6840
rect 72601 6835 72667 6838
rect 261661 6835 261727 6838
rect 62021 6762 62087 6765
rect 258165 6762 258231 6765
rect 62021 6760 258231 6762
rect 62021 6704 62026 6760
rect 62082 6704 258170 6760
rect 258226 6704 258231 6760
rect 62021 6702 258231 6704
rect 62021 6699 62087 6702
rect 258165 6699 258231 6702
rect 58433 6626 58499 6629
rect 256969 6626 257035 6629
rect 58433 6624 257035 6626
rect 58433 6568 58438 6624
rect 58494 6568 256974 6624
rect 257030 6568 257035 6624
rect 58433 6566 257035 6568
rect 58433 6563 58499 6566
rect 256969 6563 257035 6566
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect -960 6430 4170 6490
rect 54937 6490 55003 6493
rect 255773 6490 255839 6493
rect 54937 6488 255839 6490
rect 54937 6432 54942 6488
rect 54998 6432 255778 6488
rect 255834 6432 255839 6488
rect 583520 6476 584960 6566
rect 54937 6430 255839 6432
rect -960 6340 480 6430
rect 54937 6427 55003 6430
rect 255773 6427 255839 6430
rect 47853 6354 47919 6357
rect 253381 6354 253447 6357
rect 47853 6352 253447 6354
rect 47853 6296 47858 6352
rect 47914 6296 253386 6352
rect 253442 6296 253447 6352
rect 47853 6294 253447 6296
rect 47853 6291 47919 6294
rect 253381 6291 253447 6294
rect 12341 6218 12407 6221
rect 242617 6218 242683 6221
rect 12341 6216 242683 6218
rect 12341 6160 12346 6216
rect 12402 6160 242622 6216
rect 242678 6160 242683 6216
rect 12341 6158 242683 6160
rect 12341 6155 12407 6158
rect 242617 6155 242683 6158
rect 76189 6082 76255 6085
rect 262949 6082 263015 6085
rect 76189 6080 263015 6082
rect 76189 6024 76194 6080
rect 76250 6024 262954 6080
rect 263010 6024 263015 6080
rect 76189 6022 263015 6024
rect 76189 6019 76255 6022
rect 262949 6019 263015 6022
rect 109309 5130 109375 5133
rect 146937 5130 147003 5133
rect 109309 5128 147003 5130
rect 109309 5072 109314 5128
rect 109370 5072 146942 5128
rect 146998 5072 147003 5128
rect 109309 5070 147003 5072
rect 109309 5067 109375 5070
rect 146937 5067 147003 5070
rect 273897 5130 273963 5133
rect 283097 5130 283163 5133
rect 273897 5128 283163 5130
rect 273897 5072 273902 5128
rect 273958 5072 283102 5128
rect 283158 5072 283163 5128
rect 273897 5070 283163 5072
rect 273897 5067 273963 5070
rect 283097 5067 283163 5070
rect 7649 4994 7715 4997
rect 241421 4994 241487 4997
rect 7649 4992 241487 4994
rect 7649 4936 7654 4992
rect 7710 4936 241426 4992
rect 241482 4936 241487 4992
rect 7649 4934 241487 4936
rect 7649 4931 7715 4934
rect 241421 4931 241487 4934
rect 246297 4994 246363 4997
rect 286593 4994 286659 4997
rect 246297 4992 286659 4994
rect 246297 4936 246302 4992
rect 246358 4936 286598 4992
rect 286654 4936 286659 4992
rect 246297 4934 286659 4936
rect 246297 4931 246363 4934
rect 286593 4931 286659 4934
rect 55029 4858 55095 4861
rect 290181 4858 290247 4861
rect 55029 4856 290247 4858
rect 55029 4800 55034 4856
rect 55090 4800 290186 4856
rect 290242 4800 290247 4856
rect 55029 4798 290247 4800
rect 55029 4795 55095 4798
rect 290181 4795 290247 4798
rect 351177 4858 351243 4861
rect 410793 4858 410859 4861
rect 351177 4856 410859 4858
rect 351177 4800 351182 4856
rect 351238 4800 410798 4856
rect 410854 4800 410859 4856
rect 351177 4798 410859 4800
rect 351177 4795 351243 4798
rect 410793 4795 410859 4798
rect 411897 4858 411963 4861
rect 417877 4858 417943 4861
rect 411897 4856 417943 4858
rect 411897 4800 411902 4856
rect 411958 4800 417882 4856
rect 417938 4800 417943 4856
rect 411897 4798 417943 4800
rect 411897 4795 411963 4798
rect 417877 4795 417943 4798
rect 429837 4858 429903 4861
rect 435541 4858 435607 4861
rect 429837 4856 435607 4858
rect 429837 4800 429842 4856
rect 429898 4800 435546 4856
rect 435602 4800 435607 4856
rect 429837 4798 435607 4800
rect 429837 4795 429903 4798
rect 435541 4795 435607 4798
rect 450537 4858 450603 4861
rect 453297 4858 453363 4861
rect 450537 4856 453363 4858
rect 450537 4800 450542 4856
rect 450598 4800 453302 4856
rect 453358 4800 453363 4856
rect 450537 4798 453363 4800
rect 450537 4795 450603 4798
rect 453297 4795 453363 4798
rect 418797 4178 418863 4181
rect 421373 4178 421439 4181
rect 418797 4176 421439 4178
rect 418797 4120 418802 4176
rect 418858 4120 421378 4176
rect 421434 4120 421439 4176
rect 418797 4118 421439 4120
rect 418797 4115 418863 4118
rect 421373 4115 421439 4118
rect 422937 4178 423003 4181
rect 424961 4178 425027 4181
rect 422937 4176 425027 4178
rect 422937 4120 422942 4176
rect 422998 4120 424966 4176
rect 425022 4120 425027 4176
rect 422937 4118 425027 4120
rect 422937 4115 423003 4118
rect 424961 4115 425027 4118
rect 425697 4178 425763 4181
rect 428457 4178 428523 4181
rect 425697 4176 428523 4178
rect 425697 4120 425702 4176
rect 425758 4120 428462 4176
rect 428518 4120 428523 4176
rect 425697 4118 428523 4120
rect 425697 4115 425763 4118
rect 428457 4115 428523 4118
rect 436737 4178 436803 4181
rect 439129 4178 439195 4181
rect 436737 4176 439195 4178
rect 436737 4120 436742 4176
rect 436798 4120 439134 4176
rect 439190 4120 439195 4176
rect 436737 4118 439195 4120
rect 436737 4115 436803 4118
rect 439129 4115 439195 4118
rect 443637 4178 443703 4181
rect 446213 4178 446279 4181
rect 443637 4176 446279 4178
rect 443637 4120 443642 4176
rect 443698 4120 446218 4176
rect 446274 4120 446279 4176
rect 443637 4118 446279 4120
rect 443637 4115 443703 4118
rect 446213 4115 446279 4118
rect 447777 4178 447843 4181
rect 449801 4178 449867 4181
rect 447777 4176 449867 4178
rect 447777 4120 447782 4176
rect 447838 4120 449806 4176
rect 449862 4120 449867 4176
rect 447777 4118 449867 4120
rect 447777 4115 447843 4118
rect 449801 4115 449867 4118
rect 1669 4042 1735 4045
rect 7557 4042 7623 4045
rect 1669 4040 7623 4042
rect 1669 3984 1674 4040
rect 1730 3984 7562 4040
rect 7618 3984 7623 4040
rect 1669 3982 7623 3984
rect 1669 3979 1735 3982
rect 7557 3979 7623 3982
rect 244089 4042 244155 4045
rect 280981 4042 281047 4045
rect 244089 4040 281047 4042
rect 244089 3984 244094 4040
rect 244150 3984 280986 4040
rect 281042 3984 281047 4040
rect 244089 3982 281047 3984
rect 244089 3979 244155 3982
rect 280981 3979 281047 3982
rect 439497 4042 439563 4045
rect 442901 4042 442967 4045
rect 439497 4040 442967 4042
rect 439497 3984 439502 4040
rect 439558 3984 442906 4040
rect 442962 3984 442967 4040
rect 439497 3982 442967 3984
rect 439497 3979 439563 3982
rect 442901 3979 442967 3982
rect 508497 4042 508563 4045
rect 510061 4042 510127 4045
rect 508497 4040 510127 4042
rect 508497 3984 508502 4040
rect 508558 3984 510066 4040
rect 510122 3984 510127 4040
rect 508497 3982 510127 3984
rect 508497 3979 508563 3982
rect 510061 3979 510127 3982
rect 576117 4042 576183 4045
rect 577405 4042 577471 4045
rect 576117 4040 577471 4042
rect 576117 3984 576122 4040
rect 576178 3984 577410 4040
rect 577466 3984 577471 4040
rect 576117 3982 577471 3984
rect 576117 3979 576183 3982
rect 577405 3979 577471 3982
rect 118785 3906 118851 3909
rect 126237 3906 126303 3909
rect 118785 3904 126303 3906
rect 118785 3848 118790 3904
rect 118846 3848 126242 3904
rect 126298 3848 126303 3904
rect 118785 3846 126303 3848
rect 118785 3843 118851 3846
rect 126237 3843 126303 3846
rect 240501 3906 240567 3909
rect 280797 3906 280863 3909
rect 240501 3904 280863 3906
rect 240501 3848 240506 3904
rect 240562 3848 280802 3904
rect 280858 3848 280863 3904
rect 240501 3846 280863 3848
rect 240501 3843 240567 3846
rect 280797 3843 280863 3846
rect 421557 3906 421623 3909
rect 463969 3906 464035 3909
rect 421557 3904 464035 3906
rect 421557 3848 421562 3904
rect 421618 3848 463974 3904
rect 464030 3848 464035 3904
rect 421557 3846 464035 3848
rect 421557 3843 421623 3846
rect 463969 3843 464035 3846
rect 67909 3770 67975 3773
rect 101397 3770 101463 3773
rect 67909 3768 101463 3770
rect 67909 3712 67914 3768
rect 67970 3712 101402 3768
rect 101458 3712 101463 3768
rect 67909 3710 101463 3712
rect 67909 3707 67975 3710
rect 101397 3707 101463 3710
rect 119889 3770 119955 3773
rect 163497 3770 163563 3773
rect 119889 3768 163563 3770
rect 119889 3712 119894 3768
rect 119950 3712 163502 3768
rect 163558 3712 163563 3768
rect 119889 3710 163563 3712
rect 119889 3707 119955 3710
rect 163497 3707 163563 3710
rect 169569 3770 169635 3773
rect 287053 3770 287119 3773
rect 169569 3768 287119 3770
rect 169569 3712 169574 3768
rect 169630 3712 287058 3768
rect 287114 3712 287119 3768
rect 169569 3710 287119 3712
rect 169569 3707 169635 3710
rect 287053 3707 287119 3710
rect 428549 3770 428615 3773
rect 471053 3770 471119 3773
rect 428549 3768 471119 3770
rect 428549 3712 428554 3768
rect 428610 3712 471058 3768
rect 471114 3712 471119 3768
rect 428549 3710 471119 3712
rect 428549 3707 428615 3710
rect 471053 3707 471119 3710
rect 13537 3634 13603 3637
rect 119337 3634 119403 3637
rect 13537 3632 119403 3634
rect 13537 3576 13542 3632
rect 13598 3576 119342 3632
rect 119398 3576 119403 3632
rect 13537 3574 119403 3576
rect 13537 3571 13603 3574
rect 119337 3571 119403 3574
rect 124673 3634 124739 3637
rect 291193 3634 291259 3637
rect 124673 3632 291259 3634
rect 124673 3576 124678 3632
rect 124734 3576 291198 3632
rect 291254 3576 291259 3632
rect 124673 3574 291259 3576
rect 124673 3571 124739 3574
rect 291193 3571 291259 3574
rect 435357 3634 435423 3637
rect 478137 3634 478203 3637
rect 435357 3632 478203 3634
rect 435357 3576 435362 3632
rect 435418 3576 478142 3632
rect 478198 3576 478203 3632
rect 435357 3574 478203 3576
rect 435357 3571 435423 3574
rect 478137 3571 478203 3574
rect 28901 3498 28967 3501
rect 32397 3498 32463 3501
rect 28901 3496 32463 3498
rect 28901 3440 28906 3496
rect 28962 3440 32402 3496
rect 32458 3440 32463 3496
rect 28901 3438 32463 3440
rect 28901 3435 28967 3438
rect 32397 3435 32463 3438
rect 50153 3498 50219 3501
rect 51717 3498 51783 3501
rect 50153 3496 51783 3498
rect 50153 3440 50158 3496
rect 50214 3440 51722 3496
rect 51778 3440 51783 3496
rect 50153 3438 51783 3440
rect 50153 3435 50219 3438
rect 51717 3435 51783 3438
rect 57237 3498 57303 3501
rect 91737 3498 91803 3501
rect 57237 3496 91803 3498
rect 57237 3440 57242 3496
rect 57298 3440 91742 3496
rect 91798 3440 91803 3496
rect 57237 3438 91803 3440
rect 57237 3435 57303 3438
rect 91737 3435 91803 3438
rect 117589 3498 117655 3501
rect 288433 3498 288499 3501
rect 117589 3496 288499 3498
rect 117589 3440 117594 3496
rect 117650 3440 288438 3496
rect 288494 3440 288499 3496
rect 117589 3438 288499 3440
rect 117589 3435 117655 3438
rect 288433 3435 288499 3438
rect 417417 3498 417483 3501
rect 460381 3498 460447 3501
rect 417417 3496 460447 3498
rect 417417 3440 417422 3496
rect 417478 3440 460386 3496
rect 460442 3440 460447 3496
rect 417417 3438 460447 3440
rect 417417 3435 417483 3438
rect 460381 3435 460447 3438
rect 512637 3498 512703 3501
rect 513557 3498 513623 3501
rect 512637 3496 513623 3498
rect 512637 3440 512642 3496
rect 512698 3440 513562 3496
rect 513618 3440 513623 3496
rect 512637 3438 513623 3440
rect 512637 3435 512703 3438
rect 513557 3435 513623 3438
rect 562317 3498 562383 3501
rect 563237 3498 563303 3501
rect 562317 3496 563303 3498
rect 562317 3440 562322 3496
rect 562378 3440 563242 3496
rect 563298 3440 563303 3496
rect 562317 3438 563303 3440
rect 562317 3435 562383 3438
rect 563237 3435 563303 3438
rect 9949 3362 10015 3365
rect 25497 3362 25563 3365
rect 9949 3360 25563 3362
rect 9949 3304 9954 3360
rect 10010 3304 25502 3360
rect 25558 3304 25563 3360
rect 9949 3302 25563 3304
rect 9949 3299 10015 3302
rect 25497 3299 25563 3302
rect 60825 3362 60891 3365
rect 271137 3362 271203 3365
rect 272425 3362 272491 3365
rect 60825 3360 258090 3362
rect 60825 3304 60830 3360
rect 60886 3304 258090 3360
rect 60825 3302 258090 3304
rect 60825 3299 60891 3302
rect 258030 3226 258090 3302
rect 271137 3360 272491 3362
rect 271137 3304 271142 3360
rect 271198 3304 272430 3360
rect 272486 3304 272491 3360
rect 271137 3302 272491 3304
rect 271137 3299 271203 3302
rect 272425 3299 272491 3302
rect 278037 3362 278103 3365
rect 279509 3362 279575 3365
rect 278037 3360 279575 3362
rect 278037 3304 278042 3360
rect 278098 3304 279514 3360
rect 279570 3304 279575 3360
rect 278037 3302 279575 3304
rect 278037 3299 278103 3302
rect 279509 3299 279575 3302
rect 284937 3362 285003 3365
rect 371693 3362 371759 3365
rect 284937 3360 371759 3362
rect 284937 3304 284942 3360
rect 284998 3304 371698 3360
rect 371754 3304 371759 3360
rect 284937 3302 371759 3304
rect 284937 3299 285003 3302
rect 371693 3299 371759 3302
rect 442257 3362 442323 3365
rect 582189 3362 582255 3365
rect 442257 3360 582255 3362
rect 442257 3304 442262 3360
rect 442318 3304 582194 3360
rect 582250 3304 582255 3360
rect 442257 3302 582255 3304
rect 442257 3299 442323 3302
rect 582189 3299 582255 3302
rect 280061 3226 280127 3229
rect 258030 3224 280127 3226
rect 258030 3168 280066 3224
rect 280122 3168 280127 3224
rect 258030 3166 280127 3168
rect 280061 3163 280127 3166
rect 432597 3226 432663 3229
rect 474549 3226 474615 3229
rect 432597 3224 474615 3226
rect 432597 3168 432602 3224
rect 432658 3168 474554 3224
rect 474610 3168 474615 3224
rect 432597 3166 474615 3168
rect 432597 3163 432663 3166
rect 474549 3163 474615 3166
rect 414657 3090 414723 3093
rect 456885 3090 456951 3093
rect 414657 3088 456951 3090
rect 414657 3032 414662 3088
rect 414718 3032 456890 3088
rect 456946 3032 456951 3088
rect 414657 3030 456951 3032
rect 414657 3027 414723 3030
rect 456885 3027 456951 3030
rect 19425 2954 19491 2957
rect 243537 2954 243603 2957
rect 19425 2952 243603 2954
rect 19425 2896 19430 2952
rect 19486 2896 243542 2952
rect 243598 2896 243603 2952
rect 19425 2894 243603 2896
rect 19425 2891 19491 2894
rect 243537 2891 243603 2894
rect 32397 2818 32463 2821
rect 271781 2818 271847 2821
rect 32397 2816 271847 2818
rect 32397 2760 32402 2816
rect 32458 2760 271786 2816
rect 271842 2760 271847 2816
rect 32397 2758 271847 2760
rect 32397 2755 32463 2758
rect 271781 2755 271847 2758
<< via3 >>
rect 355180 683844 355244 683908
rect 57284 671196 57348 671260
rect 2820 658140 2884 658204
rect 501644 655556 501708 655620
rect 500356 654936 500420 654940
rect 500356 654880 500406 654936
rect 500406 654880 500420 654936
rect 500356 654876 500420 654880
rect 501644 654332 501708 654396
rect 500356 653380 500420 653444
rect 542676 636244 542740 636308
rect 580212 630804 580276 630868
rect 68508 626588 68572 626652
rect 291148 626316 291212 626380
rect 68692 622236 68756 622300
rect 290596 622236 290660 622300
rect 3004 619108 3068 619172
rect 541020 618564 541084 618628
rect 291700 618156 291764 618220
rect 68876 617884 68940 617948
rect 291516 614076 291580 614140
rect 70164 613532 70228 613596
rect 291332 609996 291396 610060
rect 68140 609180 68204 609244
rect 542860 607684 542924 607748
rect 543044 606324 543108 606388
rect 3372 606052 3436 606116
rect 543228 604964 543292 605028
rect 68324 604828 68388 604892
rect 68508 604420 68572 604484
rect 539364 603604 539428 603668
rect 68692 601080 68756 601084
rect 68692 601024 68706 601080
rect 68706 601024 68756 601080
rect 68692 601020 68756 601024
rect 68508 600476 68572 600540
rect 69612 596124 69676 596188
rect 63356 591772 63420 591836
rect 306972 591228 307036 591292
rect 580212 591228 580276 591292
rect 63172 587420 63236 587484
rect 69980 582524 70044 582588
rect 290780 581436 290844 581500
rect 69428 578716 69492 578780
rect 313780 577628 313844 577692
rect 66852 574364 66916 574428
rect 70164 571236 70228 571300
rect 69796 570012 69860 570076
rect 3556 566884 3620 566948
rect 65564 565660 65628 565724
rect 67404 561308 67468 561372
rect 67220 556956 67284 557020
rect 3740 553828 3804 553892
rect 3004 553420 3068 553484
rect 66116 552604 66180 552668
rect 67036 548252 67100 548316
rect 65932 543900 65996 543964
rect 66852 540908 66916 540972
rect 66852 539548 66916 539612
rect 65748 535196 65812 535260
rect 68876 531252 68940 531316
rect 68692 530844 68756 530908
rect 68876 526492 68940 526556
rect 68140 525812 68204 525876
rect 309732 524452 309796 524516
rect 68324 522956 68388 523020
rect 67956 522140 68020 522204
rect 68140 517788 68204 517852
rect 68508 517516 68572 517580
rect 289308 516156 289372 516220
rect 59860 514796 59924 514860
rect 68692 513980 68756 514044
rect 68692 513436 68756 513500
rect 68508 509084 68572 509148
rect 68876 507860 68940 507924
rect 62988 504732 63052 504796
rect 2820 502284 2884 502348
rect 3924 501740 3988 501804
rect 67956 500788 68020 500852
rect 68324 500380 68388 500444
rect 69612 496300 69676 496364
rect 69612 496028 69676 496092
rect 65564 492628 65628 492692
rect 65564 491676 65628 491740
rect 580212 484604 580276 484668
rect 291700 481068 291764 481132
rect 290596 480116 290660 480180
rect 290780 479980 290844 480044
rect 234476 479436 234540 479500
rect 543228 479436 543292 479500
rect 232268 478076 232332 478140
rect 580212 478076 580276 478140
rect 240916 477804 240980 477868
rect 291516 477940 291580 478004
rect 68324 476852 68388 476916
rect 203380 476852 203444 476916
rect 239812 476716 239876 476780
rect 542676 476716 542740 476780
rect 68508 474132 68572 474196
rect 166212 474132 166276 474196
rect 234292 473996 234356 474060
rect 543044 473996 543108 474060
rect 3740 472500 3804 472564
rect 161980 472500 162044 472564
rect 224540 472364 224604 472428
rect 224724 471956 224788 472020
rect 238340 471956 238404 472020
rect 289308 471412 289372 471476
rect 574692 471412 574756 471476
rect 3924 471140 3988 471204
rect 130332 471140 130396 471204
rect 68692 469780 68756 469844
rect 208900 469780 208964 469844
rect 291332 468692 291396 468756
rect 238524 468420 238588 468484
rect 539364 468420 539428 468484
rect 3556 467332 3620 467396
rect 282868 467332 282932 467396
rect 287100 462572 287164 462636
rect 68140 461484 68204 461548
rect 173020 461484 173084 461548
rect 235764 458764 235828 458828
rect 291148 456180 291212 456244
rect 3372 456044 3436 456108
rect 210372 456044 210436 456108
rect 238156 456044 238220 456108
rect 541020 456044 541084 456108
rect 234108 450468 234172 450532
rect 542860 450468 542924 450532
rect 227668 449516 227732 449580
rect 237236 449516 237300 449580
rect 237972 449244 238036 449308
rect 235580 446524 235644 446588
rect 57284 444212 57348 444276
rect 59860 443940 59924 444004
rect 235212 444076 235276 444140
rect 287284 443940 287348 444004
rect 224908 442308 224972 442372
rect 223988 442036 224052 442100
rect 218836 441900 218900 441964
rect 218652 441764 218716 441828
rect 221044 441628 221108 441692
rect 233924 441688 233988 441692
rect 233924 441632 233974 441688
rect 233974 441632 233988 441688
rect 233924 441628 233988 441632
rect 228404 441492 228468 441556
rect 226932 441356 226996 441420
rect 112484 441220 112548 441284
rect 280660 441220 280724 441284
rect 230980 441084 231044 441148
rect 219940 440948 220004 441012
rect 230060 440948 230124 441012
rect 112300 440540 112364 440604
rect 112852 440404 112916 440468
rect 278820 440404 278884 440468
rect 226196 440268 226260 440332
rect 227852 440268 227916 440332
rect 230428 440268 230492 440332
rect 231900 440268 231964 440332
rect 222700 440132 222764 440196
rect 227668 440132 227732 440196
rect 228220 439860 228284 439924
rect 281948 439860 282012 439924
rect 224172 439724 224236 439788
rect 281764 439724 281828 439788
rect 227116 439588 227180 439652
rect 282316 439588 282380 439652
rect 178540 439452 178604 439516
rect 221228 439316 221292 439380
rect 231532 439316 231596 439380
rect 227668 439180 227732 439244
rect 229876 439044 229940 439108
rect 239628 439044 239692 439108
rect 112668 438908 112732 438972
rect 279372 438908 279436 438972
rect 280844 438908 280908 438972
rect 278820 438636 278884 438700
rect 231164 438500 231228 438564
rect 279556 438500 279620 438564
rect 279372 437412 279436 437476
rect 281948 431564 282012 431628
rect 281764 430204 281828 430268
rect 282316 428844 282380 428908
rect 280844 426124 280908 426188
rect 280660 423404 280724 423468
rect 500172 418236 500236 418300
rect 223988 410484 224052 410548
rect 224356 409940 224420 410004
rect 239444 405996 239508 406060
rect 240180 401508 240244 401572
rect 173204 397428 173268 397492
rect 279556 396204 279620 396268
rect 287468 392124 287532 392188
rect 287652 390764 287716 390828
rect 235580 368732 235644 368796
rect 580212 365060 580276 365124
rect 235396 358396 235460 358460
rect 237972 347712 238036 347716
rect 237972 347656 237986 347712
rect 237986 347656 238036 347712
rect 237972 347652 238036 347656
rect 69980 347108 70044 347172
rect 237420 347108 237484 347172
rect 147076 345204 147140 345268
rect 69612 344932 69676 344996
rect 62988 344660 63052 344724
rect 223068 344660 223132 344724
rect 63172 344388 63236 344452
rect 63356 343980 63420 344044
rect 67404 342136 67468 342140
rect 67404 342080 67454 342136
rect 67454 342080 67468 342136
rect 67404 342076 67468 342080
rect 69796 342076 69860 342140
rect 69428 341940 69492 342004
rect 66116 341804 66180 341868
rect 66852 341668 66916 341732
rect 234660 341668 234724 341732
rect 65748 341532 65812 341596
rect 235028 341532 235092 341596
rect 65932 341396 65996 341460
rect 235580 341396 235644 341460
rect 67036 341260 67100 341324
rect 67220 341124 67284 341188
rect 65564 340988 65628 341052
rect 235212 340988 235276 341052
rect 235764 340852 235828 340916
rect 111748 339356 111812 339420
rect 280844 339084 280908 339148
rect 112852 338540 112916 338604
rect 178540 336908 178604 336972
rect 230060 335276 230124 335340
rect 230244 334112 230308 334116
rect 230244 334056 230294 334112
rect 230294 334056 230308 334112
rect 230244 334052 230308 334056
rect 219940 333644 220004 333708
rect 228404 332012 228468 332076
rect 228036 331332 228100 331396
rect 227116 330380 227180 330444
rect 299980 329020 300044 329084
rect 580212 329020 580276 329084
rect 224172 328748 224236 328812
rect 222700 327116 222764 327180
rect 239444 326300 239508 326364
rect 231532 325484 231596 325548
rect 580212 325212 580276 325276
rect 230612 324396 230676 324460
rect 112668 323852 112732 323916
rect 239812 323036 239876 323100
rect 111932 322900 111996 322964
rect 226932 322220 226996 322284
rect 112484 320588 112548 320652
rect 230980 318956 231044 319020
rect 285628 318684 285692 318748
rect 224356 318140 224420 318204
rect 229876 317324 229940 317388
rect 284340 317324 284404 317388
rect 238340 317052 238404 317116
rect 238340 316916 238404 316980
rect 224540 316508 224604 316572
rect 238156 315964 238220 316028
rect 228220 315692 228284 315756
rect 224724 315420 224788 315484
rect 280660 314604 280724 314668
rect 231900 314060 231964 314124
rect 232084 313244 232148 313308
rect 111748 312428 111812 312492
rect 544332 312020 544396 312084
rect 234108 311612 234172 311676
rect 234292 311068 234356 311132
rect 230428 310796 230492 310860
rect 234476 310524 234540 310588
rect 238524 309980 238588 310044
rect 233924 309436 233988 309500
rect 112300 309164 112364 309228
rect 222700 308892 222764 308956
rect 224172 308348 224236 308412
rect 230980 307804 231044 307868
rect 284524 307804 284588 307868
rect 234660 307668 234724 307732
rect 111932 307532 111996 307596
rect 235212 307260 235276 307324
rect 228220 306716 228284 306780
rect 48636 306172 48700 306236
rect 231348 306172 231412 306236
rect 122052 305628 122116 305692
rect 147076 305084 147140 305148
rect 173204 304540 173268 304604
rect 218836 304268 218900 304332
rect 279372 303724 279436 303788
rect 130332 303452 130396 303516
rect 161980 302908 162044 302972
rect 218652 302636 218716 302700
rect 210372 302364 210436 302428
rect 281764 302364 281828 302428
rect 221044 301004 221108 301068
rect 284708 301004 284772 301068
rect 282132 299644 282196 299708
rect 237236 298012 237300 298076
rect 221228 297740 221292 297804
rect 224908 296108 224972 296172
rect 232084 295836 232148 295900
rect 224908 295292 224972 295356
rect 238340 295292 238404 295356
rect 230244 294748 230308 294812
rect 228036 294476 228100 294540
rect 232268 294204 232332 294268
rect 284892 294204 284956 294268
rect 239628 293660 239692 293724
rect 3372 293116 3436 293180
rect 238156 293116 238220 293180
rect 227852 292844 227916 292908
rect 281580 292844 281644 292908
rect 238524 292572 238588 292636
rect 238340 292028 238404 292092
rect 239260 291484 239324 291548
rect 281028 291484 281092 291548
rect 227668 291212 227732 291276
rect 239444 290940 239508 291004
rect 239628 290396 239692 290460
rect 283052 290124 283116 290188
rect 239812 289852 239876 289916
rect 230612 289580 230676 289644
rect 231164 287948 231228 288012
rect 288388 287404 288452 287468
rect 224908 286316 224972 286380
rect 283420 286044 283484 286108
rect 226196 284684 226260 284748
rect 283236 284684 283300 284748
rect 287836 283324 287900 283388
rect 237972 283052 238036 283116
rect 237420 282916 237484 282980
rect 287284 282916 287348 282980
rect 287284 281964 287348 282028
rect 287100 281828 287164 281892
rect 237788 281420 237852 281484
rect 238156 281420 238220 281484
rect 3372 279380 3436 279444
rect 122052 279380 122116 279444
rect 235028 276796 235092 276860
rect 282868 276524 282932 276588
rect 173020 274620 173084 274684
rect 282132 274620 282196 274684
rect 208900 274076 208964 274140
rect 166212 273532 166276 273596
rect 223068 272988 223132 273052
rect 203380 272444 203444 272508
rect 580396 272172 580460 272236
rect 235580 271356 235644 271420
rect 355180 260204 355244 260268
rect 306972 258844 307036 258908
rect 320772 258844 320836 258908
rect 313780 257484 313844 257548
rect 309732 256124 309796 256188
rect 574692 254764 574756 254828
rect 3372 254084 3436 254148
rect 500172 253404 500236 253468
rect 299980 252044 300044 252108
rect 544332 250684 544396 250748
rect 320772 249324 320836 249388
rect 355180 247964 355244 248028
rect 353892 246604 353956 246668
rect 346900 245244 346964 245308
rect 500172 243884 500236 243948
rect 559420 242524 559484 242588
rect 231348 242116 231412 242180
rect 279556 241844 279620 241908
rect 287100 241436 287164 241500
rect 457300 241164 457364 241228
rect 287652 240892 287716 240956
rect 3372 240620 3436 240684
rect 283236 240620 283300 240684
rect 235396 240484 235460 240548
rect 287284 240484 287348 240548
rect 237788 240348 237852 240412
rect 284708 240076 284772 240140
rect 238524 239940 238588 240004
rect 580212 239940 580276 240004
rect 48636 239804 48700 239868
rect 287836 239804 287900 239868
rect 237972 239668 238036 239732
rect 287468 239668 287532 239732
rect 238340 238988 238404 239052
rect 580396 238988 580460 239052
rect 284892 235316 284956 235380
rect 281764 233820 281828 233884
rect 239260 232324 239324 232388
rect 279372 228244 279436 228308
rect 279556 225524 279620 225588
rect 280844 220220 280908 220284
rect 355180 218996 355244 219060
rect 281580 218588 281644 218652
rect 3556 217228 3620 217292
rect 283052 217228 283116 217292
rect 3740 215868 3804 215932
rect 283420 215868 283484 215932
rect 3372 202132 3436 202196
rect 281028 202132 281092 202196
rect 3740 201860 3804 201924
rect 239444 192476 239508 192540
rect 228220 188804 228284 188868
rect 353892 179148 353956 179212
rect 239628 152628 239692 152692
rect 288388 149772 288452 149836
rect 346900 139300 346964 139364
rect 235212 136716 235276 136780
rect 239812 112780 239876 112844
rect 500172 99452 500236 99516
rect 287100 97548 287164 97612
rect 3188 86260 3252 86324
rect 230980 86260 231044 86324
rect 3188 84628 3252 84692
rect 559420 59604 559484 59668
rect 3556 58516 3620 58580
rect 224172 45460 224236 45524
rect 280660 32540 280724 32604
rect 285628 29684 285692 29748
rect 284524 26964 284588 27028
rect 457300 19756 457364 19820
rect 3372 19348 3436 19412
rect 284340 7652 284404 7716
rect 222700 7516 222764 7580
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 677494 -8106 711002
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 -8106 677494
rect -8726 677174 -8106 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 -8106 677174
rect -8726 641494 -8106 676938
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 -8106 641494
rect -8726 641174 -8106 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 -8106 641174
rect -8726 605494 -8106 640938
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 -8106 605494
rect -8726 605174 -8106 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 -8106 605174
rect -8726 569494 -8106 604938
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 -8106 569494
rect -8726 569174 -8106 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 -8106 569174
rect -8726 533494 -8106 568938
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 -8106 533494
rect -8726 533174 -8106 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 -8106 533174
rect -8726 497494 -8106 532938
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 -8106 497494
rect -8726 497174 -8106 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 -8106 497174
rect -8726 461494 -8106 496938
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 -8106 461494
rect -8726 461174 -8106 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 -8106 461174
rect -8726 425494 -8106 460938
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 -8106 425494
rect -8726 425174 -8106 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 -8106 425174
rect -8726 389494 -8106 424938
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 -8106 389494
rect -8726 389174 -8106 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 -8106 389174
rect -8726 353494 -8106 388938
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 -8106 353494
rect -8726 353174 -8106 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 -8106 353174
rect -8726 317494 -8106 352938
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 -8106 317494
rect -8726 317174 -8106 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 -8106 317174
rect -8726 281494 -8106 316938
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 -8106 281494
rect -8726 281174 -8106 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 -8106 281174
rect -8726 245494 -8106 280938
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 -8106 245494
rect -8726 245174 -8106 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 -8106 245174
rect -8726 209494 -8106 244938
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 -8106 209494
rect -8726 209174 -8106 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 -8106 209174
rect -8726 173494 -8106 208938
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 -8106 173494
rect -8726 173174 -8106 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 -8106 173174
rect -8726 137494 -8106 172938
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 -8106 137494
rect -8726 137174 -8106 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 -8106 137174
rect -8726 101494 -8106 136938
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 -8106 101494
rect -8726 101174 -8106 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 -8106 101174
rect -8726 65494 -8106 100938
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 -8106 65494
rect -8726 65174 -8106 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 -8106 65174
rect -8726 29494 -8106 64938
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 -8106 29494
rect -8726 29174 -8106 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 -8106 29174
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 673774 -7146 710042
rect -7766 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 -7146 673774
rect -7766 673454 -7146 673538
rect -7766 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 -7146 673454
rect -7766 637774 -7146 673218
rect -7766 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 -7146 637774
rect -7766 637454 -7146 637538
rect -7766 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 -7146 637454
rect -7766 601774 -7146 637218
rect -7766 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 -7146 601774
rect -7766 601454 -7146 601538
rect -7766 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 -7146 601454
rect -7766 565774 -7146 601218
rect -7766 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 -7146 565774
rect -7766 565454 -7146 565538
rect -7766 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 -7146 565454
rect -7766 529774 -7146 565218
rect -7766 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 -7146 529774
rect -7766 529454 -7146 529538
rect -7766 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 -7146 529454
rect -7766 493774 -7146 529218
rect -7766 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 -7146 493774
rect -7766 493454 -7146 493538
rect -7766 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 -7146 493454
rect -7766 457774 -7146 493218
rect -7766 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 -7146 457774
rect -7766 457454 -7146 457538
rect -7766 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 -7146 457454
rect -7766 421774 -7146 457218
rect -7766 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 -7146 421774
rect -7766 421454 -7146 421538
rect -7766 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 -7146 421454
rect -7766 385774 -7146 421218
rect -7766 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 -7146 385774
rect -7766 385454 -7146 385538
rect -7766 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 -7146 385454
rect -7766 349774 -7146 385218
rect -7766 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 -7146 349774
rect -7766 349454 -7146 349538
rect -7766 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 -7146 349454
rect -7766 313774 -7146 349218
rect -7766 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 -7146 313774
rect -7766 313454 -7146 313538
rect -7766 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 -7146 313454
rect -7766 277774 -7146 313218
rect -7766 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 -7146 277774
rect -7766 277454 -7146 277538
rect -7766 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 -7146 277454
rect -7766 241774 -7146 277218
rect -7766 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 -7146 241774
rect -7766 241454 -7146 241538
rect -7766 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 -7146 241454
rect -7766 205774 -7146 241218
rect -7766 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 -7146 205774
rect -7766 205454 -7146 205538
rect -7766 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 -7146 205454
rect -7766 169774 -7146 205218
rect -7766 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 -7146 169774
rect -7766 169454 -7146 169538
rect -7766 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 -7146 169454
rect -7766 133774 -7146 169218
rect -7766 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 -7146 133774
rect -7766 133454 -7146 133538
rect -7766 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 -7146 133454
rect -7766 97774 -7146 133218
rect -7766 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 -7146 97774
rect -7766 97454 -7146 97538
rect -7766 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 -7146 97454
rect -7766 61774 -7146 97218
rect -7766 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 -7146 61774
rect -7766 61454 -7146 61538
rect -7766 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 -7146 61454
rect -7766 25774 -7146 61218
rect -7766 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 -7146 25774
rect -7766 25454 -7146 25538
rect -7766 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 -7146 25454
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 670054 -6186 709082
rect -6806 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 -6186 670054
rect -6806 669734 -6186 669818
rect -6806 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 -6186 669734
rect -6806 634054 -6186 669498
rect -6806 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 -6186 634054
rect -6806 633734 -6186 633818
rect -6806 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 -6186 633734
rect -6806 598054 -6186 633498
rect -6806 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 -6186 598054
rect -6806 597734 -6186 597818
rect -6806 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 -6186 597734
rect -6806 562054 -6186 597498
rect -6806 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 -6186 562054
rect -6806 561734 -6186 561818
rect -6806 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 -6186 561734
rect -6806 526054 -6186 561498
rect -6806 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 -6186 526054
rect -6806 525734 -6186 525818
rect -6806 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 -6186 525734
rect -6806 490054 -6186 525498
rect -6806 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 -6186 490054
rect -6806 489734 -6186 489818
rect -6806 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 -6186 489734
rect -6806 454054 -6186 489498
rect -6806 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 -6186 454054
rect -6806 453734 -6186 453818
rect -6806 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 -6186 453734
rect -6806 418054 -6186 453498
rect -6806 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 -6186 418054
rect -6806 417734 -6186 417818
rect -6806 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 -6186 417734
rect -6806 382054 -6186 417498
rect -6806 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 -6186 382054
rect -6806 381734 -6186 381818
rect -6806 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 -6186 381734
rect -6806 346054 -6186 381498
rect -6806 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 -6186 346054
rect -6806 345734 -6186 345818
rect -6806 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 -6186 345734
rect -6806 310054 -6186 345498
rect -6806 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 -6186 310054
rect -6806 309734 -6186 309818
rect -6806 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 -6186 309734
rect -6806 274054 -6186 309498
rect -6806 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 -6186 274054
rect -6806 273734 -6186 273818
rect -6806 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 -6186 273734
rect -6806 238054 -6186 273498
rect -6806 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 -6186 238054
rect -6806 237734 -6186 237818
rect -6806 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 -6186 237734
rect -6806 202054 -6186 237498
rect -6806 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 -6186 202054
rect -6806 201734 -6186 201818
rect -6806 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 -6186 201734
rect -6806 166054 -6186 201498
rect -6806 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 -6186 166054
rect -6806 165734 -6186 165818
rect -6806 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 -6186 165734
rect -6806 130054 -6186 165498
rect -6806 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 -6186 130054
rect -6806 129734 -6186 129818
rect -6806 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 -6186 129734
rect -6806 94054 -6186 129498
rect -6806 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 -6186 94054
rect -6806 93734 -6186 93818
rect -6806 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 -6186 93734
rect -6806 58054 -6186 93498
rect -6806 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 -6186 58054
rect -6806 57734 -6186 57818
rect -6806 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 -6186 57734
rect -6806 22054 -6186 57498
rect -6806 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 -6186 22054
rect -6806 21734 -6186 21818
rect -6806 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 -6186 21734
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 666334 -5226 708122
rect -5846 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 -5226 666334
rect -5846 666014 -5226 666098
rect -5846 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 -5226 666014
rect -5846 630334 -5226 665778
rect -5846 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 -5226 630334
rect -5846 630014 -5226 630098
rect -5846 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 -5226 630014
rect -5846 594334 -5226 629778
rect -5846 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 -5226 594334
rect -5846 594014 -5226 594098
rect -5846 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 -5226 594014
rect -5846 558334 -5226 593778
rect -5846 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 -5226 558334
rect -5846 558014 -5226 558098
rect -5846 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 -5226 558014
rect -5846 522334 -5226 557778
rect -5846 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 -5226 522334
rect -5846 522014 -5226 522098
rect -5846 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 -5226 522014
rect -5846 486334 -5226 521778
rect -5846 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 -5226 486334
rect -5846 486014 -5226 486098
rect -5846 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 -5226 486014
rect -5846 450334 -5226 485778
rect -5846 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 -5226 450334
rect -5846 450014 -5226 450098
rect -5846 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 -5226 450014
rect -5846 414334 -5226 449778
rect -5846 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 -5226 414334
rect -5846 414014 -5226 414098
rect -5846 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 -5226 414014
rect -5846 378334 -5226 413778
rect -5846 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 -5226 378334
rect -5846 378014 -5226 378098
rect -5846 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 -5226 378014
rect -5846 342334 -5226 377778
rect -5846 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 -5226 342334
rect -5846 342014 -5226 342098
rect -5846 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 -5226 342014
rect -5846 306334 -5226 341778
rect -5846 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 -5226 306334
rect -5846 306014 -5226 306098
rect -5846 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 -5226 306014
rect -5846 270334 -5226 305778
rect -5846 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 -5226 270334
rect -5846 270014 -5226 270098
rect -5846 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 -5226 270014
rect -5846 234334 -5226 269778
rect -5846 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 -5226 234334
rect -5846 234014 -5226 234098
rect -5846 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 -5226 234014
rect -5846 198334 -5226 233778
rect -5846 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 -5226 198334
rect -5846 198014 -5226 198098
rect -5846 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 -5226 198014
rect -5846 162334 -5226 197778
rect -5846 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 -5226 162334
rect -5846 162014 -5226 162098
rect -5846 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 -5226 162014
rect -5846 126334 -5226 161778
rect -5846 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 -5226 126334
rect -5846 126014 -5226 126098
rect -5846 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 -5226 126014
rect -5846 90334 -5226 125778
rect -5846 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 -5226 90334
rect -5846 90014 -5226 90098
rect -5846 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 -5226 90014
rect -5846 54334 -5226 89778
rect -5846 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 -5226 54334
rect -5846 54014 -5226 54098
rect -5846 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 -5226 54014
rect -5846 18334 -5226 53778
rect -5846 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 -5226 18334
rect -5846 18014 -5226 18098
rect -5846 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 -5226 18014
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 698614 -4266 707162
rect -4886 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 -4266 698614
rect -4886 698294 -4266 698378
rect -4886 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 -4266 698294
rect -4886 662614 -4266 698058
rect -4886 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 -4266 662614
rect -4886 662294 -4266 662378
rect -4886 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 -4266 662294
rect -4886 626614 -4266 662058
rect -4886 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 -4266 626614
rect -4886 626294 -4266 626378
rect -4886 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 -4266 626294
rect -4886 590614 -4266 626058
rect -4886 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 -4266 590614
rect -4886 590294 -4266 590378
rect -4886 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 -4266 590294
rect -4886 554614 -4266 590058
rect -4886 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 -4266 554614
rect -4886 554294 -4266 554378
rect -4886 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 -4266 554294
rect -4886 518614 -4266 554058
rect -4886 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 -4266 518614
rect -4886 518294 -4266 518378
rect -4886 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 -4266 518294
rect -4886 482614 -4266 518058
rect -4886 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 -4266 482614
rect -4886 482294 -4266 482378
rect -4886 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 -4266 482294
rect -4886 446614 -4266 482058
rect -4886 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 -4266 446614
rect -4886 446294 -4266 446378
rect -4886 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 -4266 446294
rect -4886 410614 -4266 446058
rect -4886 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 -4266 410614
rect -4886 410294 -4266 410378
rect -4886 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 -4266 410294
rect -4886 374614 -4266 410058
rect -4886 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 -4266 374614
rect -4886 374294 -4266 374378
rect -4886 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 -4266 374294
rect -4886 338614 -4266 374058
rect -4886 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 -4266 338614
rect -4886 338294 -4266 338378
rect -4886 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 -4266 338294
rect -4886 302614 -4266 338058
rect -4886 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 -4266 302614
rect -4886 302294 -4266 302378
rect -4886 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 -4266 302294
rect -4886 266614 -4266 302058
rect -4886 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 -4266 266614
rect -4886 266294 -4266 266378
rect -4886 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 -4266 266294
rect -4886 230614 -4266 266058
rect -4886 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 -4266 230614
rect -4886 230294 -4266 230378
rect -4886 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 -4266 230294
rect -4886 194614 -4266 230058
rect -4886 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 -4266 194614
rect -4886 194294 -4266 194378
rect -4886 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 -4266 194294
rect -4886 158614 -4266 194058
rect -4886 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 -4266 158614
rect -4886 158294 -4266 158378
rect -4886 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 -4266 158294
rect -4886 122614 -4266 158058
rect -4886 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 -4266 122614
rect -4886 122294 -4266 122378
rect -4886 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 -4266 122294
rect -4886 86614 -4266 122058
rect -4886 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 -4266 86614
rect -4886 86294 -4266 86378
rect -4886 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 -4266 86294
rect -4886 50614 -4266 86058
rect -4886 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 -4266 50614
rect -4886 50294 -4266 50378
rect -4886 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 -4266 50294
rect -4886 14614 -4266 50058
rect -4886 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 -4266 14614
rect -4886 14294 -4266 14378
rect -4886 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 -4266 14294
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 694894 -3306 706202
rect -3926 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 -3306 694894
rect -3926 694574 -3306 694658
rect -3926 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 -3306 694574
rect -3926 658894 -3306 694338
rect -3926 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 -3306 658894
rect -3926 658574 -3306 658658
rect -3926 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 -3306 658574
rect -3926 622894 -3306 658338
rect -3926 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 -3306 622894
rect -3926 622574 -3306 622658
rect -3926 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 -3306 622574
rect -3926 586894 -3306 622338
rect -3926 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 -3306 586894
rect -3926 586574 -3306 586658
rect -3926 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 -3306 586574
rect -3926 550894 -3306 586338
rect -3926 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 -3306 550894
rect -3926 550574 -3306 550658
rect -3926 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 -3306 550574
rect -3926 514894 -3306 550338
rect -3926 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 -3306 514894
rect -3926 514574 -3306 514658
rect -3926 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 -3306 514574
rect -3926 478894 -3306 514338
rect -3926 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 -3306 478894
rect -3926 478574 -3306 478658
rect -3926 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 -3306 478574
rect -3926 442894 -3306 478338
rect -3926 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 -3306 442894
rect -3926 442574 -3306 442658
rect -3926 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 -3306 442574
rect -3926 406894 -3306 442338
rect -3926 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 -3306 406894
rect -3926 406574 -3306 406658
rect -3926 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 -3306 406574
rect -3926 370894 -3306 406338
rect -3926 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 -3306 370894
rect -3926 370574 -3306 370658
rect -3926 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 -3306 370574
rect -3926 334894 -3306 370338
rect -3926 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 -3306 334894
rect -3926 334574 -3306 334658
rect -3926 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 -3306 334574
rect -3926 298894 -3306 334338
rect -3926 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 -3306 298894
rect -3926 298574 -3306 298658
rect -3926 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 -3306 298574
rect -3926 262894 -3306 298338
rect -3926 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 -3306 262894
rect -3926 262574 -3306 262658
rect -3926 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 -3306 262574
rect -3926 226894 -3306 262338
rect -3926 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 -3306 226894
rect -3926 226574 -3306 226658
rect -3926 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 -3306 226574
rect -3926 190894 -3306 226338
rect -3926 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 -3306 190894
rect -3926 190574 -3306 190658
rect -3926 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 -3306 190574
rect -3926 154894 -3306 190338
rect -3926 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 -3306 154894
rect -3926 154574 -3306 154658
rect -3926 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 -3306 154574
rect -3926 118894 -3306 154338
rect -3926 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 -3306 118894
rect -3926 118574 -3306 118658
rect -3926 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 -3306 118574
rect -3926 82894 -3306 118338
rect -3926 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 -3306 82894
rect -3926 82574 -3306 82658
rect -3926 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 -3306 82574
rect -3926 46894 -3306 82338
rect -3926 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 -3306 46894
rect -3926 46574 -3306 46658
rect -3926 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 -3306 46574
rect -3926 10894 -3306 46338
rect -3926 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 -3306 10894
rect -3926 10574 -3306 10658
rect -3926 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 -3306 10574
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 5514 705798 6134 711590
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 2819 658204 2885 658205
rect 2819 658140 2820 658204
rect 2884 658140 2885 658204
rect 2819 658139 2885 658140
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 2822 502349 2882 658139
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 3003 619172 3069 619173
rect 3003 619108 3004 619172
rect 3068 619108 3069 619172
rect 3003 619107 3069 619108
rect 3006 553485 3066 619107
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 3371 606116 3437 606117
rect 3371 606052 3372 606116
rect 3436 606052 3437 606116
rect 3371 606051 3437 606052
rect 3003 553484 3069 553485
rect 3003 553420 3004 553484
rect 3068 553420 3069 553484
rect 3003 553419 3069 553420
rect 2819 502348 2885 502349
rect 2819 502284 2820 502348
rect 2884 502284 2885 502348
rect 2819 502283 2885 502284
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 3374 456109 3434 606051
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 3555 566948 3621 566949
rect 3555 566884 3556 566948
rect 3620 566884 3621 566948
rect 3555 566883 3621 566884
rect 3558 467397 3618 566883
rect 3739 553892 3805 553893
rect 3739 553828 3740 553892
rect 3804 553828 3805 553892
rect 3739 553827 3805 553828
rect 3742 472565 3802 553827
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 3923 501804 3989 501805
rect 3923 501740 3924 501804
rect 3988 501740 3989 501804
rect 3923 501739 3989 501740
rect 3739 472564 3805 472565
rect 3739 472500 3740 472564
rect 3804 472500 3805 472564
rect 3739 472499 3805 472500
rect 3926 471205 3986 501739
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 3923 471204 3989 471205
rect 3923 471140 3924 471204
rect 3988 471140 3989 471204
rect 3923 471139 3989 471140
rect 3555 467396 3621 467397
rect 3555 467332 3556 467396
rect 3620 467332 3621 467396
rect 3555 467331 3621 467332
rect 3371 456108 3437 456109
rect 3371 456044 3372 456108
rect 3436 456044 3437 456108
rect 3371 456043 3437 456044
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 3371 293180 3437 293181
rect 3371 293116 3372 293180
rect 3436 293116 3437 293180
rect 3371 293115 3437 293116
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 3374 279445 3434 293115
rect 3371 279444 3437 279445
rect 3371 279380 3372 279444
rect 3436 279380 3437 279444
rect 3371 279379 3437 279380
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 3371 254148 3437 254149
rect 3371 254084 3372 254148
rect 3436 254084 3437 254148
rect 3371 254083 3437 254084
rect 3374 240685 3434 254083
rect 3371 240684 3437 240685
rect 3371 240620 3372 240684
rect 3436 240620 3437 240684
rect 3371 240619 3437 240620
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 3555 217292 3621 217293
rect 3555 217228 3556 217292
rect 3620 217228 3621 217292
rect 3555 217227 3621 217228
rect 3371 202196 3437 202197
rect 3371 202132 3372 202196
rect 3436 202132 3437 202196
rect 3371 202131 3437 202132
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 3187 86324 3253 86325
rect 3187 86260 3188 86324
rect 3252 86260 3253 86324
rect 3187 86259 3253 86260
rect 3190 84693 3250 86259
rect 3187 84692 3253 84693
rect 3187 84628 3188 84692
rect 3252 84628 3253 84692
rect 3187 84627 3253 84628
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 3374 19413 3434 202131
rect 3558 58581 3618 217227
rect 3739 215932 3805 215933
rect 3739 215868 3740 215932
rect 3804 215868 3805 215932
rect 3739 215867 3805 215868
rect 3742 201925 3802 215867
rect 3739 201924 3805 201925
rect 3739 201860 3740 201924
rect 3804 201860 3805 201924
rect 3739 201859 3805 201860
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 3555 58580 3621 58581
rect 3555 58516 3556 58580
rect 3620 58516 3621 58580
rect 3555 58515 3621 58516
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 3371 19412 3437 19413
rect 3371 19348 3372 19412
rect 3436 19348 3437 19412
rect 3371 19347 3437 19348
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -7654 6134 -1862
rect 9234 706758 9854 711590
rect 9234 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 9854 706758
rect 9234 706438 9854 706522
rect 9234 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 9854 706438
rect 9234 694894 9854 706202
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 9234 -2266 9854 10338
rect 9234 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 9854 -2266
rect 9234 -2586 9854 -2502
rect 9234 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 9854 -2586
rect 9234 -7654 9854 -2822
rect 12954 707718 13574 711590
rect 12954 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 13574 707718
rect 12954 707398 13574 707482
rect 12954 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 13574 707398
rect 12954 698614 13574 707162
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect 12954 -3226 13574 14058
rect 12954 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 13574 -3226
rect 12954 -3546 13574 -3462
rect 12954 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 13574 -3546
rect 12954 -7654 13574 -3782
rect 16674 708678 17294 711590
rect 16674 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 17294 708678
rect 16674 708358 17294 708442
rect 16674 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 17294 708358
rect 16674 666334 17294 708122
rect 16674 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 17294 666334
rect 16674 666014 17294 666098
rect 16674 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 17294 666014
rect 16674 630334 17294 665778
rect 16674 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 17294 630334
rect 16674 630014 17294 630098
rect 16674 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 17294 630014
rect 16674 594334 17294 629778
rect 16674 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 17294 594334
rect 16674 594014 17294 594098
rect 16674 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 17294 594014
rect 16674 558334 17294 593778
rect 16674 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 17294 558334
rect 16674 558014 17294 558098
rect 16674 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 17294 558014
rect 16674 522334 17294 557778
rect 16674 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 17294 522334
rect 16674 522014 17294 522098
rect 16674 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 17294 522014
rect 16674 486334 17294 521778
rect 16674 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 17294 486334
rect 16674 486014 17294 486098
rect 16674 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 17294 486014
rect 16674 450334 17294 485778
rect 16674 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 17294 450334
rect 16674 450014 17294 450098
rect 16674 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 17294 450014
rect 16674 414334 17294 449778
rect 16674 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 17294 414334
rect 16674 414014 17294 414098
rect 16674 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 17294 414014
rect 16674 378334 17294 413778
rect 16674 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 17294 378334
rect 16674 378014 17294 378098
rect 16674 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 17294 378014
rect 16674 342334 17294 377778
rect 16674 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 17294 342334
rect 16674 342014 17294 342098
rect 16674 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 17294 342014
rect 16674 306334 17294 341778
rect 16674 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 17294 306334
rect 16674 306014 17294 306098
rect 16674 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 17294 306014
rect 16674 270334 17294 305778
rect 16674 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 17294 270334
rect 16674 270014 17294 270098
rect 16674 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 17294 270014
rect 16674 234334 17294 269778
rect 16674 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 17294 234334
rect 16674 234014 17294 234098
rect 16674 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 17294 234014
rect 16674 198334 17294 233778
rect 16674 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 17294 198334
rect 16674 198014 17294 198098
rect 16674 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 17294 198014
rect 16674 162334 17294 197778
rect 16674 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 17294 162334
rect 16674 162014 17294 162098
rect 16674 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 17294 162014
rect 16674 126334 17294 161778
rect 16674 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 17294 126334
rect 16674 126014 17294 126098
rect 16674 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 17294 126014
rect 16674 90334 17294 125778
rect 16674 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 17294 90334
rect 16674 90014 17294 90098
rect 16674 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 17294 90014
rect 16674 54334 17294 89778
rect 16674 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 17294 54334
rect 16674 54014 17294 54098
rect 16674 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 17294 54014
rect 16674 18334 17294 53778
rect 16674 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 17294 18334
rect 16674 18014 17294 18098
rect 16674 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 17294 18014
rect 16674 -4186 17294 17778
rect 16674 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 17294 -4186
rect 16674 -4506 17294 -4422
rect 16674 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 17294 -4506
rect 16674 -7654 17294 -4742
rect 20394 709638 21014 711590
rect 20394 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 21014 709638
rect 20394 709318 21014 709402
rect 20394 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 21014 709318
rect 20394 670054 21014 709082
rect 20394 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 21014 670054
rect 20394 669734 21014 669818
rect 20394 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 21014 669734
rect 20394 634054 21014 669498
rect 20394 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 21014 634054
rect 20394 633734 21014 633818
rect 20394 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 21014 633734
rect 20394 598054 21014 633498
rect 20394 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 21014 598054
rect 20394 597734 21014 597818
rect 20394 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 21014 597734
rect 20394 562054 21014 597498
rect 20394 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 21014 562054
rect 20394 561734 21014 561818
rect 20394 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 21014 561734
rect 20394 526054 21014 561498
rect 20394 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 21014 526054
rect 20394 525734 21014 525818
rect 20394 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 21014 525734
rect 20394 490054 21014 525498
rect 20394 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 21014 490054
rect 20394 489734 21014 489818
rect 20394 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 21014 489734
rect 20394 454054 21014 489498
rect 20394 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 21014 454054
rect 20394 453734 21014 453818
rect 20394 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 21014 453734
rect 20394 418054 21014 453498
rect 20394 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 21014 418054
rect 20394 417734 21014 417818
rect 20394 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 21014 417734
rect 20394 382054 21014 417498
rect 20394 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 21014 382054
rect 20394 381734 21014 381818
rect 20394 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 21014 381734
rect 20394 346054 21014 381498
rect 20394 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 21014 346054
rect 20394 345734 21014 345818
rect 20394 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 21014 345734
rect 20394 310054 21014 345498
rect 20394 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 21014 310054
rect 20394 309734 21014 309818
rect 20394 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 21014 309734
rect 20394 274054 21014 309498
rect 20394 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 21014 274054
rect 20394 273734 21014 273818
rect 20394 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 21014 273734
rect 20394 238054 21014 273498
rect 20394 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 21014 238054
rect 20394 237734 21014 237818
rect 20394 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 21014 237734
rect 20394 202054 21014 237498
rect 20394 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 21014 202054
rect 20394 201734 21014 201818
rect 20394 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 21014 201734
rect 20394 166054 21014 201498
rect 20394 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 21014 166054
rect 20394 165734 21014 165818
rect 20394 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 21014 165734
rect 20394 130054 21014 165498
rect 20394 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 21014 130054
rect 20394 129734 21014 129818
rect 20394 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 21014 129734
rect 20394 94054 21014 129498
rect 20394 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 21014 94054
rect 20394 93734 21014 93818
rect 20394 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 21014 93734
rect 20394 58054 21014 93498
rect 20394 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 21014 58054
rect 20394 57734 21014 57818
rect 20394 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 21014 57734
rect 20394 22054 21014 57498
rect 20394 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 21014 22054
rect 20394 21734 21014 21818
rect 20394 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 21014 21734
rect 20394 -5146 21014 21498
rect 20394 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 21014 -5146
rect 20394 -5466 21014 -5382
rect 20394 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 21014 -5466
rect 20394 -7654 21014 -5702
rect 24114 710598 24734 711590
rect 24114 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 24734 710598
rect 24114 710278 24734 710362
rect 24114 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 24734 710278
rect 24114 673774 24734 710042
rect 24114 673538 24146 673774
rect 24382 673538 24466 673774
rect 24702 673538 24734 673774
rect 24114 673454 24734 673538
rect 24114 673218 24146 673454
rect 24382 673218 24466 673454
rect 24702 673218 24734 673454
rect 24114 637774 24734 673218
rect 24114 637538 24146 637774
rect 24382 637538 24466 637774
rect 24702 637538 24734 637774
rect 24114 637454 24734 637538
rect 24114 637218 24146 637454
rect 24382 637218 24466 637454
rect 24702 637218 24734 637454
rect 24114 601774 24734 637218
rect 24114 601538 24146 601774
rect 24382 601538 24466 601774
rect 24702 601538 24734 601774
rect 24114 601454 24734 601538
rect 24114 601218 24146 601454
rect 24382 601218 24466 601454
rect 24702 601218 24734 601454
rect 24114 565774 24734 601218
rect 24114 565538 24146 565774
rect 24382 565538 24466 565774
rect 24702 565538 24734 565774
rect 24114 565454 24734 565538
rect 24114 565218 24146 565454
rect 24382 565218 24466 565454
rect 24702 565218 24734 565454
rect 24114 529774 24734 565218
rect 24114 529538 24146 529774
rect 24382 529538 24466 529774
rect 24702 529538 24734 529774
rect 24114 529454 24734 529538
rect 24114 529218 24146 529454
rect 24382 529218 24466 529454
rect 24702 529218 24734 529454
rect 24114 493774 24734 529218
rect 24114 493538 24146 493774
rect 24382 493538 24466 493774
rect 24702 493538 24734 493774
rect 24114 493454 24734 493538
rect 24114 493218 24146 493454
rect 24382 493218 24466 493454
rect 24702 493218 24734 493454
rect 24114 457774 24734 493218
rect 24114 457538 24146 457774
rect 24382 457538 24466 457774
rect 24702 457538 24734 457774
rect 24114 457454 24734 457538
rect 24114 457218 24146 457454
rect 24382 457218 24466 457454
rect 24702 457218 24734 457454
rect 24114 421774 24734 457218
rect 24114 421538 24146 421774
rect 24382 421538 24466 421774
rect 24702 421538 24734 421774
rect 24114 421454 24734 421538
rect 24114 421218 24146 421454
rect 24382 421218 24466 421454
rect 24702 421218 24734 421454
rect 24114 385774 24734 421218
rect 24114 385538 24146 385774
rect 24382 385538 24466 385774
rect 24702 385538 24734 385774
rect 24114 385454 24734 385538
rect 24114 385218 24146 385454
rect 24382 385218 24466 385454
rect 24702 385218 24734 385454
rect 24114 349774 24734 385218
rect 24114 349538 24146 349774
rect 24382 349538 24466 349774
rect 24702 349538 24734 349774
rect 24114 349454 24734 349538
rect 24114 349218 24146 349454
rect 24382 349218 24466 349454
rect 24702 349218 24734 349454
rect 24114 313774 24734 349218
rect 24114 313538 24146 313774
rect 24382 313538 24466 313774
rect 24702 313538 24734 313774
rect 24114 313454 24734 313538
rect 24114 313218 24146 313454
rect 24382 313218 24466 313454
rect 24702 313218 24734 313454
rect 24114 277774 24734 313218
rect 24114 277538 24146 277774
rect 24382 277538 24466 277774
rect 24702 277538 24734 277774
rect 24114 277454 24734 277538
rect 24114 277218 24146 277454
rect 24382 277218 24466 277454
rect 24702 277218 24734 277454
rect 24114 241774 24734 277218
rect 24114 241538 24146 241774
rect 24382 241538 24466 241774
rect 24702 241538 24734 241774
rect 24114 241454 24734 241538
rect 24114 241218 24146 241454
rect 24382 241218 24466 241454
rect 24702 241218 24734 241454
rect 24114 205774 24734 241218
rect 24114 205538 24146 205774
rect 24382 205538 24466 205774
rect 24702 205538 24734 205774
rect 24114 205454 24734 205538
rect 24114 205218 24146 205454
rect 24382 205218 24466 205454
rect 24702 205218 24734 205454
rect 24114 169774 24734 205218
rect 24114 169538 24146 169774
rect 24382 169538 24466 169774
rect 24702 169538 24734 169774
rect 24114 169454 24734 169538
rect 24114 169218 24146 169454
rect 24382 169218 24466 169454
rect 24702 169218 24734 169454
rect 24114 133774 24734 169218
rect 24114 133538 24146 133774
rect 24382 133538 24466 133774
rect 24702 133538 24734 133774
rect 24114 133454 24734 133538
rect 24114 133218 24146 133454
rect 24382 133218 24466 133454
rect 24702 133218 24734 133454
rect 24114 97774 24734 133218
rect 24114 97538 24146 97774
rect 24382 97538 24466 97774
rect 24702 97538 24734 97774
rect 24114 97454 24734 97538
rect 24114 97218 24146 97454
rect 24382 97218 24466 97454
rect 24702 97218 24734 97454
rect 24114 61774 24734 97218
rect 24114 61538 24146 61774
rect 24382 61538 24466 61774
rect 24702 61538 24734 61774
rect 24114 61454 24734 61538
rect 24114 61218 24146 61454
rect 24382 61218 24466 61454
rect 24702 61218 24734 61454
rect 24114 25774 24734 61218
rect 24114 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 24734 25774
rect 24114 25454 24734 25538
rect 24114 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 24734 25454
rect 24114 -6106 24734 25218
rect 24114 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 24734 -6106
rect 24114 -6426 24734 -6342
rect 24114 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 24734 -6426
rect 24114 -7654 24734 -6662
rect 27834 711558 28454 711590
rect 27834 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 28454 711558
rect 27834 711238 28454 711322
rect 27834 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 28454 711238
rect 27834 677494 28454 711002
rect 27834 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 28454 677494
rect 27834 677174 28454 677258
rect 27834 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 28454 677174
rect 27834 641494 28454 676938
rect 27834 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 28454 641494
rect 27834 641174 28454 641258
rect 27834 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 28454 641174
rect 27834 605494 28454 640938
rect 27834 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 28454 605494
rect 27834 605174 28454 605258
rect 27834 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 28454 605174
rect 27834 569494 28454 604938
rect 27834 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 28454 569494
rect 27834 569174 28454 569258
rect 27834 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 28454 569174
rect 27834 533494 28454 568938
rect 27834 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 28454 533494
rect 27834 533174 28454 533258
rect 27834 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 28454 533174
rect 27834 497494 28454 532938
rect 27834 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 28454 497494
rect 27834 497174 28454 497258
rect 27834 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 28454 497174
rect 27834 461494 28454 496938
rect 27834 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 28454 461494
rect 27834 461174 28454 461258
rect 27834 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 28454 461174
rect 27834 425494 28454 460938
rect 27834 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 28454 425494
rect 27834 425174 28454 425258
rect 27834 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 28454 425174
rect 27834 389494 28454 424938
rect 27834 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 28454 389494
rect 27834 389174 28454 389258
rect 27834 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 28454 389174
rect 27834 353494 28454 388938
rect 27834 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 28454 353494
rect 27834 353174 28454 353258
rect 27834 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 28454 353174
rect 27834 317494 28454 352938
rect 27834 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 28454 317494
rect 27834 317174 28454 317258
rect 27834 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 28454 317174
rect 27834 281494 28454 316938
rect 27834 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 28454 281494
rect 27834 281174 28454 281258
rect 27834 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 28454 281174
rect 27834 245494 28454 280938
rect 27834 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 28454 245494
rect 27834 245174 28454 245258
rect 27834 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 28454 245174
rect 27834 209494 28454 244938
rect 27834 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 28454 209494
rect 27834 209174 28454 209258
rect 27834 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 28454 209174
rect 27834 173494 28454 208938
rect 27834 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 28454 173494
rect 27834 173174 28454 173258
rect 27834 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 28454 173174
rect 27834 137494 28454 172938
rect 27834 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 28454 137494
rect 27834 137174 28454 137258
rect 27834 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 28454 137174
rect 27834 101494 28454 136938
rect 27834 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 28454 101494
rect 27834 101174 28454 101258
rect 27834 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 28454 101174
rect 27834 65494 28454 100938
rect 27834 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 28454 65494
rect 27834 65174 28454 65258
rect 27834 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 28454 65174
rect 27834 29494 28454 64938
rect 27834 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 28454 29494
rect 27834 29174 28454 29258
rect 27834 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 28454 29174
rect 27834 -7066 28454 28938
rect 27834 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 28454 -7066
rect 27834 -7386 28454 -7302
rect 27834 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 28454 -7386
rect 27834 -7654 28454 -7622
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 41514 705798 42134 711590
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 691174 42134 705242
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -1306 42134 6618
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -7654 42134 -1862
rect 45234 706758 45854 711590
rect 45234 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 45854 706758
rect 45234 706438 45854 706522
rect 45234 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 45854 706438
rect 45234 694894 45854 706202
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 48954 707718 49574 711590
rect 48954 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 49574 707718
rect 48954 707398 49574 707482
rect 48954 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 49574 707398
rect 48954 698614 49574 707162
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48635 306236 48701 306237
rect 48635 306172 48636 306236
rect 48700 306172 48701 306236
rect 48635 306171 48701 306172
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 48638 239869 48698 306171
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48635 239868 48701 239869
rect 48635 239804 48636 239868
rect 48700 239804 48701 239868
rect 48635 239803 48701 239804
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -2266 45854 10338
rect 45234 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 45854 -2266
rect 45234 -2586 45854 -2502
rect 45234 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 45854 -2586
rect 45234 -7654 45854 -2822
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 48954 -3226 49574 14058
rect 48954 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 49574 -3226
rect 48954 -3546 49574 -3462
rect 48954 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 49574 -3546
rect 48954 -7654 49574 -3782
rect 52674 708678 53294 711590
rect 52674 708442 52706 708678
rect 52942 708442 53026 708678
rect 53262 708442 53294 708678
rect 52674 708358 53294 708442
rect 52674 708122 52706 708358
rect 52942 708122 53026 708358
rect 53262 708122 53294 708358
rect 52674 666334 53294 708122
rect 52674 666098 52706 666334
rect 52942 666098 53026 666334
rect 53262 666098 53294 666334
rect 52674 666014 53294 666098
rect 52674 665778 52706 666014
rect 52942 665778 53026 666014
rect 53262 665778 53294 666014
rect 52674 630334 53294 665778
rect 52674 630098 52706 630334
rect 52942 630098 53026 630334
rect 53262 630098 53294 630334
rect 52674 630014 53294 630098
rect 52674 629778 52706 630014
rect 52942 629778 53026 630014
rect 53262 629778 53294 630014
rect 52674 594334 53294 629778
rect 52674 594098 52706 594334
rect 52942 594098 53026 594334
rect 53262 594098 53294 594334
rect 52674 594014 53294 594098
rect 52674 593778 52706 594014
rect 52942 593778 53026 594014
rect 53262 593778 53294 594014
rect 52674 558334 53294 593778
rect 52674 558098 52706 558334
rect 52942 558098 53026 558334
rect 53262 558098 53294 558334
rect 52674 558014 53294 558098
rect 52674 557778 52706 558014
rect 52942 557778 53026 558014
rect 53262 557778 53294 558014
rect 52674 522334 53294 557778
rect 52674 522098 52706 522334
rect 52942 522098 53026 522334
rect 53262 522098 53294 522334
rect 52674 522014 53294 522098
rect 52674 521778 52706 522014
rect 52942 521778 53026 522014
rect 53262 521778 53294 522014
rect 52674 486334 53294 521778
rect 52674 486098 52706 486334
rect 52942 486098 53026 486334
rect 53262 486098 53294 486334
rect 52674 486014 53294 486098
rect 52674 485778 52706 486014
rect 52942 485778 53026 486014
rect 53262 485778 53294 486014
rect 52674 450334 53294 485778
rect 52674 450098 52706 450334
rect 52942 450098 53026 450334
rect 53262 450098 53294 450334
rect 52674 450014 53294 450098
rect 52674 449778 52706 450014
rect 52942 449778 53026 450014
rect 53262 449778 53294 450014
rect 52674 414334 53294 449778
rect 52674 414098 52706 414334
rect 52942 414098 53026 414334
rect 53262 414098 53294 414334
rect 52674 414014 53294 414098
rect 52674 413778 52706 414014
rect 52942 413778 53026 414014
rect 53262 413778 53294 414014
rect 52674 378334 53294 413778
rect 52674 378098 52706 378334
rect 52942 378098 53026 378334
rect 53262 378098 53294 378334
rect 52674 378014 53294 378098
rect 52674 377778 52706 378014
rect 52942 377778 53026 378014
rect 53262 377778 53294 378014
rect 52674 342334 53294 377778
rect 52674 342098 52706 342334
rect 52942 342098 53026 342334
rect 53262 342098 53294 342334
rect 52674 342014 53294 342098
rect 52674 341778 52706 342014
rect 52942 341778 53026 342014
rect 53262 341778 53294 342014
rect 52674 306334 53294 341778
rect 56394 709638 57014 711590
rect 56394 709402 56426 709638
rect 56662 709402 56746 709638
rect 56982 709402 57014 709638
rect 56394 709318 57014 709402
rect 56394 709082 56426 709318
rect 56662 709082 56746 709318
rect 56982 709082 57014 709318
rect 56394 670054 57014 709082
rect 60114 710598 60734 711590
rect 60114 710362 60146 710598
rect 60382 710362 60466 710598
rect 60702 710362 60734 710598
rect 60114 710278 60734 710362
rect 60114 710042 60146 710278
rect 60382 710042 60466 710278
rect 60702 710042 60734 710278
rect 60114 673774 60734 710042
rect 60114 673538 60146 673774
rect 60382 673538 60466 673774
rect 60702 673538 60734 673774
rect 60114 673454 60734 673538
rect 60114 673218 60146 673454
rect 60382 673218 60466 673454
rect 60702 673218 60734 673454
rect 57283 671260 57349 671261
rect 57283 671196 57284 671260
rect 57348 671196 57349 671260
rect 57283 671195 57349 671196
rect 56394 669818 56426 670054
rect 56662 669818 56746 670054
rect 56982 669818 57014 670054
rect 56394 669734 57014 669818
rect 56394 669498 56426 669734
rect 56662 669498 56746 669734
rect 56982 669498 57014 669734
rect 56394 634054 57014 669498
rect 56394 633818 56426 634054
rect 56662 633818 56746 634054
rect 56982 633818 57014 634054
rect 56394 633734 57014 633818
rect 56394 633498 56426 633734
rect 56662 633498 56746 633734
rect 56982 633498 57014 633734
rect 56394 598054 57014 633498
rect 56394 597818 56426 598054
rect 56662 597818 56746 598054
rect 56982 597818 57014 598054
rect 56394 597734 57014 597818
rect 56394 597498 56426 597734
rect 56662 597498 56746 597734
rect 56982 597498 57014 597734
rect 56394 562054 57014 597498
rect 56394 561818 56426 562054
rect 56662 561818 56746 562054
rect 56982 561818 57014 562054
rect 56394 561734 57014 561818
rect 56394 561498 56426 561734
rect 56662 561498 56746 561734
rect 56982 561498 57014 561734
rect 56394 526054 57014 561498
rect 56394 525818 56426 526054
rect 56662 525818 56746 526054
rect 56982 525818 57014 526054
rect 56394 525734 57014 525818
rect 56394 525498 56426 525734
rect 56662 525498 56746 525734
rect 56982 525498 57014 525734
rect 56394 490054 57014 525498
rect 56394 489818 56426 490054
rect 56662 489818 56746 490054
rect 56982 489818 57014 490054
rect 56394 489734 57014 489818
rect 56394 489498 56426 489734
rect 56662 489498 56746 489734
rect 56982 489498 57014 489734
rect 56394 454054 57014 489498
rect 56394 453818 56426 454054
rect 56662 453818 56746 454054
rect 56982 453818 57014 454054
rect 56394 453734 57014 453818
rect 56394 453498 56426 453734
rect 56662 453498 56746 453734
rect 56982 453498 57014 453734
rect 56394 418054 57014 453498
rect 57286 444277 57346 671195
rect 60114 637774 60734 673218
rect 60114 637538 60146 637774
rect 60382 637538 60466 637774
rect 60702 637538 60734 637774
rect 60114 637454 60734 637538
rect 60114 637218 60146 637454
rect 60382 637218 60466 637454
rect 60702 637218 60734 637454
rect 60114 601774 60734 637218
rect 60114 601538 60146 601774
rect 60382 601538 60466 601774
rect 60702 601538 60734 601774
rect 60114 601454 60734 601538
rect 60114 601218 60146 601454
rect 60382 601218 60466 601454
rect 60702 601218 60734 601454
rect 60114 565774 60734 601218
rect 63834 711558 64454 711590
rect 63834 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 64454 711558
rect 63834 711238 64454 711322
rect 63834 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 64454 711238
rect 63834 677494 64454 711002
rect 63834 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 64454 677494
rect 63834 677174 64454 677258
rect 63834 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 64454 677174
rect 63834 641494 64454 676938
rect 63834 641258 63866 641494
rect 64102 641258 64186 641494
rect 64422 641258 64454 641494
rect 63834 641174 64454 641258
rect 63834 640938 63866 641174
rect 64102 640938 64186 641174
rect 64422 640938 64454 641174
rect 63834 605494 64454 640938
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 629612 74414 650898
rect 77514 705798 78134 711590
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 691174 78134 705242
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 629257 78134 654618
rect 81234 706758 81854 711590
rect 81234 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 81854 706758
rect 81234 706438 81854 706522
rect 81234 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 81854 706438
rect 81234 694894 81854 706202
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 629257 81854 658338
rect 84954 707718 85574 711590
rect 84954 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 85574 707718
rect 84954 707398 85574 707482
rect 84954 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 85574 707398
rect 84954 698614 85574 707162
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 629257 85574 662058
rect 88674 708678 89294 711590
rect 88674 708442 88706 708678
rect 88942 708442 89026 708678
rect 89262 708442 89294 708678
rect 88674 708358 89294 708442
rect 88674 708122 88706 708358
rect 88942 708122 89026 708358
rect 89262 708122 89294 708358
rect 88674 666334 89294 708122
rect 88674 666098 88706 666334
rect 88942 666098 89026 666334
rect 89262 666098 89294 666334
rect 88674 666014 89294 666098
rect 88674 665778 88706 666014
rect 88942 665778 89026 666014
rect 89262 665778 89294 666014
rect 88674 630334 89294 665778
rect 88674 630098 88706 630334
rect 88942 630098 89026 630334
rect 89262 630098 89294 630334
rect 88674 630014 89294 630098
rect 88674 629778 88706 630014
rect 88942 629778 89026 630014
rect 89262 629778 89294 630014
rect 88674 629257 89294 629778
rect 92394 709638 93014 711590
rect 92394 709402 92426 709638
rect 92662 709402 92746 709638
rect 92982 709402 93014 709638
rect 92394 709318 93014 709402
rect 92394 709082 92426 709318
rect 92662 709082 92746 709318
rect 92982 709082 93014 709318
rect 92394 670054 93014 709082
rect 92394 669818 92426 670054
rect 92662 669818 92746 670054
rect 92982 669818 93014 670054
rect 92394 669734 93014 669818
rect 92394 669498 92426 669734
rect 92662 669498 92746 669734
rect 92982 669498 93014 669734
rect 92394 634054 93014 669498
rect 92394 633818 92426 634054
rect 92662 633818 92746 634054
rect 92982 633818 93014 634054
rect 92394 633734 93014 633818
rect 92394 633498 92426 633734
rect 92662 633498 92746 633734
rect 92982 633498 93014 633734
rect 92394 629257 93014 633498
rect 96114 710598 96734 711590
rect 96114 710362 96146 710598
rect 96382 710362 96466 710598
rect 96702 710362 96734 710598
rect 96114 710278 96734 710362
rect 96114 710042 96146 710278
rect 96382 710042 96466 710278
rect 96702 710042 96734 710278
rect 96114 673774 96734 710042
rect 96114 673538 96146 673774
rect 96382 673538 96466 673774
rect 96702 673538 96734 673774
rect 96114 673454 96734 673538
rect 96114 673218 96146 673454
rect 96382 673218 96466 673454
rect 96702 673218 96734 673454
rect 96114 637774 96734 673218
rect 96114 637538 96146 637774
rect 96382 637538 96466 637774
rect 96702 637538 96734 637774
rect 96114 637454 96734 637538
rect 96114 637218 96146 637454
rect 96382 637218 96466 637454
rect 96702 637218 96734 637454
rect 96114 629257 96734 637218
rect 99834 711558 100454 711590
rect 99834 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 100454 711558
rect 99834 711238 100454 711322
rect 99834 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 100454 711238
rect 99834 677494 100454 711002
rect 99834 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 100454 677494
rect 99834 677174 100454 677258
rect 99834 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 100454 677174
rect 99834 641494 100454 676938
rect 99834 641258 99866 641494
rect 100102 641258 100186 641494
rect 100422 641258 100454 641494
rect 99834 641174 100454 641258
rect 99834 640938 99866 641174
rect 100102 640938 100186 641174
rect 100422 640938 100454 641174
rect 99834 629257 100454 640938
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 629257 110414 650898
rect 113514 705798 114134 711590
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 691174 114134 705242
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 629257 114134 654618
rect 117234 706758 117854 711590
rect 117234 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 117854 706758
rect 117234 706438 117854 706522
rect 117234 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 117854 706438
rect 117234 694894 117854 706202
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 629257 117854 658338
rect 120954 707718 121574 711590
rect 120954 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 121574 707718
rect 120954 707398 121574 707482
rect 120954 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 121574 707398
rect 120954 698614 121574 707162
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 629257 121574 662058
rect 124674 708678 125294 711590
rect 124674 708442 124706 708678
rect 124942 708442 125026 708678
rect 125262 708442 125294 708678
rect 124674 708358 125294 708442
rect 124674 708122 124706 708358
rect 124942 708122 125026 708358
rect 125262 708122 125294 708358
rect 124674 666334 125294 708122
rect 124674 666098 124706 666334
rect 124942 666098 125026 666334
rect 125262 666098 125294 666334
rect 124674 666014 125294 666098
rect 124674 665778 124706 666014
rect 124942 665778 125026 666014
rect 125262 665778 125294 666014
rect 124674 630334 125294 665778
rect 124674 630098 124706 630334
rect 124942 630098 125026 630334
rect 125262 630098 125294 630334
rect 124674 630014 125294 630098
rect 124674 629778 124706 630014
rect 124942 629778 125026 630014
rect 125262 629778 125294 630014
rect 124674 629257 125294 629778
rect 128394 709638 129014 711590
rect 128394 709402 128426 709638
rect 128662 709402 128746 709638
rect 128982 709402 129014 709638
rect 128394 709318 129014 709402
rect 128394 709082 128426 709318
rect 128662 709082 128746 709318
rect 128982 709082 129014 709318
rect 128394 670054 129014 709082
rect 128394 669818 128426 670054
rect 128662 669818 128746 670054
rect 128982 669818 129014 670054
rect 128394 669734 129014 669818
rect 128394 669498 128426 669734
rect 128662 669498 128746 669734
rect 128982 669498 129014 669734
rect 128394 634054 129014 669498
rect 128394 633818 128426 634054
rect 128662 633818 128746 634054
rect 128982 633818 129014 634054
rect 128394 633734 129014 633818
rect 128394 633498 128426 633734
rect 128662 633498 128746 633734
rect 128982 633498 129014 633734
rect 128394 629257 129014 633498
rect 132114 710598 132734 711590
rect 132114 710362 132146 710598
rect 132382 710362 132466 710598
rect 132702 710362 132734 710598
rect 132114 710278 132734 710362
rect 132114 710042 132146 710278
rect 132382 710042 132466 710278
rect 132702 710042 132734 710278
rect 132114 673774 132734 710042
rect 132114 673538 132146 673774
rect 132382 673538 132466 673774
rect 132702 673538 132734 673774
rect 132114 673454 132734 673538
rect 132114 673218 132146 673454
rect 132382 673218 132466 673454
rect 132702 673218 132734 673454
rect 132114 637774 132734 673218
rect 132114 637538 132146 637774
rect 132382 637538 132466 637774
rect 132702 637538 132734 637774
rect 132114 637454 132734 637538
rect 132114 637218 132146 637454
rect 132382 637218 132466 637454
rect 132702 637218 132734 637454
rect 132114 629257 132734 637218
rect 135834 711558 136454 711590
rect 135834 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 136454 711558
rect 135834 711238 136454 711322
rect 135834 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 136454 711238
rect 135834 677494 136454 711002
rect 135834 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 136454 677494
rect 135834 677174 136454 677258
rect 135834 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 136454 677174
rect 135834 641494 136454 676938
rect 135834 641258 135866 641494
rect 136102 641258 136186 641494
rect 136422 641258 136454 641494
rect 135834 641174 136454 641258
rect 135834 640938 135866 641174
rect 136102 640938 136186 641174
rect 136422 640938 136454 641174
rect 135834 629612 136454 640938
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 629257 146414 650898
rect 149514 705798 150134 711590
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 691174 150134 705242
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 629257 150134 654618
rect 153234 706758 153854 711590
rect 153234 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 153854 706758
rect 153234 706438 153854 706522
rect 153234 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 153854 706438
rect 153234 694894 153854 706202
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 629257 153854 658338
rect 156954 707718 157574 711590
rect 156954 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 157574 707718
rect 156954 707398 157574 707482
rect 156954 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 157574 707398
rect 156954 698614 157574 707162
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 629257 157574 662058
rect 160674 708678 161294 711590
rect 160674 708442 160706 708678
rect 160942 708442 161026 708678
rect 161262 708442 161294 708678
rect 160674 708358 161294 708442
rect 160674 708122 160706 708358
rect 160942 708122 161026 708358
rect 161262 708122 161294 708358
rect 160674 666334 161294 708122
rect 160674 666098 160706 666334
rect 160942 666098 161026 666334
rect 161262 666098 161294 666334
rect 160674 666014 161294 666098
rect 160674 665778 160706 666014
rect 160942 665778 161026 666014
rect 161262 665778 161294 666014
rect 160674 630334 161294 665778
rect 160674 630098 160706 630334
rect 160942 630098 161026 630334
rect 161262 630098 161294 630334
rect 160674 630014 161294 630098
rect 160674 629778 160706 630014
rect 160942 629778 161026 630014
rect 161262 629778 161294 630014
rect 160674 629257 161294 629778
rect 164394 709638 165014 711590
rect 164394 709402 164426 709638
rect 164662 709402 164746 709638
rect 164982 709402 165014 709638
rect 164394 709318 165014 709402
rect 164394 709082 164426 709318
rect 164662 709082 164746 709318
rect 164982 709082 165014 709318
rect 164394 670054 165014 709082
rect 164394 669818 164426 670054
rect 164662 669818 164746 670054
rect 164982 669818 165014 670054
rect 164394 669734 165014 669818
rect 164394 669498 164426 669734
rect 164662 669498 164746 669734
rect 164982 669498 165014 669734
rect 164394 634054 165014 669498
rect 164394 633818 164426 634054
rect 164662 633818 164746 634054
rect 164982 633818 165014 634054
rect 164394 633734 165014 633818
rect 164394 633498 164426 633734
rect 164662 633498 164746 633734
rect 164982 633498 165014 633734
rect 164394 629257 165014 633498
rect 168114 710598 168734 711590
rect 168114 710362 168146 710598
rect 168382 710362 168466 710598
rect 168702 710362 168734 710598
rect 168114 710278 168734 710362
rect 168114 710042 168146 710278
rect 168382 710042 168466 710278
rect 168702 710042 168734 710278
rect 168114 673774 168734 710042
rect 168114 673538 168146 673774
rect 168382 673538 168466 673774
rect 168702 673538 168734 673774
rect 168114 673454 168734 673538
rect 168114 673218 168146 673454
rect 168382 673218 168466 673454
rect 168702 673218 168734 673454
rect 168114 637774 168734 673218
rect 168114 637538 168146 637774
rect 168382 637538 168466 637774
rect 168702 637538 168734 637774
rect 168114 637454 168734 637538
rect 168114 637218 168146 637454
rect 168382 637218 168466 637454
rect 168702 637218 168734 637454
rect 168114 629257 168734 637218
rect 171834 711558 172454 711590
rect 171834 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 172454 711558
rect 171834 711238 172454 711322
rect 171834 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 172454 711238
rect 171834 677494 172454 711002
rect 171834 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 172454 677494
rect 171834 677174 172454 677258
rect 171834 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 172454 677174
rect 171834 641494 172454 676938
rect 171834 641258 171866 641494
rect 172102 641258 172186 641494
rect 172422 641258 172454 641494
rect 171834 641174 172454 641258
rect 171834 640938 171866 641174
rect 172102 640938 172186 641174
rect 172422 640938 172454 641174
rect 171834 629257 172454 640938
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 629612 182414 650898
rect 185514 705798 186134 711590
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 691174 186134 705242
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 629257 186134 654618
rect 189234 706758 189854 711590
rect 189234 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 189854 706758
rect 189234 706438 189854 706522
rect 189234 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 189854 706438
rect 189234 694894 189854 706202
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 629257 189854 658338
rect 192954 707718 193574 711590
rect 192954 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 193574 707718
rect 192954 707398 193574 707482
rect 192954 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 193574 707398
rect 192954 698614 193574 707162
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 629257 193574 662058
rect 196674 708678 197294 711590
rect 196674 708442 196706 708678
rect 196942 708442 197026 708678
rect 197262 708442 197294 708678
rect 196674 708358 197294 708442
rect 196674 708122 196706 708358
rect 196942 708122 197026 708358
rect 197262 708122 197294 708358
rect 196674 666334 197294 708122
rect 196674 666098 196706 666334
rect 196942 666098 197026 666334
rect 197262 666098 197294 666334
rect 196674 666014 197294 666098
rect 196674 665778 196706 666014
rect 196942 665778 197026 666014
rect 197262 665778 197294 666014
rect 196674 630334 197294 665778
rect 196674 630098 196706 630334
rect 196942 630098 197026 630334
rect 197262 630098 197294 630334
rect 196674 630014 197294 630098
rect 196674 629778 196706 630014
rect 196942 629778 197026 630014
rect 197262 629778 197294 630014
rect 196674 629612 197294 629778
rect 200394 709638 201014 711590
rect 200394 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 201014 709638
rect 200394 709318 201014 709402
rect 200394 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 201014 709318
rect 200394 670054 201014 709082
rect 200394 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 201014 670054
rect 200394 669734 201014 669818
rect 200394 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 201014 669734
rect 200394 634054 201014 669498
rect 200394 633818 200426 634054
rect 200662 633818 200746 634054
rect 200982 633818 201014 634054
rect 200394 633734 201014 633818
rect 200394 633498 200426 633734
rect 200662 633498 200746 633734
rect 200982 633498 201014 633734
rect 200394 629257 201014 633498
rect 204114 710598 204734 711590
rect 204114 710362 204146 710598
rect 204382 710362 204466 710598
rect 204702 710362 204734 710598
rect 204114 710278 204734 710362
rect 204114 710042 204146 710278
rect 204382 710042 204466 710278
rect 204702 710042 204734 710278
rect 204114 673774 204734 710042
rect 204114 673538 204146 673774
rect 204382 673538 204466 673774
rect 204702 673538 204734 673774
rect 204114 673454 204734 673538
rect 204114 673218 204146 673454
rect 204382 673218 204466 673454
rect 204702 673218 204734 673454
rect 204114 637774 204734 673218
rect 204114 637538 204146 637774
rect 204382 637538 204466 637774
rect 204702 637538 204734 637774
rect 204114 637454 204734 637538
rect 204114 637218 204146 637454
rect 204382 637218 204466 637454
rect 204702 637218 204734 637454
rect 204114 629257 204734 637218
rect 207834 711558 208454 711590
rect 207834 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 208454 711558
rect 207834 711238 208454 711322
rect 207834 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 208454 711238
rect 207834 677494 208454 711002
rect 207834 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 208454 677494
rect 207834 677174 208454 677258
rect 207834 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 208454 677174
rect 207834 641494 208454 676938
rect 207834 641258 207866 641494
rect 208102 641258 208186 641494
rect 208422 641258 208454 641494
rect 207834 641174 208454 641258
rect 207834 640938 207866 641174
rect 208102 640938 208186 641174
rect 208422 640938 208454 641174
rect 207834 629257 208454 640938
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 629257 218414 650898
rect 221514 705798 222134 711590
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 691174 222134 705242
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 629257 222134 654618
rect 225234 706758 225854 711590
rect 225234 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 225854 706758
rect 225234 706438 225854 706522
rect 225234 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 225854 706438
rect 225234 694894 225854 706202
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 629257 225854 658338
rect 228954 707718 229574 711590
rect 228954 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 229574 707718
rect 228954 707398 229574 707482
rect 228954 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 229574 707398
rect 228954 698614 229574 707162
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 629257 229574 662058
rect 232674 708678 233294 711590
rect 232674 708442 232706 708678
rect 232942 708442 233026 708678
rect 233262 708442 233294 708678
rect 232674 708358 233294 708442
rect 232674 708122 232706 708358
rect 232942 708122 233026 708358
rect 233262 708122 233294 708358
rect 232674 666334 233294 708122
rect 232674 666098 232706 666334
rect 232942 666098 233026 666334
rect 233262 666098 233294 666334
rect 232674 666014 233294 666098
rect 232674 665778 232706 666014
rect 232942 665778 233026 666014
rect 233262 665778 233294 666014
rect 232674 630334 233294 665778
rect 232674 630098 232706 630334
rect 232942 630098 233026 630334
rect 233262 630098 233294 630334
rect 232674 630014 233294 630098
rect 232674 629778 232706 630014
rect 232942 629778 233026 630014
rect 233262 629778 233294 630014
rect 232674 629257 233294 629778
rect 236394 709638 237014 711590
rect 236394 709402 236426 709638
rect 236662 709402 236746 709638
rect 236982 709402 237014 709638
rect 236394 709318 237014 709402
rect 236394 709082 236426 709318
rect 236662 709082 236746 709318
rect 236982 709082 237014 709318
rect 236394 670054 237014 709082
rect 236394 669818 236426 670054
rect 236662 669818 236746 670054
rect 236982 669818 237014 670054
rect 236394 669734 237014 669818
rect 236394 669498 236426 669734
rect 236662 669498 236746 669734
rect 236982 669498 237014 669734
rect 236394 634054 237014 669498
rect 236394 633818 236426 634054
rect 236662 633818 236746 634054
rect 236982 633818 237014 634054
rect 236394 633734 237014 633818
rect 236394 633498 236426 633734
rect 236662 633498 236746 633734
rect 236982 633498 237014 633734
rect 236394 629257 237014 633498
rect 240114 710598 240734 711590
rect 240114 710362 240146 710598
rect 240382 710362 240466 710598
rect 240702 710362 240734 710598
rect 240114 710278 240734 710362
rect 240114 710042 240146 710278
rect 240382 710042 240466 710278
rect 240702 710042 240734 710278
rect 240114 673774 240734 710042
rect 240114 673538 240146 673774
rect 240382 673538 240466 673774
rect 240702 673538 240734 673774
rect 240114 673454 240734 673538
rect 240114 673218 240146 673454
rect 240382 673218 240466 673454
rect 240702 673218 240734 673454
rect 240114 637774 240734 673218
rect 240114 637538 240146 637774
rect 240382 637538 240466 637774
rect 240702 637538 240734 637774
rect 240114 637454 240734 637538
rect 240114 637218 240146 637454
rect 240382 637218 240466 637454
rect 240702 637218 240734 637454
rect 240114 629257 240734 637218
rect 243834 711558 244454 711590
rect 243834 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 244454 711558
rect 243834 711238 244454 711322
rect 243834 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 244454 711238
rect 243834 677494 244454 711002
rect 243834 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 244454 677494
rect 243834 677174 244454 677258
rect 243834 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 244454 677174
rect 243834 641494 244454 676938
rect 243834 641258 243866 641494
rect 244102 641258 244186 641494
rect 244422 641258 244454 641494
rect 243834 641174 244454 641258
rect 243834 640938 243866 641174
rect 244102 640938 244186 641174
rect 244422 640938 244454 641174
rect 243834 629257 244454 640938
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 629257 254414 650898
rect 257514 705798 258134 711590
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 691174 258134 705242
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 629257 258134 654618
rect 261234 706758 261854 711590
rect 261234 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 261854 706758
rect 261234 706438 261854 706522
rect 261234 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 261854 706438
rect 261234 694894 261854 706202
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 629257 261854 658338
rect 264954 707718 265574 711590
rect 264954 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 265574 707718
rect 264954 707398 265574 707482
rect 264954 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 265574 707398
rect 264954 698614 265574 707162
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 629257 265574 662058
rect 268674 708678 269294 711590
rect 268674 708442 268706 708678
rect 268942 708442 269026 708678
rect 269262 708442 269294 708678
rect 268674 708358 269294 708442
rect 268674 708122 268706 708358
rect 268942 708122 269026 708358
rect 269262 708122 269294 708358
rect 268674 666334 269294 708122
rect 268674 666098 268706 666334
rect 268942 666098 269026 666334
rect 269262 666098 269294 666334
rect 268674 666014 269294 666098
rect 268674 665778 268706 666014
rect 268942 665778 269026 666014
rect 269262 665778 269294 666014
rect 268674 630334 269294 665778
rect 268674 630098 268706 630334
rect 268942 630098 269026 630334
rect 269262 630098 269294 630334
rect 268674 630014 269294 630098
rect 268674 629778 268706 630014
rect 268942 629778 269026 630014
rect 269262 629778 269294 630014
rect 268674 629257 269294 629778
rect 272394 709638 273014 711590
rect 272394 709402 272426 709638
rect 272662 709402 272746 709638
rect 272982 709402 273014 709638
rect 272394 709318 273014 709402
rect 272394 709082 272426 709318
rect 272662 709082 272746 709318
rect 272982 709082 273014 709318
rect 272394 670054 273014 709082
rect 272394 669818 272426 670054
rect 272662 669818 272746 670054
rect 272982 669818 273014 670054
rect 272394 669734 273014 669818
rect 272394 669498 272426 669734
rect 272662 669498 272746 669734
rect 272982 669498 273014 669734
rect 272394 634054 273014 669498
rect 272394 633818 272426 634054
rect 272662 633818 272746 634054
rect 272982 633818 273014 634054
rect 272394 633734 273014 633818
rect 272394 633498 272426 633734
rect 272662 633498 272746 633734
rect 272982 633498 273014 633734
rect 272394 629257 273014 633498
rect 276114 710598 276734 711590
rect 276114 710362 276146 710598
rect 276382 710362 276466 710598
rect 276702 710362 276734 710598
rect 276114 710278 276734 710362
rect 276114 710042 276146 710278
rect 276382 710042 276466 710278
rect 276702 710042 276734 710278
rect 276114 673774 276734 710042
rect 276114 673538 276146 673774
rect 276382 673538 276466 673774
rect 276702 673538 276734 673774
rect 276114 673454 276734 673538
rect 276114 673218 276146 673454
rect 276382 673218 276466 673454
rect 276702 673218 276734 673454
rect 276114 637774 276734 673218
rect 276114 637538 276146 637774
rect 276382 637538 276466 637774
rect 276702 637538 276734 637774
rect 276114 637454 276734 637538
rect 276114 637218 276146 637454
rect 276382 637218 276466 637454
rect 276702 637218 276734 637454
rect 276114 629257 276734 637218
rect 279834 711558 280454 711590
rect 279834 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 280454 711558
rect 279834 711238 280454 711322
rect 279834 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 280454 711238
rect 279834 677494 280454 711002
rect 279834 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 280454 677494
rect 279834 677174 280454 677258
rect 279834 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 280454 677174
rect 279834 641494 280454 676938
rect 279834 641258 279866 641494
rect 280102 641258 280186 641494
rect 280422 641258 280454 641494
rect 279834 641174 280454 641258
rect 279834 640938 279866 641174
rect 280102 640938 280186 641174
rect 280422 640938 280454 641174
rect 279834 629257 280454 640938
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 68507 626652 68573 626653
rect 68507 626588 68508 626652
rect 68572 626588 68573 626652
rect 68507 626587 68573 626588
rect 68139 609244 68205 609245
rect 68139 609180 68140 609244
rect 68204 609180 68205 609244
rect 68139 609179 68205 609180
rect 63834 605258 63866 605494
rect 64102 605258 64186 605494
rect 64422 605258 64454 605494
rect 63834 605174 64454 605258
rect 63834 604938 63866 605174
rect 64102 604938 64186 605174
rect 64422 604938 64454 605174
rect 63355 591836 63421 591837
rect 63355 591772 63356 591836
rect 63420 591772 63421 591836
rect 63355 591771 63421 591772
rect 63171 587484 63237 587485
rect 63171 587420 63172 587484
rect 63236 587420 63237 587484
rect 63171 587419 63237 587420
rect 60114 565538 60146 565774
rect 60382 565538 60466 565774
rect 60702 565538 60734 565774
rect 60114 565454 60734 565538
rect 60114 565218 60146 565454
rect 60382 565218 60466 565454
rect 60702 565218 60734 565454
rect 60114 529774 60734 565218
rect 60114 529538 60146 529774
rect 60382 529538 60466 529774
rect 60702 529538 60734 529774
rect 60114 529454 60734 529538
rect 60114 529218 60146 529454
rect 60382 529218 60466 529454
rect 60702 529218 60734 529454
rect 59859 514860 59925 514861
rect 59859 514796 59860 514860
rect 59924 514796 59925 514860
rect 59859 514795 59925 514796
rect 57283 444276 57349 444277
rect 57283 444212 57284 444276
rect 57348 444212 57349 444276
rect 57283 444211 57349 444212
rect 59862 444005 59922 514795
rect 60114 493774 60734 529218
rect 62987 504796 63053 504797
rect 62987 504732 62988 504796
rect 63052 504732 63053 504796
rect 62987 504731 63053 504732
rect 60114 493538 60146 493774
rect 60382 493538 60466 493774
rect 60702 493538 60734 493774
rect 60114 493454 60734 493538
rect 60114 493218 60146 493454
rect 60382 493218 60466 493454
rect 60702 493218 60734 493454
rect 60114 457774 60734 493218
rect 60114 457538 60146 457774
rect 60382 457538 60466 457774
rect 60702 457538 60734 457774
rect 60114 457454 60734 457538
rect 60114 457218 60146 457454
rect 60382 457218 60466 457454
rect 60702 457218 60734 457454
rect 59859 444004 59925 444005
rect 59859 443940 59860 444004
rect 59924 443940 59925 444004
rect 59859 443939 59925 443940
rect 56394 417818 56426 418054
rect 56662 417818 56746 418054
rect 56982 417818 57014 418054
rect 56394 417734 57014 417818
rect 56394 417498 56426 417734
rect 56662 417498 56746 417734
rect 56982 417498 57014 417734
rect 56394 382054 57014 417498
rect 56394 381818 56426 382054
rect 56662 381818 56746 382054
rect 56982 381818 57014 382054
rect 56394 381734 57014 381818
rect 56394 381498 56426 381734
rect 56662 381498 56746 381734
rect 56982 381498 57014 381734
rect 56394 346054 57014 381498
rect 56394 345818 56426 346054
rect 56662 345818 56746 346054
rect 56982 345818 57014 346054
rect 56394 345734 57014 345818
rect 56394 345498 56426 345734
rect 56662 345498 56746 345734
rect 56982 345498 57014 345734
rect 54208 327454 54528 327486
rect 54208 327218 54250 327454
rect 54486 327218 54528 327454
rect 54208 327134 54528 327218
rect 54208 326898 54250 327134
rect 54486 326898 54528 327134
rect 54208 326866 54528 326898
rect 52674 306098 52706 306334
rect 52942 306098 53026 306334
rect 53262 306098 53294 306334
rect 52674 306014 53294 306098
rect 52674 305778 52706 306014
rect 52942 305778 53026 306014
rect 53262 305778 53294 306014
rect 52674 270334 53294 305778
rect 56394 310054 57014 345498
rect 60114 421774 60734 457218
rect 60114 421538 60146 421774
rect 60382 421538 60466 421774
rect 60702 421538 60734 421774
rect 60114 421454 60734 421538
rect 60114 421218 60146 421454
rect 60382 421218 60466 421454
rect 60702 421218 60734 421454
rect 60114 385774 60734 421218
rect 60114 385538 60146 385774
rect 60382 385538 60466 385774
rect 60702 385538 60734 385774
rect 60114 385454 60734 385538
rect 60114 385218 60146 385454
rect 60382 385218 60466 385454
rect 60702 385218 60734 385454
rect 60114 349774 60734 385218
rect 60114 349538 60146 349774
rect 60382 349538 60466 349774
rect 60702 349538 60734 349774
rect 60114 349454 60734 349538
rect 60114 349218 60146 349454
rect 60382 349218 60466 349454
rect 60702 349218 60734 349454
rect 60114 340449 60734 349218
rect 62990 344725 63050 504731
rect 62987 344724 63053 344725
rect 62987 344660 62988 344724
rect 63052 344660 63053 344724
rect 62987 344659 63053 344660
rect 63174 344453 63234 587419
rect 63171 344452 63237 344453
rect 63171 344388 63172 344452
rect 63236 344388 63237 344452
rect 63171 344387 63237 344388
rect 63358 344045 63418 591771
rect 63834 569494 64454 604938
rect 66851 574428 66917 574429
rect 66851 574364 66852 574428
rect 66916 574364 66917 574428
rect 66851 574363 66917 574364
rect 63834 569258 63866 569494
rect 64102 569258 64186 569494
rect 64422 569258 64454 569494
rect 63834 569174 64454 569258
rect 63834 568938 63866 569174
rect 64102 568938 64186 569174
rect 64422 568938 64454 569174
rect 63834 533494 64454 568938
rect 65563 565724 65629 565725
rect 65563 565660 65564 565724
rect 65628 565660 65629 565724
rect 65563 565659 65629 565660
rect 63834 533258 63866 533494
rect 64102 533258 64186 533494
rect 64422 533258 64454 533494
rect 63834 533174 64454 533258
rect 63834 532938 63866 533174
rect 64102 532938 64186 533174
rect 64422 532938 64454 533174
rect 63834 497494 64454 532938
rect 63834 497258 63866 497494
rect 64102 497258 64186 497494
rect 64422 497258 64454 497494
rect 63834 497174 64454 497258
rect 63834 496938 63866 497174
rect 64102 496938 64186 497174
rect 64422 496938 64454 497174
rect 63834 461494 64454 496938
rect 65566 492693 65626 565659
rect 66115 552668 66181 552669
rect 66115 552604 66116 552668
rect 66180 552604 66181 552668
rect 66115 552603 66181 552604
rect 65931 543964 65997 543965
rect 65931 543900 65932 543964
rect 65996 543900 65997 543964
rect 65931 543899 65997 543900
rect 65747 535260 65813 535261
rect 65747 535196 65748 535260
rect 65812 535196 65813 535260
rect 65747 535195 65813 535196
rect 65563 492692 65629 492693
rect 65563 492628 65564 492692
rect 65628 492628 65629 492692
rect 65563 492627 65629 492628
rect 65563 491740 65629 491741
rect 65563 491676 65564 491740
rect 65628 491676 65629 491740
rect 65563 491675 65629 491676
rect 63834 461258 63866 461494
rect 64102 461258 64186 461494
rect 64422 461258 64454 461494
rect 63834 461174 64454 461258
rect 63834 460938 63866 461174
rect 64102 460938 64186 461174
rect 64422 460938 64454 461174
rect 63834 425494 64454 460938
rect 63834 425258 63866 425494
rect 64102 425258 64186 425494
rect 64422 425258 64454 425494
rect 63834 425174 64454 425258
rect 63834 424938 63866 425174
rect 64102 424938 64186 425174
rect 64422 424938 64454 425174
rect 63834 389494 64454 424938
rect 63834 389258 63866 389494
rect 64102 389258 64186 389494
rect 64422 389258 64454 389494
rect 63834 389174 64454 389258
rect 63834 388938 63866 389174
rect 64102 388938 64186 389174
rect 64422 388938 64454 389174
rect 63834 353494 64454 388938
rect 63834 353258 63866 353494
rect 64102 353258 64186 353494
rect 64422 353258 64454 353494
rect 63834 353174 64454 353258
rect 63834 352938 63866 353174
rect 64102 352938 64186 353174
rect 64422 352938 64454 353174
rect 63355 344044 63421 344045
rect 63355 343980 63356 344044
rect 63420 343980 63421 344044
rect 63355 343979 63421 343980
rect 63834 340449 64454 352938
rect 65566 341053 65626 491675
rect 65750 341597 65810 535195
rect 65747 341596 65813 341597
rect 65747 341532 65748 341596
rect 65812 341532 65813 341596
rect 65747 341531 65813 341532
rect 65934 341461 65994 543899
rect 66118 341869 66178 552603
rect 66854 540973 66914 574363
rect 67403 561372 67469 561373
rect 67403 561308 67404 561372
rect 67468 561308 67469 561372
rect 67403 561307 67469 561308
rect 67219 557020 67285 557021
rect 67219 556956 67220 557020
rect 67284 556956 67285 557020
rect 67219 556955 67285 556956
rect 67035 548316 67101 548317
rect 67035 548252 67036 548316
rect 67100 548252 67101 548316
rect 67035 548251 67101 548252
rect 66851 540972 66917 540973
rect 66851 540908 66852 540972
rect 66916 540908 66917 540972
rect 66851 540907 66917 540908
rect 66851 539612 66917 539613
rect 66851 539548 66852 539612
rect 66916 539548 66917 539612
rect 66851 539547 66917 539548
rect 66115 341868 66181 341869
rect 66115 341804 66116 341868
rect 66180 341804 66181 341868
rect 66115 341803 66181 341804
rect 66854 341733 66914 539547
rect 66851 341732 66917 341733
rect 66851 341668 66852 341732
rect 66916 341668 66917 341732
rect 66851 341667 66917 341668
rect 65931 341460 65997 341461
rect 65931 341396 65932 341460
rect 65996 341396 65997 341460
rect 65931 341395 65997 341396
rect 67038 341325 67098 548251
rect 67035 341324 67101 341325
rect 67035 341260 67036 341324
rect 67100 341260 67101 341324
rect 67035 341259 67101 341260
rect 67222 341189 67282 556955
rect 67406 342141 67466 561307
rect 68142 525877 68202 609179
rect 68323 604892 68389 604893
rect 68323 604828 68324 604892
rect 68388 604828 68389 604892
rect 68323 604827 68389 604828
rect 68139 525876 68205 525877
rect 68139 525812 68140 525876
rect 68204 525812 68205 525876
rect 68139 525811 68205 525812
rect 68326 523021 68386 604827
rect 68510 604485 68570 626587
rect 68691 622300 68757 622301
rect 68691 622236 68692 622300
rect 68756 622236 68757 622300
rect 68691 622235 68757 622236
rect 68507 604484 68573 604485
rect 68507 604420 68508 604484
rect 68572 604420 68573 604484
rect 68507 604419 68573 604420
rect 68694 601085 68754 622235
rect 89568 619174 89888 619206
rect 89568 618938 89610 619174
rect 89846 618938 89888 619174
rect 89568 618854 89888 618938
rect 89568 618618 89610 618854
rect 89846 618618 89888 618854
rect 89568 618586 89888 618618
rect 120288 619174 120608 619206
rect 120288 618938 120330 619174
rect 120566 618938 120608 619174
rect 120288 618854 120608 618938
rect 120288 618618 120330 618854
rect 120566 618618 120608 618854
rect 120288 618586 120608 618618
rect 151008 619174 151328 619206
rect 151008 618938 151050 619174
rect 151286 618938 151328 619174
rect 151008 618854 151328 618938
rect 151008 618618 151050 618854
rect 151286 618618 151328 618854
rect 151008 618586 151328 618618
rect 181728 619174 182048 619206
rect 181728 618938 181770 619174
rect 182006 618938 182048 619174
rect 181728 618854 182048 618938
rect 181728 618618 181770 618854
rect 182006 618618 182048 618854
rect 181728 618586 182048 618618
rect 212448 619174 212768 619206
rect 212448 618938 212490 619174
rect 212726 618938 212768 619174
rect 212448 618854 212768 618938
rect 212448 618618 212490 618854
rect 212726 618618 212768 618854
rect 212448 618586 212768 618618
rect 243168 619174 243488 619206
rect 243168 618938 243210 619174
rect 243446 618938 243488 619174
rect 243168 618854 243488 618938
rect 243168 618618 243210 618854
rect 243446 618618 243488 618854
rect 243168 618586 243488 618618
rect 273888 619174 274208 619206
rect 273888 618938 273930 619174
rect 274166 618938 274208 619174
rect 273888 618854 274208 618938
rect 273888 618618 273930 618854
rect 274166 618618 274208 618854
rect 273888 618586 274208 618618
rect 68875 617948 68941 617949
rect 68875 617884 68876 617948
rect 68940 617884 68941 617948
rect 68875 617883 68941 617884
rect 68691 601084 68757 601085
rect 68691 601020 68692 601084
rect 68756 601020 68757 601084
rect 68691 601019 68757 601020
rect 68507 600540 68573 600541
rect 68507 600476 68508 600540
rect 68572 600476 68573 600540
rect 68507 600475 68573 600476
rect 68323 523020 68389 523021
rect 68323 522956 68324 523020
rect 68388 522956 68389 523020
rect 68323 522955 68389 522956
rect 67955 522204 68021 522205
rect 67955 522140 67956 522204
rect 68020 522140 68021 522204
rect 67955 522139 68021 522140
rect 67958 500853 68018 522139
rect 68139 517852 68205 517853
rect 68139 517788 68140 517852
rect 68204 517788 68205 517852
rect 68139 517787 68205 517788
rect 67955 500852 68021 500853
rect 67955 500788 67956 500852
rect 68020 500788 68021 500852
rect 67955 500787 68021 500788
rect 68142 461549 68202 517787
rect 68510 517581 68570 600475
rect 68878 531317 68938 617883
rect 74208 615454 74528 615486
rect 74208 615218 74250 615454
rect 74486 615218 74528 615454
rect 74208 615134 74528 615218
rect 74208 614898 74250 615134
rect 74486 614898 74528 615134
rect 74208 614866 74528 614898
rect 104928 615454 105248 615486
rect 104928 615218 104970 615454
rect 105206 615218 105248 615454
rect 104928 615134 105248 615218
rect 104928 614898 104970 615134
rect 105206 614898 105248 615134
rect 104928 614866 105248 614898
rect 135648 615454 135968 615486
rect 135648 615218 135690 615454
rect 135926 615218 135968 615454
rect 135648 615134 135968 615218
rect 135648 614898 135690 615134
rect 135926 614898 135968 615134
rect 135648 614866 135968 614898
rect 166368 615454 166688 615486
rect 166368 615218 166410 615454
rect 166646 615218 166688 615454
rect 166368 615134 166688 615218
rect 166368 614898 166410 615134
rect 166646 614898 166688 615134
rect 166368 614866 166688 614898
rect 197088 615454 197408 615486
rect 197088 615218 197130 615454
rect 197366 615218 197408 615454
rect 197088 615134 197408 615218
rect 197088 614898 197130 615134
rect 197366 614898 197408 615134
rect 197088 614866 197408 614898
rect 227808 615454 228128 615486
rect 227808 615218 227850 615454
rect 228086 615218 228128 615454
rect 227808 615134 228128 615218
rect 227808 614898 227850 615134
rect 228086 614898 228128 615134
rect 227808 614866 228128 614898
rect 258528 615454 258848 615486
rect 258528 615218 258570 615454
rect 258806 615218 258848 615454
rect 258528 615134 258848 615218
rect 258528 614898 258570 615134
rect 258806 614898 258848 615134
rect 258528 614866 258848 614898
rect 289794 615454 290414 650898
rect 293514 705798 294134 711590
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 691174 294134 705242
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 291147 626380 291213 626381
rect 291147 626316 291148 626380
rect 291212 626316 291213 626380
rect 291147 626315 291213 626316
rect 290595 622300 290661 622301
rect 290595 622236 290596 622300
rect 290660 622236 290661 622300
rect 290595 622235 290661 622236
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 70163 613596 70229 613597
rect 70163 613532 70164 613596
rect 70228 613532 70229 613596
rect 70163 613531 70229 613532
rect 69611 596188 69677 596189
rect 69611 596124 69612 596188
rect 69676 596124 69677 596188
rect 69611 596123 69677 596124
rect 69427 578780 69493 578781
rect 69427 578716 69428 578780
rect 69492 578716 69493 578780
rect 69427 578715 69493 578716
rect 68875 531316 68941 531317
rect 68875 531252 68876 531316
rect 68940 531252 68941 531316
rect 68875 531251 68941 531252
rect 68691 530908 68757 530909
rect 68691 530844 68692 530908
rect 68756 530844 68757 530908
rect 68691 530843 68757 530844
rect 68507 517580 68573 517581
rect 68507 517516 68508 517580
rect 68572 517516 68573 517580
rect 68507 517515 68573 517516
rect 68694 514045 68754 530843
rect 68875 526556 68941 526557
rect 68875 526492 68876 526556
rect 68940 526492 68941 526556
rect 68875 526491 68941 526492
rect 68691 514044 68757 514045
rect 68691 513980 68692 514044
rect 68756 513980 68757 514044
rect 68691 513979 68757 513980
rect 68691 513500 68757 513501
rect 68691 513436 68692 513500
rect 68756 513436 68757 513500
rect 68691 513435 68757 513436
rect 68507 509148 68573 509149
rect 68507 509084 68508 509148
rect 68572 509084 68573 509148
rect 68507 509083 68573 509084
rect 68323 500444 68389 500445
rect 68323 500380 68324 500444
rect 68388 500380 68389 500444
rect 68323 500379 68389 500380
rect 68326 476917 68386 500379
rect 68323 476916 68389 476917
rect 68323 476852 68324 476916
rect 68388 476852 68389 476916
rect 68323 476851 68389 476852
rect 68510 474197 68570 509083
rect 68507 474196 68573 474197
rect 68507 474132 68508 474196
rect 68572 474132 68573 474196
rect 68507 474131 68573 474132
rect 68694 469845 68754 513435
rect 68878 507925 68938 526491
rect 68875 507924 68941 507925
rect 68875 507860 68876 507924
rect 68940 507860 68941 507924
rect 68875 507859 68941 507860
rect 68691 469844 68757 469845
rect 68691 469780 68692 469844
rect 68756 469780 68757 469844
rect 68691 469779 68757 469780
rect 68139 461548 68205 461549
rect 68139 461484 68140 461548
rect 68204 461484 68205 461548
rect 68139 461483 68205 461484
rect 67403 342140 67469 342141
rect 67403 342076 67404 342140
rect 67468 342076 67469 342140
rect 67403 342075 67469 342076
rect 69430 342005 69490 578715
rect 69614 496365 69674 596123
rect 69979 582588 70045 582589
rect 69979 582524 69980 582588
rect 70044 582524 70045 582588
rect 69979 582523 70045 582524
rect 69795 570076 69861 570077
rect 69795 570012 69796 570076
rect 69860 570012 69861 570076
rect 69795 570011 69861 570012
rect 69611 496364 69677 496365
rect 69611 496300 69612 496364
rect 69676 496300 69677 496364
rect 69611 496299 69677 496300
rect 69611 496092 69677 496093
rect 69611 496028 69612 496092
rect 69676 496028 69677 496092
rect 69611 496027 69677 496028
rect 69614 344997 69674 496027
rect 69611 344996 69677 344997
rect 69611 344932 69612 344996
rect 69676 344932 69677 344996
rect 69611 344931 69677 344932
rect 69798 342141 69858 570011
rect 69982 347173 70042 582523
rect 70166 571301 70226 613531
rect 89568 583174 89888 583206
rect 89568 582938 89610 583174
rect 89846 582938 89888 583174
rect 89568 582854 89888 582938
rect 89568 582618 89610 582854
rect 89846 582618 89888 582854
rect 89568 582586 89888 582618
rect 120288 583174 120608 583206
rect 120288 582938 120330 583174
rect 120566 582938 120608 583174
rect 120288 582854 120608 582938
rect 120288 582618 120330 582854
rect 120566 582618 120608 582854
rect 120288 582586 120608 582618
rect 151008 583174 151328 583206
rect 151008 582938 151050 583174
rect 151286 582938 151328 583174
rect 151008 582854 151328 582938
rect 151008 582618 151050 582854
rect 151286 582618 151328 582854
rect 151008 582586 151328 582618
rect 181728 583174 182048 583206
rect 181728 582938 181770 583174
rect 182006 582938 182048 583174
rect 181728 582854 182048 582938
rect 181728 582618 181770 582854
rect 182006 582618 182048 582854
rect 181728 582586 182048 582618
rect 212448 583174 212768 583206
rect 212448 582938 212490 583174
rect 212726 582938 212768 583174
rect 212448 582854 212768 582938
rect 212448 582618 212490 582854
rect 212726 582618 212768 582854
rect 212448 582586 212768 582618
rect 243168 583174 243488 583206
rect 243168 582938 243210 583174
rect 243446 582938 243488 583174
rect 243168 582854 243488 582938
rect 243168 582618 243210 582854
rect 243446 582618 243488 582854
rect 243168 582586 243488 582618
rect 273888 583174 274208 583206
rect 273888 582938 273930 583174
rect 274166 582938 274208 583174
rect 273888 582854 274208 582938
rect 273888 582618 273930 582854
rect 274166 582618 274208 582854
rect 273888 582586 274208 582618
rect 74208 579454 74528 579486
rect 74208 579218 74250 579454
rect 74486 579218 74528 579454
rect 74208 579134 74528 579218
rect 74208 578898 74250 579134
rect 74486 578898 74528 579134
rect 74208 578866 74528 578898
rect 104928 579454 105248 579486
rect 104928 579218 104970 579454
rect 105206 579218 105248 579454
rect 104928 579134 105248 579218
rect 104928 578898 104970 579134
rect 105206 578898 105248 579134
rect 104928 578866 105248 578898
rect 135648 579454 135968 579486
rect 135648 579218 135690 579454
rect 135926 579218 135968 579454
rect 135648 579134 135968 579218
rect 135648 578898 135690 579134
rect 135926 578898 135968 579134
rect 135648 578866 135968 578898
rect 166368 579454 166688 579486
rect 166368 579218 166410 579454
rect 166646 579218 166688 579454
rect 166368 579134 166688 579218
rect 166368 578898 166410 579134
rect 166646 578898 166688 579134
rect 166368 578866 166688 578898
rect 197088 579454 197408 579486
rect 197088 579218 197130 579454
rect 197366 579218 197408 579454
rect 197088 579134 197408 579218
rect 197088 578898 197130 579134
rect 197366 578898 197408 579134
rect 197088 578866 197408 578898
rect 227808 579454 228128 579486
rect 227808 579218 227850 579454
rect 228086 579218 228128 579454
rect 227808 579134 228128 579218
rect 227808 578898 227850 579134
rect 228086 578898 228128 579134
rect 227808 578866 228128 578898
rect 258528 579454 258848 579486
rect 258528 579218 258570 579454
rect 258806 579218 258848 579454
rect 258528 579134 258848 579218
rect 258528 578898 258570 579134
rect 258806 578898 258848 579134
rect 258528 578866 258848 578898
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 70163 571300 70229 571301
rect 70163 571236 70164 571300
rect 70228 571236 70229 571300
rect 70163 571235 70229 571236
rect 89568 547174 89888 547206
rect 89568 546938 89610 547174
rect 89846 546938 89888 547174
rect 89568 546854 89888 546938
rect 89568 546618 89610 546854
rect 89846 546618 89888 546854
rect 89568 546586 89888 546618
rect 120288 547174 120608 547206
rect 120288 546938 120330 547174
rect 120566 546938 120608 547174
rect 120288 546854 120608 546938
rect 120288 546618 120330 546854
rect 120566 546618 120608 546854
rect 120288 546586 120608 546618
rect 151008 547174 151328 547206
rect 151008 546938 151050 547174
rect 151286 546938 151328 547174
rect 151008 546854 151328 546938
rect 151008 546618 151050 546854
rect 151286 546618 151328 546854
rect 151008 546586 151328 546618
rect 181728 547174 182048 547206
rect 181728 546938 181770 547174
rect 182006 546938 182048 547174
rect 181728 546854 182048 546938
rect 181728 546618 181770 546854
rect 182006 546618 182048 546854
rect 181728 546586 182048 546618
rect 212448 547174 212768 547206
rect 212448 546938 212490 547174
rect 212726 546938 212768 547174
rect 212448 546854 212768 546938
rect 212448 546618 212490 546854
rect 212726 546618 212768 546854
rect 212448 546586 212768 546618
rect 243168 547174 243488 547206
rect 243168 546938 243210 547174
rect 243446 546938 243488 547174
rect 243168 546854 243488 546938
rect 243168 546618 243210 546854
rect 243446 546618 243488 546854
rect 243168 546586 243488 546618
rect 273888 547174 274208 547206
rect 273888 546938 273930 547174
rect 274166 546938 274208 547174
rect 273888 546854 274208 546938
rect 273888 546618 273930 546854
rect 274166 546618 274208 546854
rect 273888 546586 274208 546618
rect 74208 543454 74528 543486
rect 74208 543218 74250 543454
rect 74486 543218 74528 543454
rect 74208 543134 74528 543218
rect 74208 542898 74250 543134
rect 74486 542898 74528 543134
rect 74208 542866 74528 542898
rect 104928 543454 105248 543486
rect 104928 543218 104970 543454
rect 105206 543218 105248 543454
rect 104928 543134 105248 543218
rect 104928 542898 104970 543134
rect 105206 542898 105248 543134
rect 104928 542866 105248 542898
rect 135648 543454 135968 543486
rect 135648 543218 135690 543454
rect 135926 543218 135968 543454
rect 135648 543134 135968 543218
rect 135648 542898 135690 543134
rect 135926 542898 135968 543134
rect 135648 542866 135968 542898
rect 166368 543454 166688 543486
rect 166368 543218 166410 543454
rect 166646 543218 166688 543454
rect 166368 543134 166688 543218
rect 166368 542898 166410 543134
rect 166646 542898 166688 543134
rect 166368 542866 166688 542898
rect 197088 543454 197408 543486
rect 197088 543218 197130 543454
rect 197366 543218 197408 543454
rect 197088 543134 197408 543218
rect 197088 542898 197130 543134
rect 197366 542898 197408 543134
rect 197088 542866 197408 542898
rect 227808 543454 228128 543486
rect 227808 543218 227850 543454
rect 228086 543218 228128 543454
rect 227808 543134 228128 543218
rect 227808 542898 227850 543134
rect 228086 542898 228128 543134
rect 227808 542866 228128 542898
rect 258528 543454 258848 543486
rect 258528 543218 258570 543454
rect 258806 543218 258848 543454
rect 258528 543134 258848 543218
rect 258528 542898 258570 543134
rect 258806 542898 258848 543134
rect 258528 542866 258848 542898
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289307 516220 289373 516221
rect 289307 516156 289308 516220
rect 289372 516156 289373 516220
rect 289307 516155 289373 516156
rect 89568 511174 89888 511206
rect 89568 510938 89610 511174
rect 89846 510938 89888 511174
rect 89568 510854 89888 510938
rect 89568 510618 89610 510854
rect 89846 510618 89888 510854
rect 89568 510586 89888 510618
rect 120288 511174 120608 511206
rect 120288 510938 120330 511174
rect 120566 510938 120608 511174
rect 120288 510854 120608 510938
rect 120288 510618 120330 510854
rect 120566 510618 120608 510854
rect 120288 510586 120608 510618
rect 151008 511174 151328 511206
rect 151008 510938 151050 511174
rect 151286 510938 151328 511174
rect 151008 510854 151328 510938
rect 151008 510618 151050 510854
rect 151286 510618 151328 510854
rect 151008 510586 151328 510618
rect 181728 511174 182048 511206
rect 181728 510938 181770 511174
rect 182006 510938 182048 511174
rect 181728 510854 182048 510938
rect 181728 510618 181770 510854
rect 182006 510618 182048 510854
rect 181728 510586 182048 510618
rect 212448 511174 212768 511206
rect 212448 510938 212490 511174
rect 212726 510938 212768 511174
rect 212448 510854 212768 510938
rect 212448 510618 212490 510854
rect 212726 510618 212768 510854
rect 212448 510586 212768 510618
rect 243168 511174 243488 511206
rect 243168 510938 243210 511174
rect 243446 510938 243488 511174
rect 243168 510854 243488 510938
rect 243168 510618 243210 510854
rect 243446 510618 243488 510854
rect 243168 510586 243488 510618
rect 273888 511174 274208 511206
rect 273888 510938 273930 511174
rect 274166 510938 274208 511174
rect 273888 510854 274208 510938
rect 273888 510618 273930 510854
rect 274166 510618 274208 510854
rect 273888 510586 274208 510618
rect 74208 507454 74528 507486
rect 74208 507218 74250 507454
rect 74486 507218 74528 507454
rect 74208 507134 74528 507218
rect 74208 506898 74250 507134
rect 74486 506898 74528 507134
rect 74208 506866 74528 506898
rect 104928 507454 105248 507486
rect 104928 507218 104970 507454
rect 105206 507218 105248 507454
rect 104928 507134 105248 507218
rect 104928 506898 104970 507134
rect 105206 506898 105248 507134
rect 104928 506866 105248 506898
rect 135648 507454 135968 507486
rect 135648 507218 135690 507454
rect 135926 507218 135968 507454
rect 135648 507134 135968 507218
rect 135648 506898 135690 507134
rect 135926 506898 135968 507134
rect 135648 506866 135968 506898
rect 166368 507454 166688 507486
rect 166368 507218 166410 507454
rect 166646 507218 166688 507454
rect 166368 507134 166688 507218
rect 166368 506898 166410 507134
rect 166646 506898 166688 507134
rect 166368 506866 166688 506898
rect 197088 507454 197408 507486
rect 197088 507218 197130 507454
rect 197366 507218 197408 507454
rect 197088 507134 197408 507218
rect 197088 506898 197130 507134
rect 197366 506898 197408 507134
rect 197088 506866 197408 506898
rect 227808 507454 228128 507486
rect 227808 507218 227850 507454
rect 228086 507218 228128 507454
rect 227808 507134 228128 507218
rect 227808 506898 227850 507134
rect 228086 506898 228128 507134
rect 227808 506866 228128 506898
rect 258528 507454 258848 507486
rect 258528 507218 258570 507454
rect 258806 507218 258848 507454
rect 258528 507134 258848 507218
rect 258528 506898 258570 507134
rect 258806 506898 258848 507134
rect 258528 506866 258848 506898
rect 234475 479500 234541 479501
rect 234475 479436 234476 479500
rect 234540 479436 234541 479500
rect 234475 479435 234541 479436
rect 73794 471454 74414 478303
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 69979 347172 70045 347173
rect 69979 347108 69980 347172
rect 70044 347108 70045 347172
rect 69979 347107 70045 347108
rect 69795 342140 69861 342141
rect 69795 342076 69796 342140
rect 69860 342076 69861 342140
rect 69795 342075 69861 342076
rect 69427 342004 69493 342005
rect 69427 341940 69428 342004
rect 69492 341940 69493 342004
rect 69427 341939 69493 341940
rect 67219 341188 67285 341189
rect 67219 341124 67220 341188
rect 67284 341124 67285 341188
rect 67219 341123 67285 341124
rect 65563 341052 65629 341053
rect 65563 340988 65564 341052
rect 65628 340988 65629 341052
rect 65563 340987 65629 340988
rect 73794 340449 74414 362898
rect 77514 475174 78134 478303
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 340449 78134 366618
rect 81234 442894 81854 478303
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 340449 81854 370338
rect 84954 446614 85574 478303
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 340449 85574 374058
rect 88674 450334 89294 478303
rect 88674 450098 88706 450334
rect 88942 450098 89026 450334
rect 89262 450098 89294 450334
rect 88674 450014 89294 450098
rect 88674 449778 88706 450014
rect 88942 449778 89026 450014
rect 89262 449778 89294 450014
rect 88674 414334 89294 449778
rect 88674 414098 88706 414334
rect 88942 414098 89026 414334
rect 89262 414098 89294 414334
rect 88674 414014 89294 414098
rect 88674 413778 88706 414014
rect 88942 413778 89026 414014
rect 89262 413778 89294 414014
rect 88674 378334 89294 413778
rect 88674 378098 88706 378334
rect 88942 378098 89026 378334
rect 89262 378098 89294 378334
rect 88674 378014 89294 378098
rect 88674 377778 88706 378014
rect 88942 377778 89026 378014
rect 89262 377778 89294 378014
rect 88674 342334 89294 377778
rect 88674 342098 88706 342334
rect 88942 342098 89026 342334
rect 89262 342098 89294 342334
rect 88674 342014 89294 342098
rect 88674 341778 88706 342014
rect 88942 341778 89026 342014
rect 89262 341778 89294 342014
rect 88674 340449 89294 341778
rect 92394 454054 93014 478303
rect 92394 453818 92426 454054
rect 92662 453818 92746 454054
rect 92982 453818 93014 454054
rect 92394 453734 93014 453818
rect 92394 453498 92426 453734
rect 92662 453498 92746 453734
rect 92982 453498 93014 453734
rect 92394 418054 93014 453498
rect 92394 417818 92426 418054
rect 92662 417818 92746 418054
rect 92982 417818 93014 418054
rect 92394 417734 93014 417818
rect 92394 417498 92426 417734
rect 92662 417498 92746 417734
rect 92982 417498 93014 417734
rect 92394 382054 93014 417498
rect 92394 381818 92426 382054
rect 92662 381818 92746 382054
rect 92982 381818 93014 382054
rect 92394 381734 93014 381818
rect 92394 381498 92426 381734
rect 92662 381498 92746 381734
rect 92982 381498 93014 381734
rect 92394 346054 93014 381498
rect 92394 345818 92426 346054
rect 92662 345818 92746 346054
rect 92982 345818 93014 346054
rect 92394 345734 93014 345818
rect 92394 345498 92426 345734
rect 92662 345498 92746 345734
rect 92982 345498 93014 345734
rect 92394 340449 93014 345498
rect 96114 457774 96734 478303
rect 96114 457538 96146 457774
rect 96382 457538 96466 457774
rect 96702 457538 96734 457774
rect 96114 457454 96734 457538
rect 96114 457218 96146 457454
rect 96382 457218 96466 457454
rect 96702 457218 96734 457454
rect 96114 421774 96734 457218
rect 96114 421538 96146 421774
rect 96382 421538 96466 421774
rect 96702 421538 96734 421774
rect 96114 421454 96734 421538
rect 96114 421218 96146 421454
rect 96382 421218 96466 421454
rect 96702 421218 96734 421454
rect 96114 385774 96734 421218
rect 96114 385538 96146 385774
rect 96382 385538 96466 385774
rect 96702 385538 96734 385774
rect 96114 385454 96734 385538
rect 96114 385218 96146 385454
rect 96382 385218 96466 385454
rect 96702 385218 96734 385454
rect 96114 349774 96734 385218
rect 96114 349538 96146 349774
rect 96382 349538 96466 349774
rect 96702 349538 96734 349774
rect 96114 349454 96734 349538
rect 96114 349218 96146 349454
rect 96382 349218 96466 349454
rect 96702 349218 96734 349454
rect 96114 340449 96734 349218
rect 99834 461494 100454 478303
rect 99834 461258 99866 461494
rect 100102 461258 100186 461494
rect 100422 461258 100454 461494
rect 99834 461174 100454 461258
rect 99834 460938 99866 461174
rect 100102 460938 100186 461174
rect 100422 460938 100454 461174
rect 99834 425494 100454 460938
rect 99834 425258 99866 425494
rect 100102 425258 100186 425494
rect 100422 425258 100454 425494
rect 99834 425174 100454 425258
rect 99834 424938 99866 425174
rect 100102 424938 100186 425174
rect 100422 424938 100454 425174
rect 99834 389494 100454 424938
rect 99834 389258 99866 389494
rect 100102 389258 100186 389494
rect 100422 389258 100454 389494
rect 99834 389174 100454 389258
rect 99834 388938 99866 389174
rect 100102 388938 100186 389174
rect 100422 388938 100454 389174
rect 99834 353494 100454 388938
rect 99834 353258 99866 353494
rect 100102 353258 100186 353494
rect 100422 353258 100454 353494
rect 99834 353174 100454 353258
rect 99834 352938 99866 353174
rect 100102 352938 100186 353174
rect 100422 352938 100454 353174
rect 99834 340449 100454 352938
rect 109794 471454 110414 478303
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 113514 475174 114134 478303
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 112483 441284 112549 441285
rect 112483 441220 112484 441284
rect 112548 441220 112549 441284
rect 112483 441219 112549 441220
rect 112299 440604 112365 440605
rect 112299 440540 112300 440604
rect 112364 440540 112365 440604
rect 112299 440539 112365 440540
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 399454 110414 434898
rect 109794 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 110414 399454
rect 109794 399134 110414 399218
rect 109794 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 110414 399134
rect 109794 363454 110414 398898
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 340449 110414 362898
rect 111747 339420 111813 339421
rect 111747 339356 111748 339420
rect 111812 339356 111813 339420
rect 111747 339355 111813 339356
rect 69568 331174 69888 331206
rect 69568 330938 69610 331174
rect 69846 330938 69888 331174
rect 69568 330854 69888 330938
rect 69568 330618 69610 330854
rect 69846 330618 69888 330854
rect 69568 330586 69888 330618
rect 100288 331174 100608 331206
rect 100288 330938 100330 331174
rect 100566 330938 100608 331174
rect 100288 330854 100608 330938
rect 100288 330618 100330 330854
rect 100566 330618 100608 330854
rect 100288 330586 100608 330618
rect 84928 327454 85248 327486
rect 84928 327218 84970 327454
rect 85206 327218 85248 327454
rect 84928 327134 85248 327218
rect 84928 326898 84970 327134
rect 85206 326898 85248 327134
rect 84928 326866 85248 326898
rect 111750 312493 111810 339355
rect 111931 322964 111997 322965
rect 111931 322900 111932 322964
rect 111996 322900 111997 322964
rect 111931 322899 111997 322900
rect 111747 312492 111813 312493
rect 111747 312428 111748 312492
rect 111812 312428 111813 312492
rect 111747 312427 111813 312428
rect 56394 309818 56426 310054
rect 56662 309818 56746 310054
rect 56982 309818 57014 310054
rect 56394 309734 57014 309818
rect 56394 309498 56426 309734
rect 56662 309498 56746 309734
rect 56982 309498 57014 309734
rect 54208 291454 54528 291486
rect 54208 291218 54250 291454
rect 54486 291218 54528 291454
rect 54208 291134 54528 291218
rect 54208 290898 54250 291134
rect 54486 290898 54528 291134
rect 54208 290866 54528 290898
rect 52674 270098 52706 270334
rect 52942 270098 53026 270334
rect 53262 270098 53294 270334
rect 52674 270014 53294 270098
rect 52674 269778 52706 270014
rect 52942 269778 53026 270014
rect 53262 269778 53294 270014
rect 52674 234334 53294 269778
rect 52674 234098 52706 234334
rect 52942 234098 53026 234334
rect 53262 234098 53294 234334
rect 52674 234014 53294 234098
rect 52674 233778 52706 234014
rect 52942 233778 53026 234014
rect 53262 233778 53294 234014
rect 52674 198334 53294 233778
rect 52674 198098 52706 198334
rect 52942 198098 53026 198334
rect 53262 198098 53294 198334
rect 52674 198014 53294 198098
rect 52674 197778 52706 198014
rect 52942 197778 53026 198014
rect 53262 197778 53294 198014
rect 52674 162334 53294 197778
rect 52674 162098 52706 162334
rect 52942 162098 53026 162334
rect 53262 162098 53294 162334
rect 52674 162014 53294 162098
rect 52674 161778 52706 162014
rect 52942 161778 53026 162014
rect 53262 161778 53294 162014
rect 52674 126334 53294 161778
rect 52674 126098 52706 126334
rect 52942 126098 53026 126334
rect 53262 126098 53294 126334
rect 52674 126014 53294 126098
rect 52674 125778 52706 126014
rect 52942 125778 53026 126014
rect 53262 125778 53294 126014
rect 52674 90334 53294 125778
rect 52674 90098 52706 90334
rect 52942 90098 53026 90334
rect 53262 90098 53294 90334
rect 52674 90014 53294 90098
rect 52674 89778 52706 90014
rect 52942 89778 53026 90014
rect 53262 89778 53294 90014
rect 52674 54334 53294 89778
rect 56394 274054 57014 309498
rect 111934 307597 111994 322899
rect 112302 309229 112362 440539
rect 112486 320653 112546 441219
rect 112851 440468 112917 440469
rect 112851 440404 112852 440468
rect 112916 440404 112917 440468
rect 112851 440403 112917 440404
rect 112667 438972 112733 438973
rect 112667 438908 112668 438972
rect 112732 438908 112733 438972
rect 112667 438907 112733 438908
rect 112670 323917 112730 438907
rect 112854 338605 112914 440403
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 112851 338604 112917 338605
rect 112851 338540 112852 338604
rect 112916 338540 112917 338604
rect 112851 338539 112917 338540
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 112667 323916 112733 323917
rect 112667 323852 112668 323916
rect 112732 323852 112733 323916
rect 112667 323851 112733 323852
rect 112483 320652 112549 320653
rect 112483 320588 112484 320652
rect 112548 320588 112549 320652
rect 112483 320587 112549 320588
rect 112299 309228 112365 309229
rect 112299 309164 112300 309228
rect 112364 309164 112365 309228
rect 112299 309163 112365 309164
rect 111931 307596 111997 307597
rect 111931 307532 111932 307596
rect 111996 307532 111997 307596
rect 111931 307531 111997 307532
rect 69568 295174 69888 295206
rect 69568 294938 69610 295174
rect 69846 294938 69888 295174
rect 69568 294854 69888 294938
rect 69568 294618 69610 294854
rect 69846 294618 69888 294854
rect 69568 294586 69888 294618
rect 100288 295174 100608 295206
rect 100288 294938 100330 295174
rect 100566 294938 100608 295174
rect 100288 294854 100608 294938
rect 100288 294618 100330 294854
rect 100566 294618 100608 294854
rect 100288 294586 100608 294618
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 84928 291454 85248 291486
rect 84928 291218 84970 291454
rect 85206 291218 85248 291454
rect 84928 291134 85248 291218
rect 84928 290898 84970 291134
rect 85206 290898 85248 291134
rect 84928 290866 85248 290898
rect 56394 273818 56426 274054
rect 56662 273818 56746 274054
rect 56982 273818 57014 274054
rect 56394 273734 57014 273818
rect 56394 273498 56426 273734
rect 56662 273498 56746 273734
rect 56982 273498 57014 273734
rect 56394 238054 57014 273498
rect 56394 237818 56426 238054
rect 56662 237818 56746 238054
rect 56982 237818 57014 238054
rect 56394 237734 57014 237818
rect 56394 237498 56426 237734
rect 56662 237498 56746 237734
rect 56982 237498 57014 237734
rect 56394 202054 57014 237498
rect 56394 201818 56426 202054
rect 56662 201818 56746 202054
rect 56982 201818 57014 202054
rect 56394 201734 57014 201818
rect 56394 201498 56426 201734
rect 56662 201498 56746 201734
rect 56982 201498 57014 201734
rect 56394 166054 57014 201498
rect 56394 165818 56426 166054
rect 56662 165818 56746 166054
rect 56982 165818 57014 166054
rect 56394 165734 57014 165818
rect 56394 165498 56426 165734
rect 56662 165498 56746 165734
rect 56982 165498 57014 165734
rect 56394 130054 57014 165498
rect 56394 129818 56426 130054
rect 56662 129818 56746 130054
rect 56982 129818 57014 130054
rect 56394 129734 57014 129818
rect 56394 129498 56426 129734
rect 56662 129498 56746 129734
rect 56982 129498 57014 129734
rect 56394 94054 57014 129498
rect 56394 93818 56426 94054
rect 56662 93818 56746 94054
rect 56982 93818 57014 94054
rect 56394 93734 57014 93818
rect 56394 93498 56426 93734
rect 56662 93498 56746 93734
rect 56982 93498 57014 93734
rect 55038 75454 55358 75486
rect 55038 75218 55080 75454
rect 55316 75218 55358 75454
rect 55038 75134 55358 75218
rect 55038 74898 55080 75134
rect 55316 74898 55358 75134
rect 55038 74866 55358 74898
rect 52674 54098 52706 54334
rect 52942 54098 53026 54334
rect 53262 54098 53294 54334
rect 52674 54014 53294 54098
rect 52674 53778 52706 54014
rect 52942 53778 53026 54014
rect 53262 53778 53294 54014
rect 52674 18334 53294 53778
rect 52674 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 53294 18334
rect 52674 18014 53294 18098
rect 52674 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 53294 18014
rect 52674 -4186 53294 17778
rect 52674 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 53294 -4186
rect 52674 -4506 53294 -4422
rect 52674 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 53294 -4506
rect 52674 -7654 53294 -4742
rect 56394 58054 57014 93498
rect 60114 277774 60734 278167
rect 60114 277538 60146 277774
rect 60382 277538 60466 277774
rect 60702 277538 60734 277774
rect 60114 277454 60734 277538
rect 60114 277218 60146 277454
rect 60382 277218 60466 277454
rect 60702 277218 60734 277454
rect 60114 241774 60734 277218
rect 60114 241538 60146 241774
rect 60382 241538 60466 241774
rect 60702 241538 60734 241774
rect 60114 241454 60734 241538
rect 60114 241218 60146 241454
rect 60382 241218 60466 241454
rect 60702 241218 60734 241454
rect 60114 205774 60734 241218
rect 60114 205538 60146 205774
rect 60382 205538 60466 205774
rect 60702 205538 60734 205774
rect 60114 205454 60734 205538
rect 60114 205218 60146 205454
rect 60382 205218 60466 205454
rect 60702 205218 60734 205454
rect 60114 169774 60734 205218
rect 60114 169538 60146 169774
rect 60382 169538 60466 169774
rect 60702 169538 60734 169774
rect 60114 169454 60734 169538
rect 60114 169218 60146 169454
rect 60382 169218 60466 169454
rect 60702 169218 60734 169454
rect 60114 133774 60734 169218
rect 60114 133538 60146 133774
rect 60382 133538 60466 133774
rect 60702 133538 60734 133774
rect 60114 133454 60734 133538
rect 60114 133218 60146 133454
rect 60382 133218 60466 133454
rect 60702 133218 60734 133454
rect 60114 97774 60734 133218
rect 60114 97538 60146 97774
rect 60382 97538 60466 97774
rect 60702 97538 60734 97774
rect 60114 97454 60734 97538
rect 60114 97218 60146 97454
rect 60382 97218 60466 97454
rect 60702 97218 60734 97454
rect 59132 79174 59452 79206
rect 59132 78938 59174 79174
rect 59410 78938 59452 79174
rect 59132 78854 59452 78938
rect 59132 78618 59174 78854
rect 59410 78618 59452 78854
rect 59132 78586 59452 78618
rect 56394 57818 56426 58054
rect 56662 57818 56746 58054
rect 56982 57818 57014 58054
rect 56394 57734 57014 57818
rect 56394 57498 56426 57734
rect 56662 57498 56746 57734
rect 56982 57498 57014 57734
rect 56394 22054 57014 57498
rect 56394 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 57014 22054
rect 56394 21734 57014 21818
rect 56394 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 57014 21734
rect 56394 -5146 57014 21498
rect 56394 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 57014 -5146
rect 56394 -5466 57014 -5382
rect 56394 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 57014 -5466
rect 56394 -7654 57014 -5702
rect 60114 61774 60734 97218
rect 63834 245494 64454 278167
rect 63834 245258 63866 245494
rect 64102 245258 64186 245494
rect 64422 245258 64454 245494
rect 63834 245174 64454 245258
rect 63834 244938 63866 245174
rect 64102 244938 64186 245174
rect 64422 244938 64454 245174
rect 63834 209494 64454 244938
rect 63834 209258 63866 209494
rect 64102 209258 64186 209494
rect 64422 209258 64454 209494
rect 63834 209174 64454 209258
rect 63834 208938 63866 209174
rect 64102 208938 64186 209174
rect 64422 208938 64454 209174
rect 63834 173494 64454 208938
rect 63834 173258 63866 173494
rect 64102 173258 64186 173494
rect 64422 173258 64454 173494
rect 63834 173174 64454 173258
rect 63834 172938 63866 173174
rect 64102 172938 64186 173174
rect 64422 172938 64454 173174
rect 63834 137494 64454 172938
rect 63834 137258 63866 137494
rect 64102 137258 64186 137494
rect 64422 137258 64454 137494
rect 63834 137174 64454 137258
rect 63834 136938 63866 137174
rect 64102 136938 64186 137174
rect 64422 136938 64454 137174
rect 63834 101494 64454 136938
rect 63834 101258 63866 101494
rect 64102 101258 64186 101494
rect 64422 101258 64454 101494
rect 63834 101174 64454 101258
rect 63834 100938 63866 101174
rect 64102 100938 64186 101174
rect 64422 100938 64454 101174
rect 63226 75454 63546 75486
rect 63226 75218 63268 75454
rect 63504 75218 63546 75454
rect 63226 75134 63546 75218
rect 63226 74898 63268 75134
rect 63504 74898 63546 75134
rect 63226 74866 63546 74898
rect 60114 61538 60146 61774
rect 60382 61538 60466 61774
rect 60702 61538 60734 61774
rect 60114 61454 60734 61538
rect 60114 61218 60146 61454
rect 60382 61218 60466 61454
rect 60702 61218 60734 61454
rect 60114 25774 60734 61218
rect 60114 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 60734 25774
rect 60114 25454 60734 25538
rect 60114 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 60734 25454
rect 60114 -6106 60734 25218
rect 60114 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 60734 -6106
rect 60114 -6426 60734 -6342
rect 60114 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 60734 -6426
rect 60114 -7654 60734 -6662
rect 63834 65494 64454 100938
rect 73794 255454 74414 278167
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 67320 79174 67640 79206
rect 67320 78938 67362 79174
rect 67598 78938 67640 79174
rect 67320 78854 67640 78938
rect 67320 78618 67362 78854
rect 67598 78618 67640 78854
rect 67320 78586 67640 78618
rect 71414 75454 71734 75486
rect 71414 75218 71456 75454
rect 71692 75218 71734 75454
rect 71414 75134 71734 75218
rect 71414 74898 71456 75134
rect 71692 74898 71734 75134
rect 71414 74866 71734 74898
rect 73794 75454 74414 110898
rect 77514 259174 78134 278167
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 75508 79174 75828 79206
rect 75508 78938 75550 79174
rect 75786 78938 75828 79174
rect 75508 78854 75828 78938
rect 75508 78618 75550 78854
rect 75786 78618 75828 78854
rect 75508 78586 75828 78618
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 63834 65258 63866 65494
rect 64102 65258 64186 65494
rect 64422 65258 64454 65494
rect 63834 65174 64454 65258
rect 63834 64938 63866 65174
rect 64102 64938 64186 65174
rect 64422 64938 64454 65174
rect 63834 29494 64454 64938
rect 63834 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 64454 29494
rect 63834 29174 64454 29258
rect 63834 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 64454 29174
rect 63834 -7066 64454 28938
rect 63834 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 64454 -7066
rect 63834 -7386 64454 -7302
rect 63834 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 64454 -7386
rect 63834 -7654 64454 -7622
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 77514 43174 78134 78618
rect 81234 262894 81854 278167
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 79602 75454 79922 75486
rect 79602 75218 79644 75454
rect 79880 75218 79922 75454
rect 79602 75134 79922 75218
rect 79602 74898 79644 75134
rect 79880 74898 79922 75134
rect 79602 74866 79922 74898
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -1306 78134 6618
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -7654 78134 -1862
rect 81234 46894 81854 82338
rect 84954 266614 85574 278167
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 83696 79174 84016 79206
rect 83696 78938 83738 79174
rect 83974 78938 84016 79174
rect 83696 78854 84016 78938
rect 83696 78618 83738 78854
rect 83974 78618 84016 78854
rect 83696 78586 84016 78618
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -2266 81854 10338
rect 81234 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 81854 -2266
rect 81234 -2586 81854 -2502
rect 81234 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 81854 -2586
rect 81234 -7654 81854 -2822
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 84954 -3226 85574 14058
rect 84954 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 85574 -3226
rect 84954 -3546 85574 -3462
rect 84954 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 85574 -3546
rect 84954 -7654 85574 -3782
rect 88674 270334 89294 278167
rect 88674 270098 88706 270334
rect 88942 270098 89026 270334
rect 89262 270098 89294 270334
rect 88674 270014 89294 270098
rect 88674 269778 88706 270014
rect 88942 269778 89026 270014
rect 89262 269778 89294 270014
rect 88674 234334 89294 269778
rect 88674 234098 88706 234334
rect 88942 234098 89026 234334
rect 89262 234098 89294 234334
rect 88674 234014 89294 234098
rect 88674 233778 88706 234014
rect 88942 233778 89026 234014
rect 89262 233778 89294 234014
rect 88674 198334 89294 233778
rect 88674 198098 88706 198334
rect 88942 198098 89026 198334
rect 89262 198098 89294 198334
rect 88674 198014 89294 198098
rect 88674 197778 88706 198014
rect 88942 197778 89026 198014
rect 89262 197778 89294 198014
rect 88674 162334 89294 197778
rect 88674 162098 88706 162334
rect 88942 162098 89026 162334
rect 89262 162098 89294 162334
rect 88674 162014 89294 162098
rect 88674 161778 88706 162014
rect 88942 161778 89026 162014
rect 89262 161778 89294 162014
rect 88674 126334 89294 161778
rect 88674 126098 88706 126334
rect 88942 126098 89026 126334
rect 89262 126098 89294 126334
rect 88674 126014 89294 126098
rect 88674 125778 88706 126014
rect 88942 125778 89026 126014
rect 89262 125778 89294 126014
rect 88674 90334 89294 125778
rect 88674 90098 88706 90334
rect 88942 90098 89026 90334
rect 89262 90098 89294 90334
rect 88674 90014 89294 90098
rect 88674 89778 88706 90014
rect 88942 89778 89026 90014
rect 89262 89778 89294 90014
rect 88674 54334 89294 89778
rect 88674 54098 88706 54334
rect 88942 54098 89026 54334
rect 89262 54098 89294 54334
rect 88674 54014 89294 54098
rect 88674 53778 88706 54014
rect 88942 53778 89026 54014
rect 89262 53778 89294 54014
rect 88674 18334 89294 53778
rect 88674 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 89294 18334
rect 88674 18014 89294 18098
rect 88674 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 89294 18014
rect 88674 -4186 89294 17778
rect 88674 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 89294 -4186
rect 88674 -4506 89294 -4422
rect 88674 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 89294 -4506
rect 88674 -7654 89294 -4742
rect 92394 274054 93014 278167
rect 92394 273818 92426 274054
rect 92662 273818 92746 274054
rect 92982 273818 93014 274054
rect 92394 273734 93014 273818
rect 92394 273498 92426 273734
rect 92662 273498 92746 273734
rect 92982 273498 93014 273734
rect 92394 238054 93014 273498
rect 92394 237818 92426 238054
rect 92662 237818 92746 238054
rect 92982 237818 93014 238054
rect 92394 237734 93014 237818
rect 92394 237498 92426 237734
rect 92662 237498 92746 237734
rect 92982 237498 93014 237734
rect 92394 202054 93014 237498
rect 92394 201818 92426 202054
rect 92662 201818 92746 202054
rect 92982 201818 93014 202054
rect 92394 201734 93014 201818
rect 92394 201498 92426 201734
rect 92662 201498 92746 201734
rect 92982 201498 93014 201734
rect 92394 166054 93014 201498
rect 92394 165818 92426 166054
rect 92662 165818 92746 166054
rect 92982 165818 93014 166054
rect 92394 165734 93014 165818
rect 92394 165498 92426 165734
rect 92662 165498 92746 165734
rect 92982 165498 93014 165734
rect 92394 130054 93014 165498
rect 92394 129818 92426 130054
rect 92662 129818 92746 130054
rect 92982 129818 93014 130054
rect 92394 129734 93014 129818
rect 92394 129498 92426 129734
rect 92662 129498 92746 129734
rect 92982 129498 93014 129734
rect 92394 94054 93014 129498
rect 92394 93818 92426 94054
rect 92662 93818 92746 94054
rect 92982 93818 93014 94054
rect 92394 93734 93014 93818
rect 92394 93498 92426 93734
rect 92662 93498 92746 93734
rect 92982 93498 93014 93734
rect 92394 58054 93014 93498
rect 92394 57818 92426 58054
rect 92662 57818 92746 58054
rect 92982 57818 93014 58054
rect 92394 57734 93014 57818
rect 92394 57498 92426 57734
rect 92662 57498 92746 57734
rect 92982 57498 93014 57734
rect 92394 22054 93014 57498
rect 92394 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 93014 22054
rect 92394 21734 93014 21818
rect 92394 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 93014 21734
rect 92394 -5146 93014 21498
rect 92394 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 93014 -5146
rect 92394 -5466 93014 -5382
rect 92394 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 93014 -5466
rect 92394 -7654 93014 -5702
rect 96114 277774 96734 278167
rect 96114 277538 96146 277774
rect 96382 277538 96466 277774
rect 96702 277538 96734 277774
rect 96114 277454 96734 277538
rect 96114 277218 96146 277454
rect 96382 277218 96466 277454
rect 96702 277218 96734 277454
rect 96114 241774 96734 277218
rect 96114 241538 96146 241774
rect 96382 241538 96466 241774
rect 96702 241538 96734 241774
rect 96114 241454 96734 241538
rect 96114 241218 96146 241454
rect 96382 241218 96466 241454
rect 96702 241218 96734 241454
rect 96114 205774 96734 241218
rect 96114 205538 96146 205774
rect 96382 205538 96466 205774
rect 96702 205538 96734 205774
rect 96114 205454 96734 205538
rect 96114 205218 96146 205454
rect 96382 205218 96466 205454
rect 96702 205218 96734 205454
rect 96114 169774 96734 205218
rect 96114 169538 96146 169774
rect 96382 169538 96466 169774
rect 96702 169538 96734 169774
rect 96114 169454 96734 169538
rect 96114 169218 96146 169454
rect 96382 169218 96466 169454
rect 96702 169218 96734 169454
rect 96114 133774 96734 169218
rect 96114 133538 96146 133774
rect 96382 133538 96466 133774
rect 96702 133538 96734 133774
rect 96114 133454 96734 133538
rect 96114 133218 96146 133454
rect 96382 133218 96466 133454
rect 96702 133218 96734 133454
rect 96114 97774 96734 133218
rect 96114 97538 96146 97774
rect 96382 97538 96466 97774
rect 96702 97538 96734 97774
rect 96114 97454 96734 97538
rect 96114 97218 96146 97454
rect 96382 97218 96466 97454
rect 96702 97218 96734 97454
rect 96114 61774 96734 97218
rect 96114 61538 96146 61774
rect 96382 61538 96466 61774
rect 96702 61538 96734 61774
rect 96114 61454 96734 61538
rect 96114 61218 96146 61454
rect 96382 61218 96466 61454
rect 96702 61218 96734 61454
rect 96114 25774 96734 61218
rect 96114 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 96734 25774
rect 96114 25454 96734 25538
rect 96114 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 96734 25454
rect 96114 -6106 96734 25218
rect 96114 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 96734 -6106
rect 96114 -6426 96734 -6342
rect 96114 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 96734 -6426
rect 96114 -7654 96734 -6662
rect 99834 245494 100454 278167
rect 99834 245258 99866 245494
rect 100102 245258 100186 245494
rect 100422 245258 100454 245494
rect 99834 245174 100454 245258
rect 99834 244938 99866 245174
rect 100102 244938 100186 245174
rect 100422 244938 100454 245174
rect 99834 209494 100454 244938
rect 99834 209258 99866 209494
rect 100102 209258 100186 209494
rect 100422 209258 100454 209494
rect 99834 209174 100454 209258
rect 99834 208938 99866 209174
rect 100102 208938 100186 209174
rect 100422 208938 100454 209174
rect 99834 173494 100454 208938
rect 99834 173258 99866 173494
rect 100102 173258 100186 173494
rect 100422 173258 100454 173494
rect 99834 173174 100454 173258
rect 99834 172938 99866 173174
rect 100102 172938 100186 173174
rect 100422 172938 100454 173174
rect 99834 137494 100454 172938
rect 99834 137258 99866 137494
rect 100102 137258 100186 137494
rect 100422 137258 100454 137494
rect 99834 137174 100454 137258
rect 99834 136938 99866 137174
rect 100102 136938 100186 137174
rect 100422 136938 100454 137174
rect 99834 101494 100454 136938
rect 99834 101258 99866 101494
rect 100102 101258 100186 101494
rect 100422 101258 100454 101494
rect 99834 101174 100454 101258
rect 99834 100938 99866 101174
rect 100102 100938 100186 101174
rect 100422 100938 100454 101174
rect 99834 65494 100454 100938
rect 99834 65258 99866 65494
rect 100102 65258 100186 65494
rect 100422 65258 100454 65494
rect 99834 65174 100454 65258
rect 99834 64938 99866 65174
rect 100102 64938 100186 65174
rect 100422 64938 100454 65174
rect 99834 29494 100454 64938
rect 99834 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 100454 29494
rect 99834 29174 100454 29258
rect 99834 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 100454 29174
rect 99834 -7066 100454 28938
rect 99834 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 100454 -7066
rect 99834 -7386 100454 -7302
rect 99834 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 100454 -7386
rect 99834 -7654 100454 -7622
rect 109794 255454 110414 278167
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -1306 114134 6618
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -7654 114134 -1862
rect 117234 442894 117854 478303
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -2266 117854 10338
rect 117234 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 117854 -2266
rect 117234 -2586 117854 -2502
rect 117234 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 117854 -2586
rect 117234 -7654 117854 -2822
rect 120954 446614 121574 478303
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 124674 450334 125294 478303
rect 124674 450098 124706 450334
rect 124942 450098 125026 450334
rect 125262 450098 125294 450334
rect 124674 450014 125294 450098
rect 124674 449778 124706 450014
rect 124942 449778 125026 450014
rect 125262 449778 125294 450014
rect 124674 414334 125294 449778
rect 124674 414098 124706 414334
rect 124942 414098 125026 414334
rect 125262 414098 125294 414334
rect 124674 414014 125294 414098
rect 124674 413778 124706 414014
rect 124942 413778 125026 414014
rect 125262 413778 125294 414014
rect 124674 378334 125294 413778
rect 124674 378098 124706 378334
rect 124942 378098 125026 378334
rect 125262 378098 125294 378334
rect 124674 378014 125294 378098
rect 124674 377778 124706 378014
rect 124942 377778 125026 378014
rect 125262 377778 125294 378014
rect 124674 342334 125294 377778
rect 124674 342098 124706 342334
rect 124942 342098 125026 342334
rect 125262 342098 125294 342334
rect 124674 342014 125294 342098
rect 124674 341778 124706 342014
rect 124942 341778 125026 342014
rect 125262 341778 125294 342014
rect 124674 306334 125294 341778
rect 124674 306098 124706 306334
rect 124942 306098 125026 306334
rect 125262 306098 125294 306334
rect 124674 306014 125294 306098
rect 124674 305778 124706 306014
rect 124942 305778 125026 306014
rect 125262 305778 125294 306014
rect 122051 305692 122117 305693
rect 122051 305628 122052 305692
rect 122116 305628 122117 305692
rect 122051 305627 122117 305628
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 122054 279445 122114 305627
rect 122051 279444 122117 279445
rect 122051 279380 122052 279444
rect 122116 279380 122117 279444
rect 122051 279379 122117 279380
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 120954 -3226 121574 14058
rect 120954 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 121574 -3226
rect 120954 -3546 121574 -3462
rect 120954 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 121574 -3546
rect 120954 -7654 121574 -3782
rect 124674 270334 125294 305778
rect 124674 270098 124706 270334
rect 124942 270098 125026 270334
rect 125262 270098 125294 270334
rect 124674 270014 125294 270098
rect 124674 269778 124706 270014
rect 124942 269778 125026 270014
rect 125262 269778 125294 270014
rect 124674 234334 125294 269778
rect 124674 234098 124706 234334
rect 124942 234098 125026 234334
rect 125262 234098 125294 234334
rect 124674 234014 125294 234098
rect 124674 233778 124706 234014
rect 124942 233778 125026 234014
rect 125262 233778 125294 234014
rect 124674 198334 125294 233778
rect 124674 198098 124706 198334
rect 124942 198098 125026 198334
rect 125262 198098 125294 198334
rect 124674 198014 125294 198098
rect 124674 197778 124706 198014
rect 124942 197778 125026 198014
rect 125262 197778 125294 198014
rect 124674 162334 125294 197778
rect 124674 162098 124706 162334
rect 124942 162098 125026 162334
rect 125262 162098 125294 162334
rect 124674 162014 125294 162098
rect 124674 161778 124706 162014
rect 124942 161778 125026 162014
rect 125262 161778 125294 162014
rect 124674 126334 125294 161778
rect 124674 126098 124706 126334
rect 124942 126098 125026 126334
rect 125262 126098 125294 126334
rect 124674 126014 125294 126098
rect 124674 125778 124706 126014
rect 124942 125778 125026 126014
rect 125262 125778 125294 126014
rect 124674 90334 125294 125778
rect 124674 90098 124706 90334
rect 124942 90098 125026 90334
rect 125262 90098 125294 90334
rect 124674 90014 125294 90098
rect 124674 89778 124706 90014
rect 124942 89778 125026 90014
rect 125262 89778 125294 90014
rect 124674 54334 125294 89778
rect 124674 54098 124706 54334
rect 124942 54098 125026 54334
rect 125262 54098 125294 54334
rect 124674 54014 125294 54098
rect 124674 53778 124706 54014
rect 124942 53778 125026 54014
rect 125262 53778 125294 54014
rect 124674 18334 125294 53778
rect 124674 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 125294 18334
rect 124674 18014 125294 18098
rect 124674 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 125294 18014
rect 124674 -4186 125294 17778
rect 124674 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 125294 -4186
rect 124674 -4506 125294 -4422
rect 124674 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 125294 -4506
rect 124674 -7654 125294 -4742
rect 128394 454054 129014 478303
rect 130331 471204 130397 471205
rect 130331 471140 130332 471204
rect 130396 471140 130397 471204
rect 130331 471139 130397 471140
rect 128394 453818 128426 454054
rect 128662 453818 128746 454054
rect 128982 453818 129014 454054
rect 128394 453734 129014 453818
rect 128394 453498 128426 453734
rect 128662 453498 128746 453734
rect 128982 453498 129014 453734
rect 128394 418054 129014 453498
rect 128394 417818 128426 418054
rect 128662 417818 128746 418054
rect 128982 417818 129014 418054
rect 128394 417734 129014 417818
rect 128394 417498 128426 417734
rect 128662 417498 128746 417734
rect 128982 417498 129014 417734
rect 128394 382054 129014 417498
rect 128394 381818 128426 382054
rect 128662 381818 128746 382054
rect 128982 381818 129014 382054
rect 128394 381734 129014 381818
rect 128394 381498 128426 381734
rect 128662 381498 128746 381734
rect 128982 381498 129014 381734
rect 128394 346054 129014 381498
rect 128394 345818 128426 346054
rect 128662 345818 128746 346054
rect 128982 345818 129014 346054
rect 128394 345734 129014 345818
rect 128394 345498 128426 345734
rect 128662 345498 128746 345734
rect 128982 345498 129014 345734
rect 128394 310054 129014 345498
rect 128394 309818 128426 310054
rect 128662 309818 128746 310054
rect 128982 309818 129014 310054
rect 128394 309734 129014 309818
rect 128394 309498 128426 309734
rect 128662 309498 128746 309734
rect 128982 309498 129014 309734
rect 128394 274054 129014 309498
rect 130334 303517 130394 471139
rect 132114 457774 132734 478303
rect 132114 457538 132146 457774
rect 132382 457538 132466 457774
rect 132702 457538 132734 457774
rect 132114 457454 132734 457538
rect 132114 457218 132146 457454
rect 132382 457218 132466 457454
rect 132702 457218 132734 457454
rect 132114 421774 132734 457218
rect 132114 421538 132146 421774
rect 132382 421538 132466 421774
rect 132702 421538 132734 421774
rect 132114 421454 132734 421538
rect 132114 421218 132146 421454
rect 132382 421218 132466 421454
rect 132702 421218 132734 421454
rect 132114 385774 132734 421218
rect 132114 385538 132146 385774
rect 132382 385538 132466 385774
rect 132702 385538 132734 385774
rect 132114 385454 132734 385538
rect 132114 385218 132146 385454
rect 132382 385218 132466 385454
rect 132702 385218 132734 385454
rect 132114 349774 132734 385218
rect 132114 349538 132146 349774
rect 132382 349538 132466 349774
rect 132702 349538 132734 349774
rect 132114 349454 132734 349538
rect 132114 349218 132146 349454
rect 132382 349218 132466 349454
rect 132702 349218 132734 349454
rect 132114 313774 132734 349218
rect 132114 313538 132146 313774
rect 132382 313538 132466 313774
rect 132702 313538 132734 313774
rect 132114 313454 132734 313538
rect 132114 313218 132146 313454
rect 132382 313218 132466 313454
rect 132702 313218 132734 313454
rect 130331 303516 130397 303517
rect 130331 303452 130332 303516
rect 130396 303452 130397 303516
rect 130331 303451 130397 303452
rect 128394 273818 128426 274054
rect 128662 273818 128746 274054
rect 128982 273818 129014 274054
rect 128394 273734 129014 273818
rect 128394 273498 128426 273734
rect 128662 273498 128746 273734
rect 128982 273498 129014 273734
rect 128394 238054 129014 273498
rect 128394 237818 128426 238054
rect 128662 237818 128746 238054
rect 128982 237818 129014 238054
rect 128394 237734 129014 237818
rect 128394 237498 128426 237734
rect 128662 237498 128746 237734
rect 128982 237498 129014 237734
rect 128394 202054 129014 237498
rect 128394 201818 128426 202054
rect 128662 201818 128746 202054
rect 128982 201818 129014 202054
rect 128394 201734 129014 201818
rect 128394 201498 128426 201734
rect 128662 201498 128746 201734
rect 128982 201498 129014 201734
rect 128394 166054 129014 201498
rect 128394 165818 128426 166054
rect 128662 165818 128746 166054
rect 128982 165818 129014 166054
rect 128394 165734 129014 165818
rect 128394 165498 128426 165734
rect 128662 165498 128746 165734
rect 128982 165498 129014 165734
rect 128394 130054 129014 165498
rect 128394 129818 128426 130054
rect 128662 129818 128746 130054
rect 128982 129818 129014 130054
rect 128394 129734 129014 129818
rect 128394 129498 128426 129734
rect 128662 129498 128746 129734
rect 128982 129498 129014 129734
rect 128394 94054 129014 129498
rect 128394 93818 128426 94054
rect 128662 93818 128746 94054
rect 128982 93818 129014 94054
rect 128394 93734 129014 93818
rect 128394 93498 128426 93734
rect 128662 93498 128746 93734
rect 128982 93498 129014 93734
rect 128394 58054 129014 93498
rect 128394 57818 128426 58054
rect 128662 57818 128746 58054
rect 128982 57818 129014 58054
rect 128394 57734 129014 57818
rect 128394 57498 128426 57734
rect 128662 57498 128746 57734
rect 128982 57498 129014 57734
rect 128394 22054 129014 57498
rect 128394 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 129014 22054
rect 128394 21734 129014 21818
rect 128394 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 129014 21734
rect 128394 -5146 129014 21498
rect 128394 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 129014 -5146
rect 128394 -5466 129014 -5382
rect 128394 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 129014 -5466
rect 128394 -7654 129014 -5702
rect 132114 277774 132734 313218
rect 132114 277538 132146 277774
rect 132382 277538 132466 277774
rect 132702 277538 132734 277774
rect 132114 277454 132734 277538
rect 132114 277218 132146 277454
rect 132382 277218 132466 277454
rect 132702 277218 132734 277454
rect 132114 241774 132734 277218
rect 132114 241538 132146 241774
rect 132382 241538 132466 241774
rect 132702 241538 132734 241774
rect 132114 241454 132734 241538
rect 132114 241218 132146 241454
rect 132382 241218 132466 241454
rect 132702 241218 132734 241454
rect 132114 205774 132734 241218
rect 132114 205538 132146 205774
rect 132382 205538 132466 205774
rect 132702 205538 132734 205774
rect 132114 205454 132734 205538
rect 132114 205218 132146 205454
rect 132382 205218 132466 205454
rect 132702 205218 132734 205454
rect 132114 169774 132734 205218
rect 132114 169538 132146 169774
rect 132382 169538 132466 169774
rect 132702 169538 132734 169774
rect 132114 169454 132734 169538
rect 132114 169218 132146 169454
rect 132382 169218 132466 169454
rect 132702 169218 132734 169454
rect 132114 133774 132734 169218
rect 132114 133538 132146 133774
rect 132382 133538 132466 133774
rect 132702 133538 132734 133774
rect 132114 133454 132734 133538
rect 132114 133218 132146 133454
rect 132382 133218 132466 133454
rect 132702 133218 132734 133454
rect 132114 97774 132734 133218
rect 132114 97538 132146 97774
rect 132382 97538 132466 97774
rect 132702 97538 132734 97774
rect 132114 97454 132734 97538
rect 132114 97218 132146 97454
rect 132382 97218 132466 97454
rect 132702 97218 132734 97454
rect 132114 61774 132734 97218
rect 132114 61538 132146 61774
rect 132382 61538 132466 61774
rect 132702 61538 132734 61774
rect 132114 61454 132734 61538
rect 132114 61218 132146 61454
rect 132382 61218 132466 61454
rect 132702 61218 132734 61454
rect 132114 25774 132734 61218
rect 132114 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 132734 25774
rect 132114 25454 132734 25538
rect 132114 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 132734 25454
rect 132114 -6106 132734 25218
rect 132114 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 132734 -6106
rect 132114 -6426 132734 -6342
rect 132114 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 132734 -6426
rect 132114 -7654 132734 -6662
rect 135834 461494 136454 478303
rect 135834 461258 135866 461494
rect 136102 461258 136186 461494
rect 136422 461258 136454 461494
rect 135834 461174 136454 461258
rect 135834 460938 135866 461174
rect 136102 460938 136186 461174
rect 136422 460938 136454 461174
rect 135834 425494 136454 460938
rect 135834 425258 135866 425494
rect 136102 425258 136186 425494
rect 136422 425258 136454 425494
rect 135834 425174 136454 425258
rect 135834 424938 135866 425174
rect 136102 424938 136186 425174
rect 136422 424938 136454 425174
rect 135834 389494 136454 424938
rect 135834 389258 135866 389494
rect 136102 389258 136186 389494
rect 136422 389258 136454 389494
rect 135834 389174 136454 389258
rect 135834 388938 135866 389174
rect 136102 388938 136186 389174
rect 136422 388938 136454 389174
rect 135834 353494 136454 388938
rect 135834 353258 135866 353494
rect 136102 353258 136186 353494
rect 136422 353258 136454 353494
rect 135834 353174 136454 353258
rect 135834 352938 135866 353174
rect 136102 352938 136186 353174
rect 136422 352938 136454 353174
rect 135834 317494 136454 352938
rect 135834 317258 135866 317494
rect 136102 317258 136186 317494
rect 136422 317258 136454 317494
rect 135834 317174 136454 317258
rect 135834 316938 135866 317174
rect 136102 316938 136186 317174
rect 136422 316938 136454 317174
rect 135834 281494 136454 316938
rect 135834 281258 135866 281494
rect 136102 281258 136186 281494
rect 136422 281258 136454 281494
rect 135834 281174 136454 281258
rect 135834 280938 135866 281174
rect 136102 280938 136186 281174
rect 136422 280938 136454 281174
rect 135834 245494 136454 280938
rect 135834 245258 135866 245494
rect 136102 245258 136186 245494
rect 136422 245258 136454 245494
rect 135834 245174 136454 245258
rect 135834 244938 135866 245174
rect 136102 244938 136186 245174
rect 136422 244938 136454 245174
rect 135834 209494 136454 244938
rect 135834 209258 135866 209494
rect 136102 209258 136186 209494
rect 136422 209258 136454 209494
rect 135834 209174 136454 209258
rect 135834 208938 135866 209174
rect 136102 208938 136186 209174
rect 136422 208938 136454 209174
rect 135834 173494 136454 208938
rect 135834 173258 135866 173494
rect 136102 173258 136186 173494
rect 136422 173258 136454 173494
rect 135834 173174 136454 173258
rect 135834 172938 135866 173174
rect 136102 172938 136186 173174
rect 136422 172938 136454 173174
rect 135834 137494 136454 172938
rect 135834 137258 135866 137494
rect 136102 137258 136186 137494
rect 136422 137258 136454 137494
rect 135834 137174 136454 137258
rect 135834 136938 135866 137174
rect 136102 136938 136186 137174
rect 136422 136938 136454 137174
rect 135834 101494 136454 136938
rect 135834 101258 135866 101494
rect 136102 101258 136186 101494
rect 136422 101258 136454 101494
rect 135834 101174 136454 101258
rect 135834 100938 135866 101174
rect 136102 100938 136186 101174
rect 136422 100938 136454 101174
rect 135834 65494 136454 100938
rect 135834 65258 135866 65494
rect 136102 65258 136186 65494
rect 136422 65258 136454 65494
rect 135834 65174 136454 65258
rect 135834 64938 135866 65174
rect 136102 64938 136186 65174
rect 136422 64938 136454 65174
rect 135834 29494 136454 64938
rect 135834 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 136454 29494
rect 135834 29174 136454 29258
rect 135834 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 136454 29174
rect 135834 -7066 136454 28938
rect 135834 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 136454 -7066
rect 135834 -7386 136454 -7302
rect 135834 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 136454 -7386
rect 135834 -7654 136454 -7622
rect 145794 471454 146414 478303
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 149514 475174 150134 478303
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 147075 345268 147141 345269
rect 147075 345204 147076 345268
rect 147140 345204 147141 345268
rect 147075 345203 147141 345204
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 147078 305149 147138 345203
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 147075 305148 147141 305149
rect 147075 305084 147076 305148
rect 147140 305084 147141 305148
rect 147075 305083 147141 305084
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -1306 150134 6618
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -7654 150134 -1862
rect 153234 442894 153854 478303
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -2266 153854 10338
rect 153234 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 153854 -2266
rect 153234 -2586 153854 -2502
rect 153234 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 153854 -2586
rect 153234 -7654 153854 -2822
rect 156954 446614 157574 478303
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 156954 -3226 157574 14058
rect 156954 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 157574 -3226
rect 156954 -3546 157574 -3462
rect 156954 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 157574 -3546
rect 156954 -7654 157574 -3782
rect 160674 450334 161294 478303
rect 161979 472564 162045 472565
rect 161979 472500 161980 472564
rect 162044 472500 162045 472564
rect 161979 472499 162045 472500
rect 160674 450098 160706 450334
rect 160942 450098 161026 450334
rect 161262 450098 161294 450334
rect 160674 450014 161294 450098
rect 160674 449778 160706 450014
rect 160942 449778 161026 450014
rect 161262 449778 161294 450014
rect 160674 414334 161294 449778
rect 160674 414098 160706 414334
rect 160942 414098 161026 414334
rect 161262 414098 161294 414334
rect 160674 414014 161294 414098
rect 160674 413778 160706 414014
rect 160942 413778 161026 414014
rect 161262 413778 161294 414014
rect 160674 378334 161294 413778
rect 160674 378098 160706 378334
rect 160942 378098 161026 378334
rect 161262 378098 161294 378334
rect 160674 378014 161294 378098
rect 160674 377778 160706 378014
rect 160942 377778 161026 378014
rect 161262 377778 161294 378014
rect 160674 342334 161294 377778
rect 160674 342098 160706 342334
rect 160942 342098 161026 342334
rect 161262 342098 161294 342334
rect 160674 342014 161294 342098
rect 160674 341778 160706 342014
rect 160942 341778 161026 342014
rect 161262 341778 161294 342014
rect 160674 306334 161294 341778
rect 160674 306098 160706 306334
rect 160942 306098 161026 306334
rect 161262 306098 161294 306334
rect 160674 306014 161294 306098
rect 160674 305778 160706 306014
rect 160942 305778 161026 306014
rect 161262 305778 161294 306014
rect 160674 270334 161294 305778
rect 161982 302973 162042 472499
rect 164394 454054 165014 478303
rect 166211 474196 166277 474197
rect 166211 474132 166212 474196
rect 166276 474132 166277 474196
rect 166211 474131 166277 474132
rect 164394 453818 164426 454054
rect 164662 453818 164746 454054
rect 164982 453818 165014 454054
rect 164394 453734 165014 453818
rect 164394 453498 164426 453734
rect 164662 453498 164746 453734
rect 164982 453498 165014 453734
rect 164394 418054 165014 453498
rect 164394 417818 164426 418054
rect 164662 417818 164746 418054
rect 164982 417818 165014 418054
rect 164394 417734 165014 417818
rect 164394 417498 164426 417734
rect 164662 417498 164746 417734
rect 164982 417498 165014 417734
rect 164394 382054 165014 417498
rect 164394 381818 164426 382054
rect 164662 381818 164746 382054
rect 164982 381818 165014 382054
rect 164394 381734 165014 381818
rect 164394 381498 164426 381734
rect 164662 381498 164746 381734
rect 164982 381498 165014 381734
rect 164394 346054 165014 381498
rect 164394 345818 164426 346054
rect 164662 345818 164746 346054
rect 164982 345818 165014 346054
rect 164394 345734 165014 345818
rect 164394 345498 164426 345734
rect 164662 345498 164746 345734
rect 164982 345498 165014 345734
rect 164394 310054 165014 345498
rect 164394 309818 164426 310054
rect 164662 309818 164746 310054
rect 164982 309818 165014 310054
rect 164394 309734 165014 309818
rect 164394 309498 164426 309734
rect 164662 309498 164746 309734
rect 164982 309498 165014 309734
rect 161979 302972 162045 302973
rect 161979 302908 161980 302972
rect 162044 302908 162045 302972
rect 161979 302907 162045 302908
rect 160674 270098 160706 270334
rect 160942 270098 161026 270334
rect 161262 270098 161294 270334
rect 160674 270014 161294 270098
rect 160674 269778 160706 270014
rect 160942 269778 161026 270014
rect 161262 269778 161294 270014
rect 160674 234334 161294 269778
rect 160674 234098 160706 234334
rect 160942 234098 161026 234334
rect 161262 234098 161294 234334
rect 160674 234014 161294 234098
rect 160674 233778 160706 234014
rect 160942 233778 161026 234014
rect 161262 233778 161294 234014
rect 160674 198334 161294 233778
rect 160674 198098 160706 198334
rect 160942 198098 161026 198334
rect 161262 198098 161294 198334
rect 160674 198014 161294 198098
rect 160674 197778 160706 198014
rect 160942 197778 161026 198014
rect 161262 197778 161294 198014
rect 160674 162334 161294 197778
rect 160674 162098 160706 162334
rect 160942 162098 161026 162334
rect 161262 162098 161294 162334
rect 160674 162014 161294 162098
rect 160674 161778 160706 162014
rect 160942 161778 161026 162014
rect 161262 161778 161294 162014
rect 160674 126334 161294 161778
rect 160674 126098 160706 126334
rect 160942 126098 161026 126334
rect 161262 126098 161294 126334
rect 160674 126014 161294 126098
rect 160674 125778 160706 126014
rect 160942 125778 161026 126014
rect 161262 125778 161294 126014
rect 160674 90334 161294 125778
rect 160674 90098 160706 90334
rect 160942 90098 161026 90334
rect 161262 90098 161294 90334
rect 160674 90014 161294 90098
rect 160674 89778 160706 90014
rect 160942 89778 161026 90014
rect 161262 89778 161294 90014
rect 160674 54334 161294 89778
rect 160674 54098 160706 54334
rect 160942 54098 161026 54334
rect 161262 54098 161294 54334
rect 160674 54014 161294 54098
rect 160674 53778 160706 54014
rect 160942 53778 161026 54014
rect 161262 53778 161294 54014
rect 160674 18334 161294 53778
rect 160674 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 161294 18334
rect 160674 18014 161294 18098
rect 160674 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 161294 18014
rect 160674 -4186 161294 17778
rect 160674 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 161294 -4186
rect 160674 -4506 161294 -4422
rect 160674 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 161294 -4506
rect 160674 -7654 161294 -4742
rect 164394 274054 165014 309498
rect 164394 273818 164426 274054
rect 164662 273818 164746 274054
rect 164982 273818 165014 274054
rect 164394 273734 165014 273818
rect 164394 273498 164426 273734
rect 164662 273498 164746 273734
rect 164982 273498 165014 273734
rect 166214 273597 166274 474131
rect 168114 457774 168734 478303
rect 168114 457538 168146 457774
rect 168382 457538 168466 457774
rect 168702 457538 168734 457774
rect 168114 457454 168734 457538
rect 168114 457218 168146 457454
rect 168382 457218 168466 457454
rect 168702 457218 168734 457454
rect 168114 421774 168734 457218
rect 168114 421538 168146 421774
rect 168382 421538 168466 421774
rect 168702 421538 168734 421774
rect 168114 421454 168734 421538
rect 168114 421218 168146 421454
rect 168382 421218 168466 421454
rect 168702 421218 168734 421454
rect 168114 385774 168734 421218
rect 168114 385538 168146 385774
rect 168382 385538 168466 385774
rect 168702 385538 168734 385774
rect 168114 385454 168734 385538
rect 168114 385218 168146 385454
rect 168382 385218 168466 385454
rect 168702 385218 168734 385454
rect 168114 349774 168734 385218
rect 168114 349538 168146 349774
rect 168382 349538 168466 349774
rect 168702 349538 168734 349774
rect 168114 349454 168734 349538
rect 168114 349218 168146 349454
rect 168382 349218 168466 349454
rect 168702 349218 168734 349454
rect 168114 313774 168734 349218
rect 168114 313538 168146 313774
rect 168382 313538 168466 313774
rect 168702 313538 168734 313774
rect 168114 313454 168734 313538
rect 168114 313218 168146 313454
rect 168382 313218 168466 313454
rect 168702 313218 168734 313454
rect 168114 277774 168734 313218
rect 168114 277538 168146 277774
rect 168382 277538 168466 277774
rect 168702 277538 168734 277774
rect 168114 277454 168734 277538
rect 168114 277218 168146 277454
rect 168382 277218 168466 277454
rect 168702 277218 168734 277454
rect 166211 273596 166277 273597
rect 166211 273532 166212 273596
rect 166276 273532 166277 273596
rect 166211 273531 166277 273532
rect 164394 238054 165014 273498
rect 164394 237818 164426 238054
rect 164662 237818 164746 238054
rect 164982 237818 165014 238054
rect 164394 237734 165014 237818
rect 164394 237498 164426 237734
rect 164662 237498 164746 237734
rect 164982 237498 165014 237734
rect 164394 202054 165014 237498
rect 164394 201818 164426 202054
rect 164662 201818 164746 202054
rect 164982 201818 165014 202054
rect 164394 201734 165014 201818
rect 164394 201498 164426 201734
rect 164662 201498 164746 201734
rect 164982 201498 165014 201734
rect 164394 166054 165014 201498
rect 164394 165818 164426 166054
rect 164662 165818 164746 166054
rect 164982 165818 165014 166054
rect 164394 165734 165014 165818
rect 164394 165498 164426 165734
rect 164662 165498 164746 165734
rect 164982 165498 165014 165734
rect 164394 130054 165014 165498
rect 164394 129818 164426 130054
rect 164662 129818 164746 130054
rect 164982 129818 165014 130054
rect 164394 129734 165014 129818
rect 164394 129498 164426 129734
rect 164662 129498 164746 129734
rect 164982 129498 165014 129734
rect 164394 94054 165014 129498
rect 164394 93818 164426 94054
rect 164662 93818 164746 94054
rect 164982 93818 165014 94054
rect 164394 93734 165014 93818
rect 164394 93498 164426 93734
rect 164662 93498 164746 93734
rect 164982 93498 165014 93734
rect 164394 58054 165014 93498
rect 164394 57818 164426 58054
rect 164662 57818 164746 58054
rect 164982 57818 165014 58054
rect 164394 57734 165014 57818
rect 164394 57498 164426 57734
rect 164662 57498 164746 57734
rect 164982 57498 165014 57734
rect 164394 22054 165014 57498
rect 164394 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 165014 22054
rect 164394 21734 165014 21818
rect 164394 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 165014 21734
rect 164394 -5146 165014 21498
rect 164394 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 165014 -5146
rect 164394 -5466 165014 -5382
rect 164394 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 165014 -5466
rect 164394 -7654 165014 -5702
rect 168114 241774 168734 277218
rect 168114 241538 168146 241774
rect 168382 241538 168466 241774
rect 168702 241538 168734 241774
rect 168114 241454 168734 241538
rect 168114 241218 168146 241454
rect 168382 241218 168466 241454
rect 168702 241218 168734 241454
rect 168114 205774 168734 241218
rect 168114 205538 168146 205774
rect 168382 205538 168466 205774
rect 168702 205538 168734 205774
rect 168114 205454 168734 205538
rect 168114 205218 168146 205454
rect 168382 205218 168466 205454
rect 168702 205218 168734 205454
rect 168114 169774 168734 205218
rect 168114 169538 168146 169774
rect 168382 169538 168466 169774
rect 168702 169538 168734 169774
rect 168114 169454 168734 169538
rect 168114 169218 168146 169454
rect 168382 169218 168466 169454
rect 168702 169218 168734 169454
rect 168114 133774 168734 169218
rect 168114 133538 168146 133774
rect 168382 133538 168466 133774
rect 168702 133538 168734 133774
rect 168114 133454 168734 133538
rect 168114 133218 168146 133454
rect 168382 133218 168466 133454
rect 168702 133218 168734 133454
rect 168114 97774 168734 133218
rect 168114 97538 168146 97774
rect 168382 97538 168466 97774
rect 168702 97538 168734 97774
rect 168114 97454 168734 97538
rect 168114 97218 168146 97454
rect 168382 97218 168466 97454
rect 168702 97218 168734 97454
rect 168114 61774 168734 97218
rect 168114 61538 168146 61774
rect 168382 61538 168466 61774
rect 168702 61538 168734 61774
rect 168114 61454 168734 61538
rect 168114 61218 168146 61454
rect 168382 61218 168466 61454
rect 168702 61218 168734 61454
rect 168114 25774 168734 61218
rect 168114 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 168734 25774
rect 168114 25454 168734 25538
rect 168114 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 168734 25454
rect 168114 -6106 168734 25218
rect 168114 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 168734 -6106
rect 168114 -6426 168734 -6342
rect 168114 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 168734 -6426
rect 168114 -7654 168734 -6662
rect 171834 461494 172454 478303
rect 181794 471454 182414 478303
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 171834 461258 171866 461494
rect 172102 461258 172186 461494
rect 172422 461258 172454 461494
rect 173019 461548 173085 461549
rect 173019 461484 173020 461548
rect 173084 461484 173085 461548
rect 173019 461483 173085 461484
rect 171834 461174 172454 461258
rect 171834 460938 171866 461174
rect 172102 460938 172186 461174
rect 172422 460938 172454 461174
rect 171834 425494 172454 460938
rect 171834 425258 171866 425494
rect 172102 425258 172186 425494
rect 172422 425258 172454 425494
rect 171834 425174 172454 425258
rect 171834 424938 171866 425174
rect 172102 424938 172186 425174
rect 172422 424938 172454 425174
rect 171834 389494 172454 424938
rect 171834 389258 171866 389494
rect 172102 389258 172186 389494
rect 172422 389258 172454 389494
rect 171834 389174 172454 389258
rect 171834 388938 171866 389174
rect 172102 388938 172186 389174
rect 172422 388938 172454 389174
rect 171834 353494 172454 388938
rect 171834 353258 171866 353494
rect 172102 353258 172186 353494
rect 172422 353258 172454 353494
rect 171834 353174 172454 353258
rect 171834 352938 171866 353174
rect 172102 352938 172186 353174
rect 172422 352938 172454 353174
rect 171834 317494 172454 352938
rect 171834 317258 171866 317494
rect 172102 317258 172186 317494
rect 172422 317258 172454 317494
rect 171834 317174 172454 317258
rect 171834 316938 171866 317174
rect 172102 316938 172186 317174
rect 172422 316938 172454 317174
rect 171834 281494 172454 316938
rect 171834 281258 171866 281494
rect 172102 281258 172186 281494
rect 172422 281258 172454 281494
rect 171834 281174 172454 281258
rect 171834 280938 171866 281174
rect 172102 280938 172186 281174
rect 172422 280938 172454 281174
rect 171834 245494 172454 280938
rect 173022 274685 173082 461483
rect 178539 439516 178605 439517
rect 178539 439452 178540 439516
rect 178604 439452 178605 439516
rect 178539 439451 178605 439452
rect 173203 397492 173269 397493
rect 173203 397428 173204 397492
rect 173268 397428 173269 397492
rect 173203 397427 173269 397428
rect 173206 304605 173266 397427
rect 178542 336973 178602 439451
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 178539 336972 178605 336973
rect 178539 336908 178540 336972
rect 178604 336908 178605 336972
rect 178539 336907 178605 336908
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 173203 304604 173269 304605
rect 173203 304540 173204 304604
rect 173268 304540 173269 304604
rect 173203 304539 173269 304540
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 173019 274684 173085 274685
rect 173019 274620 173020 274684
rect 173084 274620 173085 274684
rect 173019 274619 173085 274620
rect 171834 245258 171866 245494
rect 172102 245258 172186 245494
rect 172422 245258 172454 245494
rect 171834 245174 172454 245258
rect 171834 244938 171866 245174
rect 172102 244938 172186 245174
rect 172422 244938 172454 245174
rect 171834 209494 172454 244938
rect 171834 209258 171866 209494
rect 172102 209258 172186 209494
rect 172422 209258 172454 209494
rect 171834 209174 172454 209258
rect 171834 208938 171866 209174
rect 172102 208938 172186 209174
rect 172422 208938 172454 209174
rect 171834 173494 172454 208938
rect 171834 173258 171866 173494
rect 172102 173258 172186 173494
rect 172422 173258 172454 173494
rect 171834 173174 172454 173258
rect 171834 172938 171866 173174
rect 172102 172938 172186 173174
rect 172422 172938 172454 173174
rect 171834 137494 172454 172938
rect 171834 137258 171866 137494
rect 172102 137258 172186 137494
rect 172422 137258 172454 137494
rect 171834 137174 172454 137258
rect 171834 136938 171866 137174
rect 172102 136938 172186 137174
rect 172422 136938 172454 137174
rect 171834 101494 172454 136938
rect 171834 101258 171866 101494
rect 172102 101258 172186 101494
rect 172422 101258 172454 101494
rect 171834 101174 172454 101258
rect 171834 100938 171866 101174
rect 172102 100938 172186 101174
rect 172422 100938 172454 101174
rect 171834 65494 172454 100938
rect 171834 65258 171866 65494
rect 172102 65258 172186 65494
rect 172422 65258 172454 65494
rect 171834 65174 172454 65258
rect 171834 64938 171866 65174
rect 172102 64938 172186 65174
rect 172422 64938 172454 65174
rect 171834 29494 172454 64938
rect 171834 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 172454 29494
rect 171834 29174 172454 29258
rect 171834 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 172454 29174
rect 171834 -7066 172454 28938
rect 171834 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 172454 -7066
rect 171834 -7386 172454 -7302
rect 171834 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 172454 -7386
rect 171834 -7654 172454 -7622
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 185514 475174 186134 478303
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -1306 186134 6618
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -7654 186134 -1862
rect 189234 442894 189854 478303
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -2266 189854 10338
rect 189234 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 189854 -2266
rect 189234 -2586 189854 -2502
rect 189234 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 189854 -2586
rect 189234 -7654 189854 -2822
rect 192954 446614 193574 478303
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 192954 -3226 193574 14058
rect 192954 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 193574 -3226
rect 192954 -3546 193574 -3462
rect 192954 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 193574 -3546
rect 192954 -7654 193574 -3782
rect 196674 450334 197294 478303
rect 196674 450098 196706 450334
rect 196942 450098 197026 450334
rect 197262 450098 197294 450334
rect 196674 450014 197294 450098
rect 196674 449778 196706 450014
rect 196942 449778 197026 450014
rect 197262 449778 197294 450014
rect 196674 414334 197294 449778
rect 196674 414098 196706 414334
rect 196942 414098 197026 414334
rect 197262 414098 197294 414334
rect 196674 414014 197294 414098
rect 196674 413778 196706 414014
rect 196942 413778 197026 414014
rect 197262 413778 197294 414014
rect 196674 378334 197294 413778
rect 196674 378098 196706 378334
rect 196942 378098 197026 378334
rect 197262 378098 197294 378334
rect 196674 378014 197294 378098
rect 196674 377778 196706 378014
rect 196942 377778 197026 378014
rect 197262 377778 197294 378014
rect 196674 342334 197294 377778
rect 196674 342098 196706 342334
rect 196942 342098 197026 342334
rect 197262 342098 197294 342334
rect 196674 342014 197294 342098
rect 196674 341778 196706 342014
rect 196942 341778 197026 342014
rect 197262 341778 197294 342014
rect 196674 306334 197294 341778
rect 196674 306098 196706 306334
rect 196942 306098 197026 306334
rect 197262 306098 197294 306334
rect 196674 306014 197294 306098
rect 196674 305778 196706 306014
rect 196942 305778 197026 306014
rect 197262 305778 197294 306014
rect 196674 270334 197294 305778
rect 196674 270098 196706 270334
rect 196942 270098 197026 270334
rect 197262 270098 197294 270334
rect 196674 270014 197294 270098
rect 196674 269778 196706 270014
rect 196942 269778 197026 270014
rect 197262 269778 197294 270014
rect 196674 234334 197294 269778
rect 196674 234098 196706 234334
rect 196942 234098 197026 234334
rect 197262 234098 197294 234334
rect 196674 234014 197294 234098
rect 196674 233778 196706 234014
rect 196942 233778 197026 234014
rect 197262 233778 197294 234014
rect 196674 198334 197294 233778
rect 196674 198098 196706 198334
rect 196942 198098 197026 198334
rect 197262 198098 197294 198334
rect 196674 198014 197294 198098
rect 196674 197778 196706 198014
rect 196942 197778 197026 198014
rect 197262 197778 197294 198014
rect 196674 162334 197294 197778
rect 196674 162098 196706 162334
rect 196942 162098 197026 162334
rect 197262 162098 197294 162334
rect 196674 162014 197294 162098
rect 196674 161778 196706 162014
rect 196942 161778 197026 162014
rect 197262 161778 197294 162014
rect 196674 126334 197294 161778
rect 196674 126098 196706 126334
rect 196942 126098 197026 126334
rect 197262 126098 197294 126334
rect 196674 126014 197294 126098
rect 196674 125778 196706 126014
rect 196942 125778 197026 126014
rect 197262 125778 197294 126014
rect 196674 90334 197294 125778
rect 196674 90098 196706 90334
rect 196942 90098 197026 90334
rect 197262 90098 197294 90334
rect 196674 90014 197294 90098
rect 196674 89778 196706 90014
rect 196942 89778 197026 90014
rect 197262 89778 197294 90014
rect 196674 54334 197294 89778
rect 196674 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 197294 54334
rect 196674 54014 197294 54098
rect 196674 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 197294 54014
rect 196674 18334 197294 53778
rect 196674 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 197294 18334
rect 196674 18014 197294 18098
rect 196674 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 197294 18014
rect 196674 -4186 197294 17778
rect 196674 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 197294 -4186
rect 196674 -4506 197294 -4422
rect 196674 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 197294 -4506
rect 196674 -7654 197294 -4742
rect 200394 454054 201014 478303
rect 203379 476916 203445 476917
rect 203379 476852 203380 476916
rect 203444 476852 203445 476916
rect 203379 476851 203445 476852
rect 200394 453818 200426 454054
rect 200662 453818 200746 454054
rect 200982 453818 201014 454054
rect 200394 453734 201014 453818
rect 200394 453498 200426 453734
rect 200662 453498 200746 453734
rect 200982 453498 201014 453734
rect 200394 418054 201014 453498
rect 200394 417818 200426 418054
rect 200662 417818 200746 418054
rect 200982 417818 201014 418054
rect 200394 417734 201014 417818
rect 200394 417498 200426 417734
rect 200662 417498 200746 417734
rect 200982 417498 201014 417734
rect 200394 382054 201014 417498
rect 200394 381818 200426 382054
rect 200662 381818 200746 382054
rect 200982 381818 201014 382054
rect 200394 381734 201014 381818
rect 200394 381498 200426 381734
rect 200662 381498 200746 381734
rect 200982 381498 201014 381734
rect 200394 346054 201014 381498
rect 200394 345818 200426 346054
rect 200662 345818 200746 346054
rect 200982 345818 201014 346054
rect 200394 345734 201014 345818
rect 200394 345498 200426 345734
rect 200662 345498 200746 345734
rect 200982 345498 201014 345734
rect 200394 310054 201014 345498
rect 200394 309818 200426 310054
rect 200662 309818 200746 310054
rect 200982 309818 201014 310054
rect 200394 309734 201014 309818
rect 200394 309498 200426 309734
rect 200662 309498 200746 309734
rect 200982 309498 201014 309734
rect 200394 274054 201014 309498
rect 200394 273818 200426 274054
rect 200662 273818 200746 274054
rect 200982 273818 201014 274054
rect 200394 273734 201014 273818
rect 200394 273498 200426 273734
rect 200662 273498 200746 273734
rect 200982 273498 201014 273734
rect 200394 238054 201014 273498
rect 203382 272509 203442 476851
rect 204114 457774 204734 478303
rect 204114 457538 204146 457774
rect 204382 457538 204466 457774
rect 204702 457538 204734 457774
rect 204114 457454 204734 457538
rect 204114 457218 204146 457454
rect 204382 457218 204466 457454
rect 204702 457218 204734 457454
rect 204114 421774 204734 457218
rect 204114 421538 204146 421774
rect 204382 421538 204466 421774
rect 204702 421538 204734 421774
rect 204114 421454 204734 421538
rect 204114 421218 204146 421454
rect 204382 421218 204466 421454
rect 204702 421218 204734 421454
rect 204114 385774 204734 421218
rect 204114 385538 204146 385774
rect 204382 385538 204466 385774
rect 204702 385538 204734 385774
rect 204114 385454 204734 385538
rect 204114 385218 204146 385454
rect 204382 385218 204466 385454
rect 204702 385218 204734 385454
rect 204114 349774 204734 385218
rect 204114 349538 204146 349774
rect 204382 349538 204466 349774
rect 204702 349538 204734 349774
rect 204114 349454 204734 349538
rect 204114 349218 204146 349454
rect 204382 349218 204466 349454
rect 204702 349218 204734 349454
rect 204114 313774 204734 349218
rect 204114 313538 204146 313774
rect 204382 313538 204466 313774
rect 204702 313538 204734 313774
rect 204114 313454 204734 313538
rect 204114 313218 204146 313454
rect 204382 313218 204466 313454
rect 204702 313218 204734 313454
rect 204114 277774 204734 313218
rect 204114 277538 204146 277774
rect 204382 277538 204466 277774
rect 204702 277538 204734 277774
rect 204114 277454 204734 277538
rect 204114 277218 204146 277454
rect 204382 277218 204466 277454
rect 204702 277218 204734 277454
rect 203379 272508 203445 272509
rect 203379 272444 203380 272508
rect 203444 272444 203445 272508
rect 203379 272443 203445 272444
rect 200394 237818 200426 238054
rect 200662 237818 200746 238054
rect 200982 237818 201014 238054
rect 200394 237734 201014 237818
rect 200394 237498 200426 237734
rect 200662 237498 200746 237734
rect 200982 237498 201014 237734
rect 200394 202054 201014 237498
rect 200394 201818 200426 202054
rect 200662 201818 200746 202054
rect 200982 201818 201014 202054
rect 200394 201734 201014 201818
rect 200394 201498 200426 201734
rect 200662 201498 200746 201734
rect 200982 201498 201014 201734
rect 200394 166054 201014 201498
rect 200394 165818 200426 166054
rect 200662 165818 200746 166054
rect 200982 165818 201014 166054
rect 200394 165734 201014 165818
rect 200394 165498 200426 165734
rect 200662 165498 200746 165734
rect 200982 165498 201014 165734
rect 200394 130054 201014 165498
rect 200394 129818 200426 130054
rect 200662 129818 200746 130054
rect 200982 129818 201014 130054
rect 200394 129734 201014 129818
rect 200394 129498 200426 129734
rect 200662 129498 200746 129734
rect 200982 129498 201014 129734
rect 200394 94054 201014 129498
rect 200394 93818 200426 94054
rect 200662 93818 200746 94054
rect 200982 93818 201014 94054
rect 200394 93734 201014 93818
rect 200394 93498 200426 93734
rect 200662 93498 200746 93734
rect 200982 93498 201014 93734
rect 200394 58054 201014 93498
rect 200394 57818 200426 58054
rect 200662 57818 200746 58054
rect 200982 57818 201014 58054
rect 200394 57734 201014 57818
rect 200394 57498 200426 57734
rect 200662 57498 200746 57734
rect 200982 57498 201014 57734
rect 200394 22054 201014 57498
rect 200394 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 201014 22054
rect 200394 21734 201014 21818
rect 200394 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 201014 21734
rect 200394 -5146 201014 21498
rect 200394 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 201014 -5146
rect 200394 -5466 201014 -5382
rect 200394 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 201014 -5466
rect 200394 -7654 201014 -5702
rect 204114 241774 204734 277218
rect 204114 241538 204146 241774
rect 204382 241538 204466 241774
rect 204702 241538 204734 241774
rect 204114 241454 204734 241538
rect 204114 241218 204146 241454
rect 204382 241218 204466 241454
rect 204702 241218 204734 241454
rect 204114 205774 204734 241218
rect 204114 205538 204146 205774
rect 204382 205538 204466 205774
rect 204702 205538 204734 205774
rect 204114 205454 204734 205538
rect 204114 205218 204146 205454
rect 204382 205218 204466 205454
rect 204702 205218 204734 205454
rect 204114 169774 204734 205218
rect 204114 169538 204146 169774
rect 204382 169538 204466 169774
rect 204702 169538 204734 169774
rect 204114 169454 204734 169538
rect 204114 169218 204146 169454
rect 204382 169218 204466 169454
rect 204702 169218 204734 169454
rect 204114 133774 204734 169218
rect 204114 133538 204146 133774
rect 204382 133538 204466 133774
rect 204702 133538 204734 133774
rect 204114 133454 204734 133538
rect 204114 133218 204146 133454
rect 204382 133218 204466 133454
rect 204702 133218 204734 133454
rect 204114 97774 204734 133218
rect 204114 97538 204146 97774
rect 204382 97538 204466 97774
rect 204702 97538 204734 97774
rect 204114 97454 204734 97538
rect 204114 97218 204146 97454
rect 204382 97218 204466 97454
rect 204702 97218 204734 97454
rect 204114 61774 204734 97218
rect 204114 61538 204146 61774
rect 204382 61538 204466 61774
rect 204702 61538 204734 61774
rect 204114 61454 204734 61538
rect 204114 61218 204146 61454
rect 204382 61218 204466 61454
rect 204702 61218 204734 61454
rect 204114 25774 204734 61218
rect 204114 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 204734 25774
rect 204114 25454 204734 25538
rect 204114 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 204734 25454
rect 204114 -6106 204734 25218
rect 204114 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 204734 -6106
rect 204114 -6426 204734 -6342
rect 204114 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 204734 -6426
rect 204114 -7654 204734 -6662
rect 207834 461494 208454 478303
rect 217794 471454 218414 478303
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 208899 469844 208965 469845
rect 208899 469780 208900 469844
rect 208964 469780 208965 469844
rect 208899 469779 208965 469780
rect 207834 461258 207866 461494
rect 208102 461258 208186 461494
rect 208422 461258 208454 461494
rect 207834 461174 208454 461258
rect 207834 460938 207866 461174
rect 208102 460938 208186 461174
rect 208422 460938 208454 461174
rect 207834 425494 208454 460938
rect 207834 425258 207866 425494
rect 208102 425258 208186 425494
rect 208422 425258 208454 425494
rect 207834 425174 208454 425258
rect 207834 424938 207866 425174
rect 208102 424938 208186 425174
rect 208422 424938 208454 425174
rect 207834 389494 208454 424938
rect 207834 389258 207866 389494
rect 208102 389258 208186 389494
rect 208422 389258 208454 389494
rect 207834 389174 208454 389258
rect 207834 388938 207866 389174
rect 208102 388938 208186 389174
rect 208422 388938 208454 389174
rect 207834 353494 208454 388938
rect 207834 353258 207866 353494
rect 208102 353258 208186 353494
rect 208422 353258 208454 353494
rect 207834 353174 208454 353258
rect 207834 352938 207866 353174
rect 208102 352938 208186 353174
rect 208422 352938 208454 353174
rect 207834 317494 208454 352938
rect 207834 317258 207866 317494
rect 208102 317258 208186 317494
rect 208422 317258 208454 317494
rect 207834 317174 208454 317258
rect 207834 316938 207866 317174
rect 208102 316938 208186 317174
rect 208422 316938 208454 317174
rect 207834 281494 208454 316938
rect 207834 281258 207866 281494
rect 208102 281258 208186 281494
rect 208422 281258 208454 281494
rect 207834 281174 208454 281258
rect 207834 280938 207866 281174
rect 208102 280938 208186 281174
rect 208422 280938 208454 281174
rect 207834 245494 208454 280938
rect 208902 274141 208962 469779
rect 210371 456108 210437 456109
rect 210371 456044 210372 456108
rect 210436 456044 210437 456108
rect 210371 456043 210437 456044
rect 210374 302429 210434 456043
rect 217794 435454 218414 470898
rect 221514 475174 222134 478303
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 218835 441964 218901 441965
rect 218835 441900 218836 441964
rect 218900 441900 218901 441964
rect 218835 441899 218901 441900
rect 218651 441828 218717 441829
rect 218651 441764 218652 441828
rect 218716 441764 218717 441828
rect 218651 441763 218717 441764
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 210371 302428 210437 302429
rect 210371 302364 210372 302428
rect 210436 302364 210437 302428
rect 210371 302363 210437 302364
rect 217794 291454 218414 326898
rect 218654 302701 218714 441763
rect 218838 304333 218898 441899
rect 221043 441692 221109 441693
rect 221043 441628 221044 441692
rect 221108 441628 221109 441692
rect 221043 441627 221109 441628
rect 219939 441012 220005 441013
rect 219939 440948 219940 441012
rect 220004 440948 220005 441012
rect 219939 440947 220005 440948
rect 219942 333709 220002 440947
rect 219939 333708 220005 333709
rect 219939 333644 219940 333708
rect 220004 333644 220005 333708
rect 219939 333643 220005 333644
rect 218835 304332 218901 304333
rect 218835 304268 218836 304332
rect 218900 304268 218901 304332
rect 218835 304267 218901 304268
rect 218651 302700 218717 302701
rect 218651 302636 218652 302700
rect 218716 302636 218717 302700
rect 218651 302635 218717 302636
rect 221046 301069 221106 441627
rect 221227 439380 221293 439381
rect 221227 439316 221228 439380
rect 221292 439316 221293 439380
rect 221227 439315 221293 439316
rect 221043 301068 221109 301069
rect 221043 301004 221044 301068
rect 221108 301004 221109 301068
rect 221043 301003 221109 301004
rect 221230 297805 221290 439315
rect 221514 439174 222134 474618
rect 224539 472428 224605 472429
rect 224539 472364 224540 472428
rect 224604 472364 224605 472428
rect 224539 472363 224605 472364
rect 223987 442100 224053 442101
rect 223987 442036 223988 442100
rect 224052 442036 224053 442100
rect 223987 442035 224053 442036
rect 222699 440196 222765 440197
rect 222699 440132 222700 440196
rect 222764 440132 222765 440196
rect 222699 440131 222765 440132
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221227 297804 221293 297805
rect 221227 297740 221228 297804
rect 221292 297740 221293 297804
rect 221227 297739 221293 297740
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 208899 274140 208965 274141
rect 208899 274076 208900 274140
rect 208964 274076 208965 274140
rect 208899 274075 208965 274076
rect 207834 245258 207866 245494
rect 208102 245258 208186 245494
rect 208422 245258 208454 245494
rect 207834 245174 208454 245258
rect 207834 244938 207866 245174
rect 208102 244938 208186 245174
rect 208422 244938 208454 245174
rect 207834 209494 208454 244938
rect 207834 209258 207866 209494
rect 208102 209258 208186 209494
rect 208422 209258 208454 209494
rect 207834 209174 208454 209258
rect 207834 208938 207866 209174
rect 208102 208938 208186 209174
rect 208422 208938 208454 209174
rect 207834 173494 208454 208938
rect 207834 173258 207866 173494
rect 208102 173258 208186 173494
rect 208422 173258 208454 173494
rect 207834 173174 208454 173258
rect 207834 172938 207866 173174
rect 208102 172938 208186 173174
rect 208422 172938 208454 173174
rect 207834 137494 208454 172938
rect 207834 137258 207866 137494
rect 208102 137258 208186 137494
rect 208422 137258 208454 137494
rect 207834 137174 208454 137258
rect 207834 136938 207866 137174
rect 208102 136938 208186 137174
rect 208422 136938 208454 137174
rect 207834 101494 208454 136938
rect 207834 101258 207866 101494
rect 208102 101258 208186 101494
rect 208422 101258 208454 101494
rect 207834 101174 208454 101258
rect 207834 100938 207866 101174
rect 208102 100938 208186 101174
rect 208422 100938 208454 101174
rect 207834 65494 208454 100938
rect 207834 65258 207866 65494
rect 208102 65258 208186 65494
rect 208422 65258 208454 65494
rect 207834 65174 208454 65258
rect 207834 64938 207866 65174
rect 208102 64938 208186 65174
rect 208422 64938 208454 65174
rect 207834 29494 208454 64938
rect 207834 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 208454 29494
rect 207834 29174 208454 29258
rect 207834 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 208454 29174
rect 207834 -7066 208454 28938
rect 207834 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 208454 -7066
rect 207834 -7386 208454 -7302
rect 207834 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 208454 -7386
rect 207834 -7654 208454 -7622
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 221514 295174 222134 330618
rect 222702 327181 222762 440131
rect 223990 410549 224050 442035
rect 224171 439788 224237 439789
rect 224171 439724 224172 439788
rect 224236 439724 224237 439788
rect 224171 439723 224237 439724
rect 223987 410548 224053 410549
rect 223987 410484 223988 410548
rect 224052 410484 224053 410548
rect 223987 410483 224053 410484
rect 223067 344724 223133 344725
rect 223067 344660 223068 344724
rect 223132 344660 223133 344724
rect 223067 344659 223133 344660
rect 222699 327180 222765 327181
rect 222699 327116 222700 327180
rect 222764 327116 222765 327180
rect 222699 327115 222765 327116
rect 222699 308956 222765 308957
rect 222699 308892 222700 308956
rect 222764 308892 222765 308956
rect 222699 308891 222765 308892
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 223174 222134 258618
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 222702 7581 222762 308891
rect 223070 273053 223130 344659
rect 224174 328813 224234 439723
rect 224355 410004 224421 410005
rect 224355 409940 224356 410004
rect 224420 409940 224421 410004
rect 224355 409939 224421 409940
rect 224171 328812 224237 328813
rect 224171 328748 224172 328812
rect 224236 328748 224237 328812
rect 224171 328747 224237 328748
rect 224358 318205 224418 409939
rect 224355 318204 224421 318205
rect 224355 318140 224356 318204
rect 224420 318140 224421 318204
rect 224355 318139 224421 318140
rect 224542 316573 224602 472363
rect 224723 472020 224789 472021
rect 224723 471956 224724 472020
rect 224788 471956 224789 472020
rect 224723 471955 224789 471956
rect 224539 316572 224605 316573
rect 224539 316508 224540 316572
rect 224604 316508 224605 316572
rect 224539 316507 224605 316508
rect 224726 315485 224786 471955
rect 225234 442894 225854 478303
rect 227667 449580 227733 449581
rect 227667 449516 227668 449580
rect 227732 449516 227733 449580
rect 227667 449515 227733 449516
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 224907 442372 224973 442373
rect 224907 442308 224908 442372
rect 224972 442370 224973 442372
rect 224972 442310 225154 442370
rect 224972 442308 224973 442310
rect 224907 442307 224973 442308
rect 225094 437490 225154 442310
rect 224910 437430 225154 437490
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 224723 315484 224789 315485
rect 224723 315420 224724 315484
rect 224788 315420 224789 315484
rect 224723 315419 224789 315420
rect 224171 308412 224237 308413
rect 224171 308348 224172 308412
rect 224236 308348 224237 308412
rect 224171 308347 224237 308348
rect 223067 273052 223133 273053
rect 223067 272988 223068 273052
rect 223132 272988 223133 273052
rect 223067 272987 223133 272988
rect 224174 45525 224234 308347
rect 224910 296173 224970 437430
rect 225234 406894 225854 442338
rect 226931 441420 226997 441421
rect 226931 441356 226932 441420
rect 226996 441356 226997 441420
rect 226931 441355 226997 441356
rect 226195 440332 226261 440333
rect 226195 440268 226196 440332
rect 226260 440268 226261 440332
rect 226195 440267 226261 440268
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 224907 296172 224973 296173
rect 224907 296108 224908 296172
rect 224972 296108 224973 296172
rect 224907 296107 224973 296108
rect 224907 295356 224973 295357
rect 224907 295292 224908 295356
rect 224972 295292 224973 295356
rect 224907 295291 224973 295292
rect 224910 286381 224970 295291
rect 224907 286380 224973 286381
rect 224907 286316 224908 286380
rect 224972 286316 224973 286380
rect 224907 286315 224973 286316
rect 225234 262894 225854 298338
rect 226198 284749 226258 440267
rect 226934 322285 226994 441355
rect 227670 440197 227730 449515
rect 228954 446614 229574 478303
rect 232267 478140 232333 478141
rect 232267 478076 232268 478140
rect 232332 478076 232333 478140
rect 232267 478075 232333 478076
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228403 441556 228469 441557
rect 228403 441492 228404 441556
rect 228468 441492 228469 441556
rect 228403 441491 228469 441492
rect 227851 440332 227917 440333
rect 227851 440268 227852 440332
rect 227916 440268 227917 440332
rect 227851 440267 227917 440268
rect 227667 440196 227733 440197
rect 227667 440132 227668 440196
rect 227732 440132 227733 440196
rect 227667 440131 227733 440132
rect 227115 439652 227181 439653
rect 227115 439588 227116 439652
rect 227180 439588 227181 439652
rect 227115 439587 227181 439588
rect 227118 330445 227178 439587
rect 227667 439244 227733 439245
rect 227667 439180 227668 439244
rect 227732 439180 227733 439244
rect 227667 439179 227733 439180
rect 227115 330444 227181 330445
rect 227115 330380 227116 330444
rect 227180 330380 227181 330444
rect 227115 330379 227181 330380
rect 226931 322284 226997 322285
rect 226931 322220 226932 322284
rect 226996 322220 226997 322284
rect 226931 322219 226997 322220
rect 227670 291277 227730 439179
rect 227854 292909 227914 440267
rect 228219 439924 228285 439925
rect 228219 439860 228220 439924
rect 228284 439860 228285 439924
rect 228219 439859 228285 439860
rect 228035 331396 228101 331397
rect 228035 331332 228036 331396
rect 228100 331332 228101 331396
rect 228035 331331 228101 331332
rect 228038 294541 228098 331331
rect 228222 315757 228282 439859
rect 228406 332077 228466 441491
rect 228954 410614 229574 446058
rect 230979 441148 231045 441149
rect 230979 441084 230980 441148
rect 231044 441084 231045 441148
rect 230979 441083 231045 441084
rect 230059 441012 230125 441013
rect 230059 440948 230060 441012
rect 230124 440948 230125 441012
rect 230059 440947 230125 440948
rect 229875 439108 229941 439109
rect 229875 439044 229876 439108
rect 229940 439044 229941 439108
rect 229875 439043 229941 439044
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228403 332076 228469 332077
rect 228403 332012 228404 332076
rect 228468 332012 228469 332076
rect 228403 332011 228469 332012
rect 228219 315756 228285 315757
rect 228219 315692 228220 315756
rect 228284 315692 228285 315756
rect 228219 315691 228285 315692
rect 228219 306780 228285 306781
rect 228219 306716 228220 306780
rect 228284 306716 228285 306780
rect 228219 306715 228285 306716
rect 228035 294540 228101 294541
rect 228035 294476 228036 294540
rect 228100 294476 228101 294540
rect 228035 294475 228101 294476
rect 227851 292908 227917 292909
rect 227851 292844 227852 292908
rect 227916 292844 227917 292908
rect 227851 292843 227917 292844
rect 227667 291276 227733 291277
rect 227667 291212 227668 291276
rect 227732 291212 227733 291276
rect 227667 291211 227733 291212
rect 226195 284748 226261 284749
rect 226195 284684 226196 284748
rect 226260 284684 226261 284748
rect 226195 284683 226261 284684
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 226894 225854 262338
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 154894 225854 190338
rect 228222 188869 228282 306715
rect 228954 302614 229574 338058
rect 229878 317389 229938 439043
rect 230062 335341 230122 440947
rect 230427 440332 230493 440333
rect 230427 440268 230428 440332
rect 230492 440268 230493 440332
rect 230427 440267 230493 440268
rect 230059 335340 230125 335341
rect 230059 335276 230060 335340
rect 230124 335276 230125 335340
rect 230059 335275 230125 335276
rect 230243 334116 230309 334117
rect 230243 334052 230244 334116
rect 230308 334052 230309 334116
rect 230243 334051 230309 334052
rect 229875 317388 229941 317389
rect 229875 317324 229876 317388
rect 229940 317324 229941 317388
rect 229875 317323 229941 317324
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 266614 229574 302058
rect 230246 294813 230306 334051
rect 230430 310861 230490 440267
rect 230611 324460 230677 324461
rect 230611 324396 230612 324460
rect 230676 324396 230677 324460
rect 230611 324395 230677 324396
rect 230427 310860 230493 310861
rect 230427 310796 230428 310860
rect 230492 310796 230493 310860
rect 230427 310795 230493 310796
rect 230243 294812 230309 294813
rect 230243 294748 230244 294812
rect 230308 294748 230309 294812
rect 230243 294747 230309 294748
rect 230614 289645 230674 324395
rect 230982 319021 231042 441083
rect 231899 440332 231965 440333
rect 231899 440268 231900 440332
rect 231964 440268 231965 440332
rect 231899 440267 231965 440268
rect 231531 439380 231597 439381
rect 231531 439316 231532 439380
rect 231596 439316 231597 439380
rect 231531 439315 231597 439316
rect 231163 438564 231229 438565
rect 231163 438500 231164 438564
rect 231228 438500 231229 438564
rect 231163 438499 231229 438500
rect 230979 319020 231045 319021
rect 230979 318956 230980 319020
rect 231044 318956 231045 319020
rect 230979 318955 231045 318956
rect 230979 307868 231045 307869
rect 230979 307804 230980 307868
rect 231044 307804 231045 307868
rect 230979 307803 231045 307804
rect 230611 289644 230677 289645
rect 230611 289580 230612 289644
rect 230676 289580 230677 289644
rect 230611 289579 230677 289580
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 230614 229574 266058
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228219 188868 228285 188869
rect 228219 188804 228220 188868
rect 228284 188804 228285 188868
rect 228219 188803 228285 188804
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 118894 225854 154338
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 82894 225854 118338
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 224171 45524 224237 45525
rect 224171 45460 224172 45524
rect 224236 45460 224237 45524
rect 224171 45459 224237 45460
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 222699 7580 222765 7581
rect 222699 7516 222700 7580
rect 222764 7516 222765 7580
rect 222699 7515 222765 7516
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -7654 222134 -1862
rect 225234 -2266 225854 10338
rect 225234 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 225854 -2266
rect 225234 -2586 225854 -2502
rect 225234 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 225854 -2586
rect 225234 -7654 225854 -2822
rect 228954 158614 229574 194058
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 230982 86325 231042 307803
rect 231166 288013 231226 438499
rect 231534 325549 231594 439315
rect 231531 325548 231597 325549
rect 231531 325484 231532 325548
rect 231596 325484 231597 325548
rect 231531 325483 231597 325484
rect 231902 314125 231962 440267
rect 231899 314124 231965 314125
rect 231899 314060 231900 314124
rect 231964 314060 231965 314124
rect 231899 314059 231965 314060
rect 232083 313308 232149 313309
rect 232083 313244 232084 313308
rect 232148 313244 232149 313308
rect 232083 313243 232149 313244
rect 231347 306236 231413 306237
rect 231347 306172 231348 306236
rect 231412 306172 231413 306236
rect 231347 306171 231413 306172
rect 231163 288012 231229 288013
rect 231163 287948 231164 288012
rect 231228 287948 231229 288012
rect 231163 287947 231229 287948
rect 231350 242181 231410 306171
rect 232086 295901 232146 313243
rect 232083 295900 232149 295901
rect 232083 295836 232084 295900
rect 232148 295836 232149 295900
rect 232083 295835 232149 295836
rect 232270 294269 232330 478075
rect 232674 450334 233294 478303
rect 234291 474060 234357 474061
rect 234291 473996 234292 474060
rect 234356 473996 234357 474060
rect 234291 473995 234357 473996
rect 234107 450532 234173 450533
rect 234107 450468 234108 450532
rect 234172 450468 234173 450532
rect 234107 450467 234173 450468
rect 232674 450098 232706 450334
rect 232942 450098 233026 450334
rect 233262 450098 233294 450334
rect 232674 450014 233294 450098
rect 232674 449778 232706 450014
rect 232942 449778 233026 450014
rect 233262 449778 233294 450014
rect 232674 414334 233294 449778
rect 233923 441692 233989 441693
rect 233923 441628 233924 441692
rect 233988 441628 233989 441692
rect 233923 441627 233989 441628
rect 232674 414098 232706 414334
rect 232942 414098 233026 414334
rect 233262 414098 233294 414334
rect 232674 414014 233294 414098
rect 232674 413778 232706 414014
rect 232942 413778 233026 414014
rect 233262 413778 233294 414014
rect 232674 378334 233294 413778
rect 232674 378098 232706 378334
rect 232942 378098 233026 378334
rect 233262 378098 233294 378334
rect 232674 378014 233294 378098
rect 232674 377778 232706 378014
rect 232942 377778 233026 378014
rect 233262 377778 233294 378014
rect 232674 342334 233294 377778
rect 232674 342098 232706 342334
rect 232942 342098 233026 342334
rect 233262 342098 233294 342334
rect 232674 342014 233294 342098
rect 232674 341778 232706 342014
rect 232942 341778 233026 342014
rect 233262 341778 233294 342014
rect 232674 306334 233294 341778
rect 233926 309501 233986 441627
rect 234110 311677 234170 450467
rect 234107 311676 234173 311677
rect 234107 311612 234108 311676
rect 234172 311612 234173 311676
rect 234107 311611 234173 311612
rect 234294 311133 234354 473995
rect 234291 311132 234357 311133
rect 234291 311068 234292 311132
rect 234356 311068 234357 311132
rect 234291 311067 234357 311068
rect 234478 310589 234538 479435
rect 235763 458828 235829 458829
rect 235763 458764 235764 458828
rect 235828 458764 235829 458828
rect 235763 458763 235829 458764
rect 235579 446588 235645 446589
rect 235579 446524 235580 446588
rect 235644 446524 235645 446588
rect 235579 446523 235645 446524
rect 235211 444140 235277 444141
rect 235211 444076 235212 444140
rect 235276 444076 235277 444140
rect 235211 444075 235277 444076
rect 234659 341732 234725 341733
rect 234659 341668 234660 341732
rect 234724 341668 234725 341732
rect 234659 341667 234725 341668
rect 234475 310588 234541 310589
rect 234475 310524 234476 310588
rect 234540 310524 234541 310588
rect 234475 310523 234541 310524
rect 233923 309500 233989 309501
rect 233923 309436 233924 309500
rect 233988 309436 233989 309500
rect 233923 309435 233989 309436
rect 234662 307733 234722 341667
rect 235027 341596 235093 341597
rect 235027 341532 235028 341596
rect 235092 341532 235093 341596
rect 235027 341531 235093 341532
rect 234659 307732 234725 307733
rect 234659 307668 234660 307732
rect 234724 307668 234725 307732
rect 234659 307667 234725 307668
rect 232674 306098 232706 306334
rect 232942 306098 233026 306334
rect 233262 306098 233294 306334
rect 232674 306014 233294 306098
rect 232674 305778 232706 306014
rect 232942 305778 233026 306014
rect 233262 305778 233294 306014
rect 232267 294268 232333 294269
rect 232267 294204 232268 294268
rect 232332 294204 232333 294268
rect 232267 294203 232333 294204
rect 232674 270334 233294 305778
rect 235030 276861 235090 341531
rect 235214 341053 235274 444075
rect 235582 368797 235642 446523
rect 235579 368796 235645 368797
rect 235579 368732 235580 368796
rect 235644 368732 235645 368796
rect 235579 368731 235645 368732
rect 235395 358460 235461 358461
rect 235395 358396 235396 358460
rect 235460 358396 235461 358460
rect 235395 358395 235461 358396
rect 235211 341052 235277 341053
rect 235211 340988 235212 341052
rect 235276 340988 235277 341052
rect 235211 340987 235277 340988
rect 235211 307324 235277 307325
rect 235211 307260 235212 307324
rect 235276 307260 235277 307324
rect 235211 307259 235277 307260
rect 235027 276860 235093 276861
rect 235027 276796 235028 276860
rect 235092 276796 235093 276860
rect 235027 276795 235093 276796
rect 232674 270098 232706 270334
rect 232942 270098 233026 270334
rect 233262 270098 233294 270334
rect 232674 270014 233294 270098
rect 232674 269778 232706 270014
rect 232942 269778 233026 270014
rect 233262 269778 233294 270014
rect 231347 242180 231413 242181
rect 231347 242116 231348 242180
rect 231412 242116 231413 242180
rect 231347 242115 231413 242116
rect 232674 234334 233294 269778
rect 232674 234098 232706 234334
rect 232942 234098 233026 234334
rect 233262 234098 233294 234334
rect 232674 234014 233294 234098
rect 232674 233778 232706 234014
rect 232942 233778 233026 234014
rect 233262 233778 233294 234014
rect 232674 198334 233294 233778
rect 232674 198098 232706 198334
rect 232942 198098 233026 198334
rect 233262 198098 233294 198334
rect 232674 198014 233294 198098
rect 232674 197778 232706 198014
rect 232942 197778 233026 198014
rect 233262 197778 233294 198014
rect 232674 162334 233294 197778
rect 232674 162098 232706 162334
rect 232942 162098 233026 162334
rect 233262 162098 233294 162334
rect 232674 162014 233294 162098
rect 232674 161778 232706 162014
rect 232942 161778 233026 162014
rect 233262 161778 233294 162014
rect 232674 126334 233294 161778
rect 235214 136781 235274 307259
rect 235398 240549 235458 358395
rect 235579 341460 235645 341461
rect 235579 341396 235580 341460
rect 235644 341396 235645 341460
rect 235579 341395 235645 341396
rect 235582 271421 235642 341395
rect 235766 340917 235826 458763
rect 236394 454054 237014 478303
rect 239811 476780 239877 476781
rect 239811 476716 239812 476780
rect 239876 476716 239877 476780
rect 239811 476715 239877 476716
rect 238339 472020 238405 472021
rect 238339 471956 238340 472020
rect 238404 471956 238405 472020
rect 238339 471955 238405 471956
rect 238155 456108 238221 456109
rect 238155 456044 238156 456108
rect 238220 456044 238221 456108
rect 238155 456043 238221 456044
rect 236394 453818 236426 454054
rect 236662 453818 236746 454054
rect 236982 453818 237014 454054
rect 236394 453734 237014 453818
rect 236394 453498 236426 453734
rect 236662 453498 236746 453734
rect 236982 453498 237014 453734
rect 236394 418054 237014 453498
rect 237235 449580 237301 449581
rect 237235 449516 237236 449580
rect 237300 449516 237301 449580
rect 237235 449515 237301 449516
rect 236394 417818 236426 418054
rect 236662 417818 236746 418054
rect 236982 417818 237014 418054
rect 236394 417734 237014 417818
rect 236394 417498 236426 417734
rect 236662 417498 236746 417734
rect 236982 417498 237014 417734
rect 236394 382054 237014 417498
rect 236394 381818 236426 382054
rect 236662 381818 236746 382054
rect 236982 381818 237014 382054
rect 236394 381734 237014 381818
rect 236394 381498 236426 381734
rect 236662 381498 236746 381734
rect 236982 381498 237014 381734
rect 236394 346054 237014 381498
rect 236394 345818 236426 346054
rect 236662 345818 236746 346054
rect 236982 345818 237014 346054
rect 236394 345734 237014 345818
rect 236394 345498 236426 345734
rect 236662 345498 236746 345734
rect 236982 345498 237014 345734
rect 235763 340916 235829 340917
rect 235763 340852 235764 340916
rect 235828 340852 235829 340916
rect 235763 340851 235829 340852
rect 236394 310054 237014 345498
rect 236394 309818 236426 310054
rect 236662 309818 236746 310054
rect 236982 309818 237014 310054
rect 236394 309734 237014 309818
rect 236394 309498 236426 309734
rect 236662 309498 236746 309734
rect 236982 309498 237014 309734
rect 236394 274054 237014 309498
rect 237238 298077 237298 449515
rect 237971 449308 238037 449309
rect 237971 449244 237972 449308
rect 238036 449244 238037 449308
rect 237971 449243 238037 449244
rect 237974 347717 238034 449243
rect 237971 347716 238037 347717
rect 237971 347652 237972 347716
rect 238036 347652 238037 347716
rect 237971 347651 238037 347652
rect 237419 347172 237485 347173
rect 237419 347108 237420 347172
rect 237484 347108 237485 347172
rect 237419 347107 237485 347108
rect 237235 298076 237301 298077
rect 237235 298012 237236 298076
rect 237300 298012 237301 298076
rect 237235 298011 237301 298012
rect 237422 282981 237482 347107
rect 238158 316029 238218 456043
rect 238342 317117 238402 471955
rect 238523 468484 238589 468485
rect 238523 468420 238524 468484
rect 238588 468420 238589 468484
rect 238523 468419 238589 468420
rect 238339 317116 238405 317117
rect 238339 317052 238340 317116
rect 238404 317052 238405 317116
rect 238339 317051 238405 317052
rect 238339 316980 238405 316981
rect 238339 316916 238340 316980
rect 238404 316916 238405 316980
rect 238339 316915 238405 316916
rect 238155 316028 238221 316029
rect 238155 315964 238156 316028
rect 238220 315964 238221 316028
rect 238155 315963 238221 315964
rect 238342 295357 238402 316915
rect 238526 310045 238586 468419
rect 239627 439108 239693 439109
rect 239627 439044 239628 439108
rect 239692 439044 239693 439108
rect 239627 439043 239693 439044
rect 239443 406060 239509 406061
rect 239443 405996 239444 406060
rect 239508 405996 239509 406060
rect 239443 405995 239509 405996
rect 239446 326365 239506 405995
rect 239443 326364 239509 326365
rect 239443 326300 239444 326364
rect 239508 326300 239509 326364
rect 239443 326299 239509 326300
rect 238523 310044 238589 310045
rect 238523 309980 238524 310044
rect 238588 309980 238589 310044
rect 238523 309979 238589 309980
rect 238339 295356 238405 295357
rect 238339 295292 238340 295356
rect 238404 295292 238405 295356
rect 238339 295291 238405 295292
rect 239630 293725 239690 439043
rect 239814 323101 239874 476715
rect 240114 457774 240734 478303
rect 240915 477868 240981 477869
rect 240915 477804 240916 477868
rect 240980 477804 240981 477868
rect 240915 477803 240981 477804
rect 240114 457538 240146 457774
rect 240382 457538 240466 457774
rect 240702 457538 240734 457774
rect 240114 457454 240734 457538
rect 240114 457218 240146 457454
rect 240382 457218 240466 457454
rect 240702 457218 240734 457454
rect 240114 421774 240734 457218
rect 240114 421538 240146 421774
rect 240382 421538 240466 421774
rect 240702 421538 240734 421774
rect 240114 421454 240734 421538
rect 240114 421218 240146 421454
rect 240382 421218 240466 421454
rect 240702 421218 240734 421454
rect 240114 402313 240734 421218
rect 240179 401572 240245 401573
rect 240179 401508 240180 401572
rect 240244 401570 240245 401572
rect 240918 401570 240978 477803
rect 253794 471454 254414 478303
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 244208 435454 244528 435486
rect 244208 435218 244250 435454
rect 244486 435218 244528 435454
rect 244208 435134 244528 435218
rect 244208 434898 244250 435134
rect 244486 434898 244528 435134
rect 244208 434866 244528 434898
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 402313 254414 434898
rect 257514 475174 258134 478303
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 261234 442894 261854 478303
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 402313 258134 402618
rect 259568 403174 259888 403206
rect 259568 402938 259610 403174
rect 259846 402938 259888 403174
rect 259568 402854 259888 402938
rect 259568 402618 259610 402854
rect 259846 402618 259888 402854
rect 259568 402586 259888 402618
rect 261234 402313 261854 406338
rect 264954 446614 265574 478303
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 402313 265574 410058
rect 268674 450334 269294 478303
rect 268674 450098 268706 450334
rect 268942 450098 269026 450334
rect 269262 450098 269294 450334
rect 268674 450014 269294 450098
rect 268674 449778 268706 450014
rect 268942 449778 269026 450014
rect 269262 449778 269294 450014
rect 268674 414334 269294 449778
rect 268674 414098 268706 414334
rect 268942 414098 269026 414334
rect 269262 414098 269294 414334
rect 268674 414014 269294 414098
rect 268674 413778 268706 414014
rect 268942 413778 269026 414014
rect 269262 413778 269294 414014
rect 268674 402313 269294 413778
rect 272394 454054 273014 478303
rect 272394 453818 272426 454054
rect 272662 453818 272746 454054
rect 272982 453818 273014 454054
rect 272394 453734 273014 453818
rect 272394 453498 272426 453734
rect 272662 453498 272746 453734
rect 272982 453498 273014 453734
rect 272394 418054 273014 453498
rect 276114 457774 276734 478303
rect 276114 457538 276146 457774
rect 276382 457538 276466 457774
rect 276702 457538 276734 457774
rect 276114 457454 276734 457538
rect 276114 457218 276146 457454
rect 276382 457218 276466 457454
rect 276702 457218 276734 457454
rect 274928 435454 275248 435486
rect 274928 435218 274970 435454
rect 275206 435218 275248 435454
rect 274928 435134 275248 435218
rect 274928 434898 274970 435134
rect 275206 434898 275248 435134
rect 274928 434866 275248 434898
rect 272394 417818 272426 418054
rect 272662 417818 272746 418054
rect 272982 417818 273014 418054
rect 272394 417734 273014 417818
rect 272394 417498 272426 417734
rect 272662 417498 272746 417734
rect 272982 417498 273014 417734
rect 272394 402313 273014 417498
rect 276114 421774 276734 457218
rect 279834 461494 280454 478303
rect 289310 471477 289370 516155
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289307 471476 289373 471477
rect 289307 471412 289308 471476
rect 289372 471412 289373 471476
rect 289307 471411 289373 471412
rect 289794 471454 290414 506898
rect 290598 480181 290658 622235
rect 290779 581500 290845 581501
rect 290779 581436 290780 581500
rect 290844 581436 290845 581500
rect 290779 581435 290845 581436
rect 290595 480180 290661 480181
rect 290595 480116 290596 480180
rect 290660 480116 290661 480180
rect 290595 480115 290661 480116
rect 290782 480045 290842 581435
rect 290779 480044 290845 480045
rect 290779 479980 290780 480044
rect 290844 479980 290845 480044
rect 290779 479979 290845 479980
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 282867 467396 282933 467397
rect 282867 467332 282868 467396
rect 282932 467332 282933 467396
rect 282867 467331 282933 467332
rect 279834 461258 279866 461494
rect 280102 461258 280186 461494
rect 280422 461258 280454 461494
rect 279834 461174 280454 461258
rect 279834 460938 279866 461174
rect 280102 460938 280186 461174
rect 280422 460938 280454 461174
rect 278819 440468 278885 440469
rect 278819 440404 278820 440468
rect 278884 440404 278885 440468
rect 278819 440403 278885 440404
rect 278822 438701 278882 440403
rect 279371 438972 279437 438973
rect 279371 438908 279372 438972
rect 279436 438908 279437 438972
rect 279371 438907 279437 438908
rect 278819 438700 278885 438701
rect 278819 438636 278820 438700
rect 278884 438636 278885 438700
rect 278819 438635 278885 438636
rect 279374 437477 279434 438907
rect 279555 438564 279621 438565
rect 279555 438500 279556 438564
rect 279620 438500 279621 438564
rect 279555 438499 279621 438500
rect 279371 437476 279437 437477
rect 279371 437412 279372 437476
rect 279436 437412 279437 437476
rect 279371 437411 279437 437412
rect 276114 421538 276146 421774
rect 276382 421538 276466 421774
rect 276702 421538 276734 421774
rect 276114 421454 276734 421538
rect 276114 421218 276146 421454
rect 276382 421218 276466 421454
rect 276702 421218 276734 421454
rect 276114 402313 276734 421218
rect 240244 401510 240978 401570
rect 240244 401508 240245 401510
rect 240179 401507 240245 401508
rect 244208 399454 244528 399486
rect 244208 399218 244250 399454
rect 244486 399218 244528 399454
rect 244208 399134 244528 399218
rect 244208 398898 244250 399134
rect 244486 398898 244528 399134
rect 244208 398866 244528 398898
rect 274928 399454 275248 399486
rect 274928 399218 274970 399454
rect 275206 399218 275248 399454
rect 274928 399134 275248 399218
rect 274928 398898 274970 399134
rect 275206 398898 275248 399134
rect 274928 398866 275248 398898
rect 279558 396269 279618 438499
rect 279834 425494 280454 460938
rect 280659 441284 280725 441285
rect 280659 441220 280660 441284
rect 280724 441220 280725 441284
rect 280659 441219 280725 441220
rect 279834 425258 279866 425494
rect 280102 425258 280186 425494
rect 280422 425258 280454 425494
rect 279834 425174 280454 425258
rect 279834 424938 279866 425174
rect 280102 424938 280186 425174
rect 280422 424938 280454 425174
rect 279555 396268 279621 396269
rect 279555 396204 279556 396268
rect 279620 396204 279621 396268
rect 279555 396203 279621 396204
rect 279834 389494 280454 424938
rect 280662 423469 280722 441219
rect 281947 439924 282013 439925
rect 281947 439860 281948 439924
rect 282012 439860 282013 439924
rect 281947 439859 282013 439860
rect 281763 439788 281829 439789
rect 281763 439724 281764 439788
rect 281828 439724 281829 439788
rect 281763 439723 281829 439724
rect 280843 438972 280909 438973
rect 280843 438908 280844 438972
rect 280908 438908 280909 438972
rect 280843 438907 280909 438908
rect 280846 426189 280906 438907
rect 281766 430269 281826 439723
rect 281950 431629 282010 439859
rect 282315 439652 282381 439653
rect 282315 439588 282316 439652
rect 282380 439588 282381 439652
rect 282315 439587 282381 439588
rect 281947 431628 282013 431629
rect 281947 431564 281948 431628
rect 282012 431564 282013 431628
rect 281947 431563 282013 431564
rect 281763 430268 281829 430269
rect 281763 430204 281764 430268
rect 281828 430204 281829 430268
rect 281763 430203 281829 430204
rect 282318 428909 282378 439587
rect 282315 428908 282381 428909
rect 282315 428844 282316 428908
rect 282380 428844 282381 428908
rect 282315 428843 282381 428844
rect 280843 426188 280909 426189
rect 280843 426124 280844 426188
rect 280908 426124 280909 426188
rect 280843 426123 280909 426124
rect 280659 423468 280725 423469
rect 280659 423404 280660 423468
rect 280724 423404 280725 423468
rect 280659 423403 280725 423404
rect 279834 389258 279866 389494
rect 280102 389258 280186 389494
rect 280422 389258 280454 389494
rect 279834 389174 280454 389258
rect 279834 388938 279866 389174
rect 280102 388938 280186 389174
rect 280422 388938 280454 389174
rect 259568 367174 259888 367206
rect 259568 366938 259610 367174
rect 259846 366938 259888 367174
rect 259568 366854 259888 366938
rect 259568 366618 259610 366854
rect 259846 366618 259888 366854
rect 259568 366586 259888 366618
rect 244208 363454 244528 363486
rect 244208 363218 244250 363454
rect 244486 363218 244528 363454
rect 244208 363134 244528 363218
rect 244208 362898 244250 363134
rect 244486 362898 244528 363134
rect 244208 362866 244528 362898
rect 274928 363454 275248 363486
rect 274928 363218 274970 363454
rect 275206 363218 275248 363454
rect 274928 363134 275248 363218
rect 274928 362898 274970 363134
rect 275206 362898 275248 363134
rect 274928 362866 275248 362898
rect 279834 353494 280454 388938
rect 279834 353258 279866 353494
rect 280102 353258 280186 353494
rect 280422 353258 280454 353494
rect 279834 353174 280454 353258
rect 279834 352938 279866 353174
rect 280102 352938 280186 353174
rect 280422 352938 280454 353174
rect 259568 331174 259888 331206
rect 259568 330938 259610 331174
rect 259846 330938 259888 331174
rect 259568 330854 259888 330938
rect 259568 330618 259610 330854
rect 259846 330618 259888 330854
rect 259568 330586 259888 330618
rect 244208 327454 244528 327486
rect 244208 327218 244250 327454
rect 244486 327218 244528 327454
rect 244208 327134 244528 327218
rect 244208 326898 244250 327134
rect 244486 326898 244528 327134
rect 244208 326866 244528 326898
rect 274928 327454 275248 327486
rect 274928 327218 274970 327454
rect 275206 327218 275248 327454
rect 274928 327134 275248 327218
rect 274928 326898 274970 327134
rect 275206 326898 275248 327134
rect 274928 326866 275248 326898
rect 239811 323100 239877 323101
rect 239811 323036 239812 323100
rect 239876 323036 239877 323100
rect 239811 323035 239877 323036
rect 279834 317494 280454 352938
rect 280843 339148 280909 339149
rect 280843 339084 280844 339148
rect 280908 339084 280909 339148
rect 280843 339083 280909 339084
rect 279834 317258 279866 317494
rect 280102 317258 280186 317494
rect 280422 317258 280454 317494
rect 279834 317174 280454 317258
rect 279834 316938 279866 317174
rect 280102 316938 280186 317174
rect 280422 316938 280454 317174
rect 279371 303788 279437 303789
rect 279371 303724 279372 303788
rect 279436 303724 279437 303788
rect 279371 303723 279437 303724
rect 259568 295174 259888 295206
rect 259568 294938 259610 295174
rect 259846 294938 259888 295174
rect 259568 294854 259888 294938
rect 259568 294618 259610 294854
rect 259846 294618 259888 294854
rect 259568 294586 259888 294618
rect 239627 293724 239693 293725
rect 239627 293660 239628 293724
rect 239692 293660 239693 293724
rect 239627 293659 239693 293660
rect 238155 293180 238221 293181
rect 238155 293116 238156 293180
rect 238220 293116 238221 293180
rect 238155 293115 238221 293116
rect 237971 283116 238037 283117
rect 237971 283052 237972 283116
rect 238036 283052 238037 283116
rect 237971 283051 238037 283052
rect 237419 282980 237485 282981
rect 237419 282916 237420 282980
rect 237484 282916 237485 282980
rect 237419 282915 237485 282916
rect 237787 281484 237853 281485
rect 237787 281420 237788 281484
rect 237852 281420 237853 281484
rect 237787 281419 237853 281420
rect 236394 273818 236426 274054
rect 236662 273818 236746 274054
rect 236982 273818 237014 274054
rect 236394 273734 237014 273818
rect 236394 273498 236426 273734
rect 236662 273498 236746 273734
rect 236982 273498 237014 273734
rect 235579 271420 235645 271421
rect 235579 271356 235580 271420
rect 235644 271356 235645 271420
rect 235579 271355 235645 271356
rect 235395 240548 235461 240549
rect 235395 240484 235396 240548
rect 235460 240484 235461 240548
rect 235395 240483 235461 240484
rect 236394 238054 237014 273498
rect 237790 240413 237850 281419
rect 237787 240412 237853 240413
rect 237787 240348 237788 240412
rect 237852 240348 237853 240412
rect 237787 240347 237853 240348
rect 237974 239733 238034 283051
rect 238158 281485 238218 293115
rect 238523 292636 238589 292637
rect 238523 292572 238524 292636
rect 238588 292572 238589 292636
rect 238523 292571 238589 292572
rect 238339 292092 238405 292093
rect 238339 292028 238340 292092
rect 238404 292028 238405 292092
rect 238339 292027 238405 292028
rect 238155 281484 238221 281485
rect 238155 281420 238156 281484
rect 238220 281420 238221 281484
rect 238155 281419 238221 281420
rect 237971 239732 238037 239733
rect 237971 239668 237972 239732
rect 238036 239668 238037 239732
rect 237971 239667 238037 239668
rect 238342 239053 238402 292027
rect 238526 240005 238586 292571
rect 239259 291548 239325 291549
rect 239259 291484 239260 291548
rect 239324 291484 239325 291548
rect 239259 291483 239325 291484
rect 238523 240004 238589 240005
rect 238523 239940 238524 240004
rect 238588 239940 238589 240004
rect 238523 239939 238589 239940
rect 238339 239052 238405 239053
rect 238339 238988 238340 239052
rect 238404 238988 238405 239052
rect 238339 238987 238405 238988
rect 236394 237818 236426 238054
rect 236662 237818 236746 238054
rect 236982 237818 237014 238054
rect 236394 237734 237014 237818
rect 236394 237498 236426 237734
rect 236662 237498 236746 237734
rect 236982 237498 237014 237734
rect 236394 202054 237014 237498
rect 239262 232389 239322 291483
rect 244208 291454 244528 291486
rect 244208 291218 244250 291454
rect 244486 291218 244528 291454
rect 244208 291134 244528 291218
rect 239443 291004 239509 291005
rect 239443 290940 239444 291004
rect 239508 290940 239509 291004
rect 239443 290939 239509 290940
rect 239259 232388 239325 232389
rect 239259 232324 239260 232388
rect 239324 232324 239325 232388
rect 239259 232323 239325 232324
rect 236394 201818 236426 202054
rect 236662 201818 236746 202054
rect 236982 201818 237014 202054
rect 236394 201734 237014 201818
rect 236394 201498 236426 201734
rect 236662 201498 236746 201734
rect 236982 201498 237014 201734
rect 236394 166054 237014 201498
rect 239446 192541 239506 290939
rect 244208 290898 244250 291134
rect 244486 290898 244528 291134
rect 244208 290866 244528 290898
rect 274928 291454 275248 291486
rect 274928 291218 274970 291454
rect 275206 291218 275248 291454
rect 274928 291134 275248 291218
rect 274928 290898 274970 291134
rect 275206 290898 275248 291134
rect 274928 290866 275248 290898
rect 239627 290460 239693 290461
rect 239627 290396 239628 290460
rect 239692 290396 239693 290460
rect 239627 290395 239693 290396
rect 239443 192540 239509 192541
rect 239443 192476 239444 192540
rect 239508 192476 239509 192540
rect 239443 192475 239509 192476
rect 236394 165818 236426 166054
rect 236662 165818 236746 166054
rect 236982 165818 237014 166054
rect 236394 165734 237014 165818
rect 236394 165498 236426 165734
rect 236662 165498 236746 165734
rect 236982 165498 237014 165734
rect 235211 136780 235277 136781
rect 235211 136716 235212 136780
rect 235276 136716 235277 136780
rect 235211 136715 235277 136716
rect 232674 126098 232706 126334
rect 232942 126098 233026 126334
rect 233262 126098 233294 126334
rect 232674 126014 233294 126098
rect 232674 125778 232706 126014
rect 232942 125778 233026 126014
rect 233262 125778 233294 126014
rect 232674 90334 233294 125778
rect 232674 90098 232706 90334
rect 232942 90098 233026 90334
rect 233262 90098 233294 90334
rect 232674 90014 233294 90098
rect 232674 89778 232706 90014
rect 232942 89778 233026 90014
rect 233262 89778 233294 90014
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 230979 86324 231045 86325
rect 230979 86260 230980 86324
rect 231044 86260 231045 86324
rect 230979 86259 231045 86260
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 228954 -3226 229574 14058
rect 228954 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 229574 -3226
rect 228954 -3546 229574 -3462
rect 228954 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 229574 -3546
rect 228954 -7654 229574 -3782
rect 232674 54334 233294 89778
rect 232674 54098 232706 54334
rect 232942 54098 233026 54334
rect 233262 54098 233294 54334
rect 232674 54014 233294 54098
rect 232674 53778 232706 54014
rect 232942 53778 233026 54014
rect 233262 53778 233294 54014
rect 232674 18334 233294 53778
rect 232674 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 233294 18334
rect 232674 18014 233294 18098
rect 232674 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 233294 18014
rect 232674 -4186 233294 17778
rect 232674 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 233294 -4186
rect 232674 -4506 233294 -4422
rect 232674 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 233294 -4506
rect 232674 -7654 233294 -4742
rect 236394 130054 237014 165498
rect 239630 152693 239690 290395
rect 239811 289916 239877 289917
rect 239811 289852 239812 289916
rect 239876 289852 239877 289916
rect 239811 289851 239877 289852
rect 239627 152692 239693 152693
rect 239627 152628 239628 152692
rect 239692 152628 239693 152692
rect 239627 152627 239693 152628
rect 236394 129818 236426 130054
rect 236662 129818 236746 130054
rect 236982 129818 237014 130054
rect 236394 129734 237014 129818
rect 236394 129498 236426 129734
rect 236662 129498 236746 129734
rect 236982 129498 237014 129734
rect 236394 94054 237014 129498
rect 239814 112845 239874 289851
rect 259568 259174 259888 259206
rect 259568 258938 259610 259174
rect 259846 258938 259888 259174
rect 259568 258854 259888 258938
rect 259568 258618 259610 258854
rect 259846 258618 259888 258854
rect 259568 258586 259888 258618
rect 244208 255454 244528 255486
rect 244208 255218 244250 255454
rect 244486 255218 244528 255454
rect 244208 255134 244528 255218
rect 244208 254898 244250 255134
rect 244486 254898 244528 255134
rect 244208 254866 244528 254898
rect 274928 255454 275248 255486
rect 274928 255218 274970 255454
rect 275206 255218 275248 255454
rect 274928 255134 275248 255218
rect 274928 254898 274970 255134
rect 275206 254898 275248 255134
rect 274928 254866 275248 254898
rect 240114 205774 240734 241295
rect 240114 205538 240146 205774
rect 240382 205538 240466 205774
rect 240702 205538 240734 205774
rect 240114 205454 240734 205538
rect 240114 205218 240146 205454
rect 240382 205218 240466 205454
rect 240702 205218 240734 205454
rect 240114 169774 240734 205218
rect 240114 169538 240146 169774
rect 240382 169538 240466 169774
rect 240702 169538 240734 169774
rect 240114 169454 240734 169538
rect 240114 169218 240146 169454
rect 240382 169218 240466 169454
rect 240702 169218 240734 169454
rect 240114 133774 240734 169218
rect 240114 133538 240146 133774
rect 240382 133538 240466 133774
rect 240702 133538 240734 133774
rect 240114 133454 240734 133538
rect 240114 133218 240146 133454
rect 240382 133218 240466 133454
rect 240702 133218 240734 133454
rect 239811 112844 239877 112845
rect 239811 112780 239812 112844
rect 239876 112780 239877 112844
rect 239811 112779 239877 112780
rect 236394 93818 236426 94054
rect 236662 93818 236746 94054
rect 236982 93818 237014 94054
rect 236394 93734 237014 93818
rect 236394 93498 236426 93734
rect 236662 93498 236746 93734
rect 236982 93498 237014 93734
rect 236394 58054 237014 93498
rect 236394 57818 236426 58054
rect 236662 57818 236746 58054
rect 236982 57818 237014 58054
rect 236394 57734 237014 57818
rect 236394 57498 236426 57734
rect 236662 57498 236746 57734
rect 236982 57498 237014 57734
rect 236394 22054 237014 57498
rect 236394 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 237014 22054
rect 236394 21734 237014 21818
rect 236394 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 237014 21734
rect 236394 -5146 237014 21498
rect 236394 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 237014 -5146
rect 236394 -5466 237014 -5382
rect 236394 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 237014 -5466
rect 236394 -7654 237014 -5702
rect 240114 97774 240734 133218
rect 240114 97538 240146 97774
rect 240382 97538 240466 97774
rect 240702 97538 240734 97774
rect 240114 97454 240734 97538
rect 240114 97218 240146 97454
rect 240382 97218 240466 97454
rect 240702 97218 240734 97454
rect 240114 61774 240734 97218
rect 240114 61538 240146 61774
rect 240382 61538 240466 61774
rect 240702 61538 240734 61774
rect 240114 61454 240734 61538
rect 240114 61218 240146 61454
rect 240382 61218 240466 61454
rect 240702 61218 240734 61454
rect 240114 25774 240734 61218
rect 240114 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 240734 25774
rect 240114 25454 240734 25538
rect 240114 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 240734 25454
rect 240114 -6106 240734 25218
rect 240114 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 240734 -6106
rect 240114 -6426 240734 -6342
rect 240114 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 240734 -6426
rect 240114 -7654 240734 -6662
rect 243834 209494 244454 239988
rect 243834 209258 243866 209494
rect 244102 209258 244186 209494
rect 244422 209258 244454 209494
rect 243834 209174 244454 209258
rect 243834 208938 243866 209174
rect 244102 208938 244186 209174
rect 244422 208938 244454 209174
rect 243834 173494 244454 208938
rect 243834 173258 243866 173494
rect 244102 173258 244186 173494
rect 244422 173258 244454 173494
rect 243834 173174 244454 173258
rect 243834 172938 243866 173174
rect 244102 172938 244186 173174
rect 244422 172938 244454 173174
rect 243834 137494 244454 172938
rect 243834 137258 243866 137494
rect 244102 137258 244186 137494
rect 244422 137258 244454 137494
rect 243834 137174 244454 137258
rect 243834 136938 243866 137174
rect 244102 136938 244186 137174
rect 244422 136938 244454 137174
rect 243834 101494 244454 136938
rect 243834 101258 243866 101494
rect 244102 101258 244186 101494
rect 244422 101258 244454 101494
rect 243834 101174 244454 101258
rect 243834 100938 243866 101174
rect 244102 100938 244186 101174
rect 244422 100938 244454 101174
rect 243834 65494 244454 100938
rect 243834 65258 243866 65494
rect 244102 65258 244186 65494
rect 244422 65258 244454 65494
rect 243834 65174 244454 65258
rect 243834 64938 243866 65174
rect 244102 64938 244186 65174
rect 244422 64938 244454 65174
rect 243834 29494 244454 64938
rect 243834 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 244454 29494
rect 243834 29174 244454 29258
rect 243834 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 244454 29174
rect 243834 -7066 244454 28938
rect 243834 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 244454 -7066
rect 243834 -7386 244454 -7302
rect 243834 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 244454 -7386
rect 243834 -7654 244454 -7622
rect 253794 219454 254414 241295
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 257514 223174 258134 241295
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -1306 258134 6618
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -7654 258134 -1862
rect 261234 226894 261854 241295
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -2266 261854 10338
rect 261234 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 261854 -2266
rect 261234 -2586 261854 -2502
rect 261234 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 261854 -2586
rect 261234 -7654 261854 -2822
rect 264954 230614 265574 241295
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 264954 -3226 265574 14058
rect 264954 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 265574 -3226
rect 264954 -3546 265574 -3462
rect 264954 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 265574 -3546
rect 264954 -7654 265574 -3782
rect 268674 234334 269294 241295
rect 268674 234098 268706 234334
rect 268942 234098 269026 234334
rect 269262 234098 269294 234334
rect 268674 234014 269294 234098
rect 268674 233778 268706 234014
rect 268942 233778 269026 234014
rect 269262 233778 269294 234014
rect 268674 198334 269294 233778
rect 268674 198098 268706 198334
rect 268942 198098 269026 198334
rect 269262 198098 269294 198334
rect 268674 198014 269294 198098
rect 268674 197778 268706 198014
rect 268942 197778 269026 198014
rect 269262 197778 269294 198014
rect 268674 162334 269294 197778
rect 268674 162098 268706 162334
rect 268942 162098 269026 162334
rect 269262 162098 269294 162334
rect 268674 162014 269294 162098
rect 268674 161778 268706 162014
rect 268942 161778 269026 162014
rect 269262 161778 269294 162014
rect 268674 126334 269294 161778
rect 268674 126098 268706 126334
rect 268942 126098 269026 126334
rect 269262 126098 269294 126334
rect 268674 126014 269294 126098
rect 268674 125778 268706 126014
rect 268942 125778 269026 126014
rect 269262 125778 269294 126014
rect 268674 90334 269294 125778
rect 268674 90098 268706 90334
rect 268942 90098 269026 90334
rect 269262 90098 269294 90334
rect 268674 90014 269294 90098
rect 268674 89778 268706 90014
rect 268942 89778 269026 90014
rect 269262 89778 269294 90014
rect 268674 54334 269294 89778
rect 268674 54098 268706 54334
rect 268942 54098 269026 54334
rect 269262 54098 269294 54334
rect 268674 54014 269294 54098
rect 268674 53778 268706 54014
rect 268942 53778 269026 54014
rect 269262 53778 269294 54014
rect 268674 18334 269294 53778
rect 268674 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 269294 18334
rect 268674 18014 269294 18098
rect 268674 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 269294 18014
rect 268674 -4186 269294 17778
rect 268674 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 269294 -4186
rect 268674 -4506 269294 -4422
rect 268674 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 269294 -4506
rect 268674 -7654 269294 -4742
rect 272394 238054 273014 241295
rect 272394 237818 272426 238054
rect 272662 237818 272746 238054
rect 272982 237818 273014 238054
rect 272394 237734 273014 237818
rect 272394 237498 272426 237734
rect 272662 237498 272746 237734
rect 272982 237498 273014 237734
rect 272394 202054 273014 237498
rect 272394 201818 272426 202054
rect 272662 201818 272746 202054
rect 272982 201818 273014 202054
rect 272394 201734 273014 201818
rect 272394 201498 272426 201734
rect 272662 201498 272746 201734
rect 272982 201498 273014 201734
rect 272394 166054 273014 201498
rect 272394 165818 272426 166054
rect 272662 165818 272746 166054
rect 272982 165818 273014 166054
rect 272394 165734 273014 165818
rect 272394 165498 272426 165734
rect 272662 165498 272746 165734
rect 272982 165498 273014 165734
rect 272394 130054 273014 165498
rect 272394 129818 272426 130054
rect 272662 129818 272746 130054
rect 272982 129818 273014 130054
rect 272394 129734 273014 129818
rect 272394 129498 272426 129734
rect 272662 129498 272746 129734
rect 272982 129498 273014 129734
rect 272394 94054 273014 129498
rect 272394 93818 272426 94054
rect 272662 93818 272746 94054
rect 272982 93818 273014 94054
rect 272394 93734 273014 93818
rect 272394 93498 272426 93734
rect 272662 93498 272746 93734
rect 272982 93498 273014 93734
rect 272394 58054 273014 93498
rect 272394 57818 272426 58054
rect 272662 57818 272746 58054
rect 272982 57818 273014 58054
rect 272394 57734 273014 57818
rect 272394 57498 272426 57734
rect 272662 57498 272746 57734
rect 272982 57498 273014 57734
rect 272394 22054 273014 57498
rect 272394 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 273014 22054
rect 272394 21734 273014 21818
rect 272394 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 273014 21734
rect 272394 -5146 273014 21498
rect 272394 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 273014 -5146
rect 272394 -5466 273014 -5382
rect 272394 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 273014 -5466
rect 272394 -7654 273014 -5702
rect 276114 205774 276734 241295
rect 279374 228309 279434 303723
rect 279834 281494 280454 316938
rect 280659 314668 280725 314669
rect 280659 314604 280660 314668
rect 280724 314604 280725 314668
rect 280659 314603 280725 314604
rect 279834 281258 279866 281494
rect 280102 281258 280186 281494
rect 280422 281258 280454 281494
rect 279834 281174 280454 281258
rect 279834 280938 279866 281174
rect 280102 280938 280186 281174
rect 280422 280938 280454 281174
rect 279834 245494 280454 280938
rect 279834 245258 279866 245494
rect 280102 245258 280186 245494
rect 280422 245258 280454 245494
rect 279834 245174 280454 245258
rect 279834 244938 279866 245174
rect 280102 244938 280186 245174
rect 280422 244938 280454 245174
rect 279555 241908 279621 241909
rect 279555 241844 279556 241908
rect 279620 241844 279621 241908
rect 279555 241843 279621 241844
rect 279371 228308 279437 228309
rect 279371 228244 279372 228308
rect 279436 228244 279437 228308
rect 279371 228243 279437 228244
rect 279558 225589 279618 241843
rect 279555 225588 279621 225589
rect 279555 225524 279556 225588
rect 279620 225524 279621 225588
rect 279555 225523 279621 225524
rect 276114 205538 276146 205774
rect 276382 205538 276466 205774
rect 276702 205538 276734 205774
rect 276114 205454 276734 205538
rect 276114 205218 276146 205454
rect 276382 205218 276466 205454
rect 276702 205218 276734 205454
rect 276114 169774 276734 205218
rect 276114 169538 276146 169774
rect 276382 169538 276466 169774
rect 276702 169538 276734 169774
rect 276114 169454 276734 169538
rect 276114 169218 276146 169454
rect 276382 169218 276466 169454
rect 276702 169218 276734 169454
rect 276114 133774 276734 169218
rect 276114 133538 276146 133774
rect 276382 133538 276466 133774
rect 276702 133538 276734 133774
rect 276114 133454 276734 133538
rect 276114 133218 276146 133454
rect 276382 133218 276466 133454
rect 276702 133218 276734 133454
rect 276114 97774 276734 133218
rect 276114 97538 276146 97774
rect 276382 97538 276466 97774
rect 276702 97538 276734 97774
rect 276114 97454 276734 97538
rect 276114 97218 276146 97454
rect 276382 97218 276466 97454
rect 276702 97218 276734 97454
rect 276114 61774 276734 97218
rect 276114 61538 276146 61774
rect 276382 61538 276466 61774
rect 276702 61538 276734 61774
rect 276114 61454 276734 61538
rect 276114 61218 276146 61454
rect 276382 61218 276466 61454
rect 276702 61218 276734 61454
rect 276114 25774 276734 61218
rect 276114 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 276734 25774
rect 276114 25454 276734 25538
rect 276114 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 276734 25454
rect 276114 -6106 276734 25218
rect 276114 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 276734 -6106
rect 276114 -6426 276734 -6342
rect 276114 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 276734 -6426
rect 276114 -7654 276734 -6662
rect 279834 209494 280454 244938
rect 279834 209258 279866 209494
rect 280102 209258 280186 209494
rect 280422 209258 280454 209494
rect 279834 209174 280454 209258
rect 279834 208938 279866 209174
rect 280102 208938 280186 209174
rect 280422 208938 280454 209174
rect 279834 173494 280454 208938
rect 279834 173258 279866 173494
rect 280102 173258 280186 173494
rect 280422 173258 280454 173494
rect 279834 173174 280454 173258
rect 279834 172938 279866 173174
rect 280102 172938 280186 173174
rect 280422 172938 280454 173174
rect 279834 137494 280454 172938
rect 279834 137258 279866 137494
rect 280102 137258 280186 137494
rect 280422 137258 280454 137494
rect 279834 137174 280454 137258
rect 279834 136938 279866 137174
rect 280102 136938 280186 137174
rect 280422 136938 280454 137174
rect 279834 101494 280454 136938
rect 279834 101258 279866 101494
rect 280102 101258 280186 101494
rect 280422 101258 280454 101494
rect 279834 101174 280454 101258
rect 279834 100938 279866 101174
rect 280102 100938 280186 101174
rect 280422 100938 280454 101174
rect 279834 65494 280454 100938
rect 279834 65258 279866 65494
rect 280102 65258 280186 65494
rect 280422 65258 280454 65494
rect 279834 65174 280454 65258
rect 279834 64938 279866 65174
rect 280102 64938 280186 65174
rect 280422 64938 280454 65174
rect 279834 29494 280454 64938
rect 280662 32605 280722 314603
rect 280846 220285 280906 339083
rect 281763 302428 281829 302429
rect 281763 302364 281764 302428
rect 281828 302364 281829 302428
rect 281763 302363 281829 302364
rect 281579 292908 281645 292909
rect 281579 292844 281580 292908
rect 281644 292844 281645 292908
rect 281579 292843 281645 292844
rect 281027 291548 281093 291549
rect 281027 291484 281028 291548
rect 281092 291484 281093 291548
rect 281027 291483 281093 291484
rect 280843 220284 280909 220285
rect 280843 220220 280844 220284
rect 280908 220220 280909 220284
rect 280843 220219 280909 220220
rect 281030 202197 281090 291483
rect 281582 218653 281642 292843
rect 281766 233885 281826 302363
rect 282131 299708 282197 299709
rect 282131 299644 282132 299708
rect 282196 299644 282197 299708
rect 282131 299643 282197 299644
rect 282134 274685 282194 299643
rect 282870 276589 282930 467331
rect 287099 462636 287165 462637
rect 287099 462572 287100 462636
rect 287164 462572 287165 462636
rect 287099 462571 287165 462572
rect 285627 318748 285693 318749
rect 285627 318684 285628 318748
rect 285692 318684 285693 318748
rect 285627 318683 285693 318684
rect 284339 317388 284405 317389
rect 284339 317324 284340 317388
rect 284404 317324 284405 317388
rect 284339 317323 284405 317324
rect 283051 290188 283117 290189
rect 283051 290124 283052 290188
rect 283116 290124 283117 290188
rect 283051 290123 283117 290124
rect 282867 276588 282933 276589
rect 282867 276524 282868 276588
rect 282932 276524 282933 276588
rect 282867 276523 282933 276524
rect 282131 274684 282197 274685
rect 282131 274620 282132 274684
rect 282196 274620 282197 274684
rect 282131 274619 282197 274620
rect 281763 233884 281829 233885
rect 281763 233820 281764 233884
rect 281828 233820 281829 233884
rect 281763 233819 281829 233820
rect 281579 218652 281645 218653
rect 281579 218588 281580 218652
rect 281644 218588 281645 218652
rect 281579 218587 281645 218588
rect 283054 217293 283114 290123
rect 283419 286108 283485 286109
rect 283419 286044 283420 286108
rect 283484 286044 283485 286108
rect 283419 286043 283485 286044
rect 283235 284748 283301 284749
rect 283235 284684 283236 284748
rect 283300 284684 283301 284748
rect 283235 284683 283301 284684
rect 283238 240685 283298 284683
rect 283235 240684 283301 240685
rect 283235 240620 283236 240684
rect 283300 240620 283301 240684
rect 283235 240619 283301 240620
rect 283051 217292 283117 217293
rect 283051 217228 283052 217292
rect 283116 217228 283117 217292
rect 283051 217227 283117 217228
rect 283422 215933 283482 286043
rect 283419 215932 283485 215933
rect 283419 215868 283420 215932
rect 283484 215868 283485 215932
rect 283419 215867 283485 215868
rect 281027 202196 281093 202197
rect 281027 202132 281028 202196
rect 281092 202132 281093 202196
rect 281027 202131 281093 202132
rect 280659 32604 280725 32605
rect 280659 32540 280660 32604
rect 280724 32540 280725 32604
rect 280659 32539 280725 32540
rect 279834 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 280454 29494
rect 279834 29174 280454 29258
rect 279834 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 280454 29174
rect 279834 -7066 280454 28938
rect 284342 7717 284402 317323
rect 284523 307868 284589 307869
rect 284523 307804 284524 307868
rect 284588 307804 284589 307868
rect 284523 307803 284589 307804
rect 284526 27029 284586 307803
rect 284707 301068 284773 301069
rect 284707 301004 284708 301068
rect 284772 301004 284773 301068
rect 284707 301003 284773 301004
rect 284710 240141 284770 301003
rect 284891 294268 284957 294269
rect 284891 294204 284892 294268
rect 284956 294204 284957 294268
rect 284891 294203 284957 294204
rect 284707 240140 284773 240141
rect 284707 240076 284708 240140
rect 284772 240076 284773 240140
rect 284707 240075 284773 240076
rect 284894 235381 284954 294203
rect 284891 235380 284957 235381
rect 284891 235316 284892 235380
rect 284956 235316 284957 235380
rect 284891 235315 284957 235316
rect 285630 29749 285690 318683
rect 287102 281893 287162 462571
rect 287283 444004 287349 444005
rect 287283 443940 287284 444004
rect 287348 443940 287349 444004
rect 287283 443939 287349 443940
rect 287286 282981 287346 443939
rect 289794 435454 290414 470898
rect 291150 456245 291210 626315
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 291699 618220 291765 618221
rect 291699 618156 291700 618220
rect 291764 618156 291765 618220
rect 291699 618155 291765 618156
rect 291515 614140 291581 614141
rect 291515 614076 291516 614140
rect 291580 614076 291581 614140
rect 291515 614075 291581 614076
rect 291331 610060 291397 610061
rect 291331 609996 291332 610060
rect 291396 609996 291397 610060
rect 291331 609995 291397 609996
rect 291334 468757 291394 609995
rect 291518 478005 291578 614075
rect 291702 481133 291762 618155
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 291699 481132 291765 481133
rect 291699 481068 291700 481132
rect 291764 481068 291765 481132
rect 291699 481067 291765 481068
rect 291515 478004 291581 478005
rect 291515 477940 291516 478004
rect 291580 477940 291581 478004
rect 291515 477939 291581 477940
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 291331 468756 291397 468757
rect 291331 468692 291332 468756
rect 291396 468692 291397 468756
rect 291331 468691 291397 468692
rect 291147 456244 291213 456245
rect 291147 456180 291148 456244
rect 291212 456180 291213 456244
rect 291147 456179 291213 456180
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 287467 392188 287533 392189
rect 287467 392124 287468 392188
rect 287532 392124 287533 392188
rect 287467 392123 287533 392124
rect 287283 282980 287349 282981
rect 287283 282916 287284 282980
rect 287348 282916 287349 282980
rect 287283 282915 287349 282916
rect 287283 282028 287349 282029
rect 287283 281964 287284 282028
rect 287348 281964 287349 282028
rect 287283 281963 287349 281964
rect 287099 281892 287165 281893
rect 287099 281828 287100 281892
rect 287164 281828 287165 281892
rect 287099 281827 287165 281828
rect 287099 241500 287165 241501
rect 287099 241436 287100 241500
rect 287164 241436 287165 241500
rect 287099 241435 287165 241436
rect 287102 97613 287162 241435
rect 287286 240549 287346 281963
rect 287283 240548 287349 240549
rect 287283 240484 287284 240548
rect 287348 240484 287349 240548
rect 287283 240483 287349 240484
rect 287470 239733 287530 392123
rect 287651 390828 287717 390829
rect 287651 390764 287652 390828
rect 287716 390764 287717 390828
rect 287651 390763 287717 390764
rect 287654 240957 287714 390763
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 288387 287468 288453 287469
rect 288387 287404 288388 287468
rect 288452 287404 288453 287468
rect 288387 287403 288453 287404
rect 287835 283388 287901 283389
rect 287835 283324 287836 283388
rect 287900 283324 287901 283388
rect 287835 283323 287901 283324
rect 287651 240956 287717 240957
rect 287651 240892 287652 240956
rect 287716 240892 287717 240956
rect 287651 240891 287717 240892
rect 287838 239869 287898 283323
rect 287835 239868 287901 239869
rect 287835 239804 287836 239868
rect 287900 239804 287901 239868
rect 287835 239803 287901 239804
rect 287467 239732 287533 239733
rect 287467 239668 287468 239732
rect 287532 239668 287533 239732
rect 287467 239667 287533 239668
rect 288390 149837 288450 287403
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 288387 149836 288453 149837
rect 288387 149772 288388 149836
rect 288452 149772 288453 149836
rect 288387 149771 288453 149772
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 287099 97612 287165 97613
rect 287099 97548 287100 97612
rect 287164 97548 287165 97612
rect 287099 97547 287165 97548
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 285627 29748 285693 29749
rect 285627 29684 285628 29748
rect 285692 29684 285693 29748
rect 285627 29683 285693 29684
rect 284523 27028 284589 27029
rect 284523 26964 284524 27028
rect 284588 26964 284589 27028
rect 284523 26963 284589 26964
rect 284339 7716 284405 7717
rect 284339 7652 284340 7716
rect 284404 7652 284405 7716
rect 284339 7651 284405 7652
rect 279834 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 280454 -7066
rect 279834 -7386 280454 -7302
rect 279834 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 280454 -7386
rect 279834 -7654 280454 -7622
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -7654 294134 -1862
rect 297234 706758 297854 711590
rect 297234 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 297854 706758
rect 297234 706438 297854 706522
rect 297234 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 297854 706438
rect 297234 694894 297854 706202
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 300954 707718 301574 711590
rect 300954 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 301574 707718
rect 300954 707398 301574 707482
rect 300954 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 301574 707398
rect 300954 698614 301574 707162
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 299979 329084 300045 329085
rect 299979 329020 299980 329084
rect 300044 329020 300045 329084
rect 299979 329019 300045 329020
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 299982 252109 300042 329019
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 299979 252108 300045 252109
rect 299979 252044 299980 252108
rect 300044 252044 300045 252108
rect 299979 252043 300045 252044
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -2266 297854 10338
rect 297234 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 297854 -2266
rect 297234 -2586 297854 -2502
rect 297234 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 297854 -2586
rect 297234 -7654 297854 -2822
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 300954 -3226 301574 14058
rect 300954 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 301574 -3226
rect 300954 -3546 301574 -3462
rect 300954 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 301574 -3546
rect 300954 -7654 301574 -3782
rect 304674 708678 305294 711590
rect 304674 708442 304706 708678
rect 304942 708442 305026 708678
rect 305262 708442 305294 708678
rect 304674 708358 305294 708442
rect 304674 708122 304706 708358
rect 304942 708122 305026 708358
rect 305262 708122 305294 708358
rect 304674 666334 305294 708122
rect 304674 666098 304706 666334
rect 304942 666098 305026 666334
rect 305262 666098 305294 666334
rect 304674 666014 305294 666098
rect 304674 665778 304706 666014
rect 304942 665778 305026 666014
rect 305262 665778 305294 666014
rect 304674 630334 305294 665778
rect 304674 630098 304706 630334
rect 304942 630098 305026 630334
rect 305262 630098 305294 630334
rect 304674 630014 305294 630098
rect 304674 629778 304706 630014
rect 304942 629778 305026 630014
rect 305262 629778 305294 630014
rect 304674 594334 305294 629778
rect 304674 594098 304706 594334
rect 304942 594098 305026 594334
rect 305262 594098 305294 594334
rect 304674 594014 305294 594098
rect 304674 593778 304706 594014
rect 304942 593778 305026 594014
rect 305262 593778 305294 594014
rect 304674 558334 305294 593778
rect 308394 709638 309014 711590
rect 308394 709402 308426 709638
rect 308662 709402 308746 709638
rect 308982 709402 309014 709638
rect 308394 709318 309014 709402
rect 308394 709082 308426 709318
rect 308662 709082 308746 709318
rect 308982 709082 309014 709318
rect 308394 670054 309014 709082
rect 308394 669818 308426 670054
rect 308662 669818 308746 670054
rect 308982 669818 309014 670054
rect 308394 669734 309014 669818
rect 308394 669498 308426 669734
rect 308662 669498 308746 669734
rect 308982 669498 309014 669734
rect 308394 634054 309014 669498
rect 308394 633818 308426 634054
rect 308662 633818 308746 634054
rect 308982 633818 309014 634054
rect 308394 633734 309014 633818
rect 308394 633498 308426 633734
rect 308662 633498 308746 633734
rect 308982 633498 309014 633734
rect 308394 598054 309014 633498
rect 308394 597818 308426 598054
rect 308662 597818 308746 598054
rect 308982 597818 309014 598054
rect 308394 597734 309014 597818
rect 308394 597498 308426 597734
rect 308662 597498 308746 597734
rect 308982 597498 309014 597734
rect 306971 591292 307037 591293
rect 306971 591228 306972 591292
rect 307036 591228 307037 591292
rect 306971 591227 307037 591228
rect 304674 558098 304706 558334
rect 304942 558098 305026 558334
rect 305262 558098 305294 558334
rect 304674 558014 305294 558098
rect 304674 557778 304706 558014
rect 304942 557778 305026 558014
rect 305262 557778 305294 558014
rect 304674 522334 305294 557778
rect 304674 522098 304706 522334
rect 304942 522098 305026 522334
rect 305262 522098 305294 522334
rect 304674 522014 305294 522098
rect 304674 521778 304706 522014
rect 304942 521778 305026 522014
rect 305262 521778 305294 522014
rect 304674 486334 305294 521778
rect 304674 486098 304706 486334
rect 304942 486098 305026 486334
rect 305262 486098 305294 486334
rect 304674 486014 305294 486098
rect 304674 485778 304706 486014
rect 304942 485778 305026 486014
rect 305262 485778 305294 486014
rect 304674 450334 305294 485778
rect 304674 450098 304706 450334
rect 304942 450098 305026 450334
rect 305262 450098 305294 450334
rect 304674 450014 305294 450098
rect 304674 449778 304706 450014
rect 304942 449778 305026 450014
rect 305262 449778 305294 450014
rect 304674 414334 305294 449778
rect 304674 414098 304706 414334
rect 304942 414098 305026 414334
rect 305262 414098 305294 414334
rect 304674 414014 305294 414098
rect 304674 413778 304706 414014
rect 304942 413778 305026 414014
rect 305262 413778 305294 414014
rect 304674 378334 305294 413778
rect 304674 378098 304706 378334
rect 304942 378098 305026 378334
rect 305262 378098 305294 378334
rect 304674 378014 305294 378098
rect 304674 377778 304706 378014
rect 304942 377778 305026 378014
rect 305262 377778 305294 378014
rect 304674 342334 305294 377778
rect 304674 342098 304706 342334
rect 304942 342098 305026 342334
rect 305262 342098 305294 342334
rect 304674 342014 305294 342098
rect 304674 341778 304706 342014
rect 304942 341778 305026 342014
rect 305262 341778 305294 342014
rect 304674 306334 305294 341778
rect 304674 306098 304706 306334
rect 304942 306098 305026 306334
rect 305262 306098 305294 306334
rect 304674 306014 305294 306098
rect 304674 305778 304706 306014
rect 304942 305778 305026 306014
rect 305262 305778 305294 306014
rect 304674 270334 305294 305778
rect 304674 270098 304706 270334
rect 304942 270098 305026 270334
rect 305262 270098 305294 270334
rect 304674 270014 305294 270098
rect 304674 269778 304706 270014
rect 304942 269778 305026 270014
rect 305262 269778 305294 270014
rect 304674 234334 305294 269778
rect 306974 258909 307034 591227
rect 308394 562054 309014 597498
rect 308394 561818 308426 562054
rect 308662 561818 308746 562054
rect 308982 561818 309014 562054
rect 308394 561734 309014 561818
rect 308394 561498 308426 561734
rect 308662 561498 308746 561734
rect 308982 561498 309014 561734
rect 308394 526054 309014 561498
rect 308394 525818 308426 526054
rect 308662 525818 308746 526054
rect 308982 525818 309014 526054
rect 308394 525734 309014 525818
rect 308394 525498 308426 525734
rect 308662 525498 308746 525734
rect 308982 525498 309014 525734
rect 308394 490054 309014 525498
rect 312114 710598 312734 711590
rect 312114 710362 312146 710598
rect 312382 710362 312466 710598
rect 312702 710362 312734 710598
rect 312114 710278 312734 710362
rect 312114 710042 312146 710278
rect 312382 710042 312466 710278
rect 312702 710042 312734 710278
rect 312114 673774 312734 710042
rect 312114 673538 312146 673774
rect 312382 673538 312466 673774
rect 312702 673538 312734 673774
rect 312114 673454 312734 673538
rect 312114 673218 312146 673454
rect 312382 673218 312466 673454
rect 312702 673218 312734 673454
rect 312114 637774 312734 673218
rect 312114 637538 312146 637774
rect 312382 637538 312466 637774
rect 312702 637538 312734 637774
rect 312114 637454 312734 637538
rect 312114 637218 312146 637454
rect 312382 637218 312466 637454
rect 312702 637218 312734 637454
rect 312114 601774 312734 637218
rect 312114 601538 312146 601774
rect 312382 601538 312466 601774
rect 312702 601538 312734 601774
rect 312114 601454 312734 601538
rect 312114 601218 312146 601454
rect 312382 601218 312466 601454
rect 312702 601218 312734 601454
rect 312114 565774 312734 601218
rect 315834 711558 316454 711590
rect 315834 711322 315866 711558
rect 316102 711322 316186 711558
rect 316422 711322 316454 711558
rect 315834 711238 316454 711322
rect 315834 711002 315866 711238
rect 316102 711002 316186 711238
rect 316422 711002 316454 711238
rect 315834 677494 316454 711002
rect 315834 677258 315866 677494
rect 316102 677258 316186 677494
rect 316422 677258 316454 677494
rect 315834 677174 316454 677258
rect 315834 676938 315866 677174
rect 316102 676938 316186 677174
rect 316422 676938 316454 677174
rect 315834 641494 316454 676938
rect 315834 641258 315866 641494
rect 316102 641258 316186 641494
rect 316422 641258 316454 641494
rect 315834 641174 316454 641258
rect 315834 640938 315866 641174
rect 316102 640938 316186 641174
rect 316422 640938 316454 641174
rect 315834 605494 316454 640938
rect 315834 605258 315866 605494
rect 316102 605258 316186 605494
rect 316422 605258 316454 605494
rect 315834 605174 316454 605258
rect 315834 604938 315866 605174
rect 316102 604938 316186 605174
rect 316422 604938 316454 605174
rect 313779 577692 313845 577693
rect 313779 577628 313780 577692
rect 313844 577628 313845 577692
rect 313779 577627 313845 577628
rect 312114 565538 312146 565774
rect 312382 565538 312466 565774
rect 312702 565538 312734 565774
rect 312114 565454 312734 565538
rect 312114 565218 312146 565454
rect 312382 565218 312466 565454
rect 312702 565218 312734 565454
rect 312114 529774 312734 565218
rect 312114 529538 312146 529774
rect 312382 529538 312466 529774
rect 312702 529538 312734 529774
rect 312114 529454 312734 529538
rect 312114 529218 312146 529454
rect 312382 529218 312466 529454
rect 312702 529218 312734 529454
rect 309731 524516 309797 524517
rect 309731 524452 309732 524516
rect 309796 524452 309797 524516
rect 309731 524451 309797 524452
rect 308394 489818 308426 490054
rect 308662 489818 308746 490054
rect 308982 489818 309014 490054
rect 308394 489734 309014 489818
rect 308394 489498 308426 489734
rect 308662 489498 308746 489734
rect 308982 489498 309014 489734
rect 308394 454054 309014 489498
rect 308394 453818 308426 454054
rect 308662 453818 308746 454054
rect 308982 453818 309014 454054
rect 308394 453734 309014 453818
rect 308394 453498 308426 453734
rect 308662 453498 308746 453734
rect 308982 453498 309014 453734
rect 308394 418054 309014 453498
rect 308394 417818 308426 418054
rect 308662 417818 308746 418054
rect 308982 417818 309014 418054
rect 308394 417734 309014 417818
rect 308394 417498 308426 417734
rect 308662 417498 308746 417734
rect 308982 417498 309014 417734
rect 308394 382054 309014 417498
rect 308394 381818 308426 382054
rect 308662 381818 308746 382054
rect 308982 381818 309014 382054
rect 308394 381734 309014 381818
rect 308394 381498 308426 381734
rect 308662 381498 308746 381734
rect 308982 381498 309014 381734
rect 308394 346054 309014 381498
rect 308394 345818 308426 346054
rect 308662 345818 308746 346054
rect 308982 345818 309014 346054
rect 308394 345734 309014 345818
rect 308394 345498 308426 345734
rect 308662 345498 308746 345734
rect 308982 345498 309014 345734
rect 308394 310054 309014 345498
rect 308394 309818 308426 310054
rect 308662 309818 308746 310054
rect 308982 309818 309014 310054
rect 308394 309734 309014 309818
rect 308394 309498 308426 309734
rect 308662 309498 308746 309734
rect 308982 309498 309014 309734
rect 308394 274054 309014 309498
rect 308394 273818 308426 274054
rect 308662 273818 308746 274054
rect 308982 273818 309014 274054
rect 308394 273734 309014 273818
rect 308394 273498 308426 273734
rect 308662 273498 308746 273734
rect 308982 273498 309014 273734
rect 306971 258908 307037 258909
rect 306971 258844 306972 258908
rect 307036 258844 307037 258908
rect 306971 258843 307037 258844
rect 304674 234098 304706 234334
rect 304942 234098 305026 234334
rect 305262 234098 305294 234334
rect 304674 234014 305294 234098
rect 304674 233778 304706 234014
rect 304942 233778 305026 234014
rect 305262 233778 305294 234014
rect 304674 198334 305294 233778
rect 304674 198098 304706 198334
rect 304942 198098 305026 198334
rect 305262 198098 305294 198334
rect 304674 198014 305294 198098
rect 304674 197778 304706 198014
rect 304942 197778 305026 198014
rect 305262 197778 305294 198014
rect 304674 162334 305294 197778
rect 304674 162098 304706 162334
rect 304942 162098 305026 162334
rect 305262 162098 305294 162334
rect 304674 162014 305294 162098
rect 304674 161778 304706 162014
rect 304942 161778 305026 162014
rect 305262 161778 305294 162014
rect 304674 126334 305294 161778
rect 304674 126098 304706 126334
rect 304942 126098 305026 126334
rect 305262 126098 305294 126334
rect 304674 126014 305294 126098
rect 304674 125778 304706 126014
rect 304942 125778 305026 126014
rect 305262 125778 305294 126014
rect 304674 90334 305294 125778
rect 304674 90098 304706 90334
rect 304942 90098 305026 90334
rect 305262 90098 305294 90334
rect 304674 90014 305294 90098
rect 304674 89778 304706 90014
rect 304942 89778 305026 90014
rect 305262 89778 305294 90014
rect 304674 54334 305294 89778
rect 304674 54098 304706 54334
rect 304942 54098 305026 54334
rect 305262 54098 305294 54334
rect 304674 54014 305294 54098
rect 304674 53778 304706 54014
rect 304942 53778 305026 54014
rect 305262 53778 305294 54014
rect 304674 18334 305294 53778
rect 304674 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 305294 18334
rect 304674 18014 305294 18098
rect 304674 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 305294 18014
rect 304674 -4186 305294 17778
rect 304674 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 305294 -4186
rect 304674 -4506 305294 -4422
rect 304674 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 305294 -4506
rect 304674 -7654 305294 -4742
rect 308394 238054 309014 273498
rect 309734 256189 309794 524451
rect 312114 493774 312734 529218
rect 312114 493538 312146 493774
rect 312382 493538 312466 493774
rect 312702 493538 312734 493774
rect 312114 493454 312734 493538
rect 312114 493218 312146 493454
rect 312382 493218 312466 493454
rect 312702 493218 312734 493454
rect 312114 457774 312734 493218
rect 312114 457538 312146 457774
rect 312382 457538 312466 457774
rect 312702 457538 312734 457774
rect 312114 457454 312734 457538
rect 312114 457218 312146 457454
rect 312382 457218 312466 457454
rect 312702 457218 312734 457454
rect 312114 421774 312734 457218
rect 312114 421538 312146 421774
rect 312382 421538 312466 421774
rect 312702 421538 312734 421774
rect 312114 421454 312734 421538
rect 312114 421218 312146 421454
rect 312382 421218 312466 421454
rect 312702 421218 312734 421454
rect 312114 385774 312734 421218
rect 312114 385538 312146 385774
rect 312382 385538 312466 385774
rect 312702 385538 312734 385774
rect 312114 385454 312734 385538
rect 312114 385218 312146 385454
rect 312382 385218 312466 385454
rect 312702 385218 312734 385454
rect 312114 349774 312734 385218
rect 312114 349538 312146 349774
rect 312382 349538 312466 349774
rect 312702 349538 312734 349774
rect 312114 349454 312734 349538
rect 312114 349218 312146 349454
rect 312382 349218 312466 349454
rect 312702 349218 312734 349454
rect 312114 313774 312734 349218
rect 312114 313538 312146 313774
rect 312382 313538 312466 313774
rect 312702 313538 312734 313774
rect 312114 313454 312734 313538
rect 312114 313218 312146 313454
rect 312382 313218 312466 313454
rect 312702 313218 312734 313454
rect 312114 277774 312734 313218
rect 312114 277538 312146 277774
rect 312382 277538 312466 277774
rect 312702 277538 312734 277774
rect 312114 277454 312734 277538
rect 312114 277218 312146 277454
rect 312382 277218 312466 277454
rect 312702 277218 312734 277454
rect 309731 256188 309797 256189
rect 309731 256124 309732 256188
rect 309796 256124 309797 256188
rect 309731 256123 309797 256124
rect 308394 237818 308426 238054
rect 308662 237818 308746 238054
rect 308982 237818 309014 238054
rect 308394 237734 309014 237818
rect 308394 237498 308426 237734
rect 308662 237498 308746 237734
rect 308982 237498 309014 237734
rect 308394 202054 309014 237498
rect 308394 201818 308426 202054
rect 308662 201818 308746 202054
rect 308982 201818 309014 202054
rect 308394 201734 309014 201818
rect 308394 201498 308426 201734
rect 308662 201498 308746 201734
rect 308982 201498 309014 201734
rect 308394 166054 309014 201498
rect 308394 165818 308426 166054
rect 308662 165818 308746 166054
rect 308982 165818 309014 166054
rect 308394 165734 309014 165818
rect 308394 165498 308426 165734
rect 308662 165498 308746 165734
rect 308982 165498 309014 165734
rect 308394 130054 309014 165498
rect 308394 129818 308426 130054
rect 308662 129818 308746 130054
rect 308982 129818 309014 130054
rect 308394 129734 309014 129818
rect 308394 129498 308426 129734
rect 308662 129498 308746 129734
rect 308982 129498 309014 129734
rect 308394 94054 309014 129498
rect 308394 93818 308426 94054
rect 308662 93818 308746 94054
rect 308982 93818 309014 94054
rect 308394 93734 309014 93818
rect 308394 93498 308426 93734
rect 308662 93498 308746 93734
rect 308982 93498 309014 93734
rect 308394 58054 309014 93498
rect 308394 57818 308426 58054
rect 308662 57818 308746 58054
rect 308982 57818 309014 58054
rect 308394 57734 309014 57818
rect 308394 57498 308426 57734
rect 308662 57498 308746 57734
rect 308982 57498 309014 57734
rect 308394 22054 309014 57498
rect 308394 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 309014 22054
rect 308394 21734 309014 21818
rect 308394 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 309014 21734
rect 308394 -5146 309014 21498
rect 308394 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 309014 -5146
rect 308394 -5466 309014 -5382
rect 308394 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 309014 -5466
rect 308394 -7654 309014 -5702
rect 312114 241774 312734 277218
rect 313782 257549 313842 577627
rect 315834 569494 316454 604938
rect 315834 569258 315866 569494
rect 316102 569258 316186 569494
rect 316422 569258 316454 569494
rect 315834 569174 316454 569258
rect 315834 568938 315866 569174
rect 316102 568938 316186 569174
rect 316422 568938 316454 569174
rect 315834 533494 316454 568938
rect 315834 533258 315866 533494
rect 316102 533258 316186 533494
rect 316422 533258 316454 533494
rect 315834 533174 316454 533258
rect 315834 532938 315866 533174
rect 316102 532938 316186 533174
rect 316422 532938 316454 533174
rect 315834 497494 316454 532938
rect 315834 497258 315866 497494
rect 316102 497258 316186 497494
rect 316422 497258 316454 497494
rect 315834 497174 316454 497258
rect 315834 496938 315866 497174
rect 316102 496938 316186 497174
rect 316422 496938 316454 497174
rect 315834 461494 316454 496938
rect 315834 461258 315866 461494
rect 316102 461258 316186 461494
rect 316422 461258 316454 461494
rect 315834 461174 316454 461258
rect 315834 460938 315866 461174
rect 316102 460938 316186 461174
rect 316422 460938 316454 461174
rect 315834 425494 316454 460938
rect 315834 425258 315866 425494
rect 316102 425258 316186 425494
rect 316422 425258 316454 425494
rect 315834 425174 316454 425258
rect 315834 424938 315866 425174
rect 316102 424938 316186 425174
rect 316422 424938 316454 425174
rect 315834 389494 316454 424938
rect 315834 389258 315866 389494
rect 316102 389258 316186 389494
rect 316422 389258 316454 389494
rect 315834 389174 316454 389258
rect 315834 388938 315866 389174
rect 316102 388938 316186 389174
rect 316422 388938 316454 389174
rect 315834 353494 316454 388938
rect 315834 353258 315866 353494
rect 316102 353258 316186 353494
rect 316422 353258 316454 353494
rect 315834 353174 316454 353258
rect 315834 352938 315866 353174
rect 316102 352938 316186 353174
rect 316422 352938 316454 353174
rect 315834 317494 316454 352938
rect 315834 317258 315866 317494
rect 316102 317258 316186 317494
rect 316422 317258 316454 317494
rect 315834 317174 316454 317258
rect 315834 316938 315866 317174
rect 316102 316938 316186 317174
rect 316422 316938 316454 317174
rect 315834 281494 316454 316938
rect 315834 281258 315866 281494
rect 316102 281258 316186 281494
rect 316422 281258 316454 281494
rect 315834 281174 316454 281258
rect 315834 280938 315866 281174
rect 316102 280938 316186 281174
rect 316422 280938 316454 281174
rect 313779 257548 313845 257549
rect 313779 257484 313780 257548
rect 313844 257484 313845 257548
rect 313779 257483 313845 257484
rect 312114 241538 312146 241774
rect 312382 241538 312466 241774
rect 312702 241538 312734 241774
rect 312114 241454 312734 241538
rect 312114 241218 312146 241454
rect 312382 241218 312466 241454
rect 312702 241218 312734 241454
rect 312114 205774 312734 241218
rect 312114 205538 312146 205774
rect 312382 205538 312466 205774
rect 312702 205538 312734 205774
rect 312114 205454 312734 205538
rect 312114 205218 312146 205454
rect 312382 205218 312466 205454
rect 312702 205218 312734 205454
rect 312114 169774 312734 205218
rect 312114 169538 312146 169774
rect 312382 169538 312466 169774
rect 312702 169538 312734 169774
rect 312114 169454 312734 169538
rect 312114 169218 312146 169454
rect 312382 169218 312466 169454
rect 312702 169218 312734 169454
rect 312114 133774 312734 169218
rect 312114 133538 312146 133774
rect 312382 133538 312466 133774
rect 312702 133538 312734 133774
rect 312114 133454 312734 133538
rect 312114 133218 312146 133454
rect 312382 133218 312466 133454
rect 312702 133218 312734 133454
rect 312114 97774 312734 133218
rect 312114 97538 312146 97774
rect 312382 97538 312466 97774
rect 312702 97538 312734 97774
rect 312114 97454 312734 97538
rect 312114 97218 312146 97454
rect 312382 97218 312466 97454
rect 312702 97218 312734 97454
rect 312114 61774 312734 97218
rect 312114 61538 312146 61774
rect 312382 61538 312466 61774
rect 312702 61538 312734 61774
rect 312114 61454 312734 61538
rect 312114 61218 312146 61454
rect 312382 61218 312466 61454
rect 312702 61218 312734 61454
rect 312114 25774 312734 61218
rect 312114 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 312734 25774
rect 312114 25454 312734 25538
rect 312114 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 312734 25454
rect 312114 -6106 312734 25218
rect 312114 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 312734 -6106
rect 312114 -6426 312734 -6342
rect 312114 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 312734 -6426
rect 312114 -7654 312734 -6662
rect 315834 245494 316454 280938
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 320771 258908 320837 258909
rect 320771 258844 320772 258908
rect 320836 258844 320837 258908
rect 320771 258843 320837 258844
rect 320774 249389 320834 258843
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 320771 249388 320837 249389
rect 320771 249324 320772 249388
rect 320836 249324 320837 249388
rect 320771 249323 320837 249324
rect 315834 245258 315866 245494
rect 316102 245258 316186 245494
rect 316422 245258 316454 245494
rect 315834 245174 316454 245258
rect 315834 244938 315866 245174
rect 316102 244938 316186 245174
rect 316422 244938 316454 245174
rect 315834 209494 316454 244938
rect 315834 209258 315866 209494
rect 316102 209258 316186 209494
rect 316422 209258 316454 209494
rect 315834 209174 316454 209258
rect 315834 208938 315866 209174
rect 316102 208938 316186 209174
rect 316422 208938 316454 209174
rect 315834 173494 316454 208938
rect 315834 173258 315866 173494
rect 316102 173258 316186 173494
rect 316422 173258 316454 173494
rect 315834 173174 316454 173258
rect 315834 172938 315866 173174
rect 316102 172938 316186 173174
rect 316422 172938 316454 173174
rect 315834 137494 316454 172938
rect 315834 137258 315866 137494
rect 316102 137258 316186 137494
rect 316422 137258 316454 137494
rect 315834 137174 316454 137258
rect 315834 136938 315866 137174
rect 316102 136938 316186 137174
rect 316422 136938 316454 137174
rect 315834 101494 316454 136938
rect 315834 101258 315866 101494
rect 316102 101258 316186 101494
rect 316422 101258 316454 101494
rect 315834 101174 316454 101258
rect 315834 100938 315866 101174
rect 316102 100938 316186 101174
rect 316422 100938 316454 101174
rect 315834 65494 316454 100938
rect 315834 65258 315866 65494
rect 316102 65258 316186 65494
rect 316422 65258 316454 65494
rect 315834 65174 316454 65258
rect 315834 64938 315866 65174
rect 316102 64938 316186 65174
rect 316422 64938 316454 65174
rect 315834 29494 316454 64938
rect 315834 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 316454 29494
rect 315834 29174 316454 29258
rect 315834 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 316454 29174
rect 315834 -7066 316454 28938
rect 315834 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 316454 -7066
rect 315834 -7386 316454 -7302
rect 315834 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 316454 -7386
rect 315834 -7654 316454 -7622
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 329514 705798 330134 711590
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 691174 330134 705242
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -1306 330134 6618
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -7654 330134 -1862
rect 333234 706758 333854 711590
rect 333234 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 333854 706758
rect 333234 706438 333854 706522
rect 333234 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 333854 706438
rect 333234 694894 333854 706202
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -2266 333854 10338
rect 333234 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 333854 -2266
rect 333234 -2586 333854 -2502
rect 333234 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 333854 -2586
rect 333234 -7654 333854 -2822
rect 336954 707718 337574 711590
rect 336954 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 337574 707718
rect 336954 707398 337574 707482
rect 336954 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 337574 707398
rect 336954 698614 337574 707162
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 336954 -3226 337574 14058
rect 336954 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 337574 -3226
rect 336954 -3546 337574 -3462
rect 336954 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 337574 -3546
rect 336954 -7654 337574 -3782
rect 340674 708678 341294 711590
rect 340674 708442 340706 708678
rect 340942 708442 341026 708678
rect 341262 708442 341294 708678
rect 340674 708358 341294 708442
rect 340674 708122 340706 708358
rect 340942 708122 341026 708358
rect 341262 708122 341294 708358
rect 340674 666334 341294 708122
rect 340674 666098 340706 666334
rect 340942 666098 341026 666334
rect 341262 666098 341294 666334
rect 340674 666014 341294 666098
rect 340674 665778 340706 666014
rect 340942 665778 341026 666014
rect 341262 665778 341294 666014
rect 340674 630334 341294 665778
rect 340674 630098 340706 630334
rect 340942 630098 341026 630334
rect 341262 630098 341294 630334
rect 340674 630014 341294 630098
rect 340674 629778 340706 630014
rect 340942 629778 341026 630014
rect 341262 629778 341294 630014
rect 340674 594334 341294 629778
rect 340674 594098 340706 594334
rect 340942 594098 341026 594334
rect 341262 594098 341294 594334
rect 340674 594014 341294 594098
rect 340674 593778 340706 594014
rect 340942 593778 341026 594014
rect 341262 593778 341294 594014
rect 340674 558334 341294 593778
rect 340674 558098 340706 558334
rect 340942 558098 341026 558334
rect 341262 558098 341294 558334
rect 340674 558014 341294 558098
rect 340674 557778 340706 558014
rect 340942 557778 341026 558014
rect 341262 557778 341294 558014
rect 340674 522334 341294 557778
rect 340674 522098 340706 522334
rect 340942 522098 341026 522334
rect 341262 522098 341294 522334
rect 340674 522014 341294 522098
rect 340674 521778 340706 522014
rect 340942 521778 341026 522014
rect 341262 521778 341294 522014
rect 340674 486334 341294 521778
rect 340674 486098 340706 486334
rect 340942 486098 341026 486334
rect 341262 486098 341294 486334
rect 340674 486014 341294 486098
rect 340674 485778 340706 486014
rect 340942 485778 341026 486014
rect 341262 485778 341294 486014
rect 340674 450334 341294 485778
rect 340674 450098 340706 450334
rect 340942 450098 341026 450334
rect 341262 450098 341294 450334
rect 340674 450014 341294 450098
rect 340674 449778 340706 450014
rect 340942 449778 341026 450014
rect 341262 449778 341294 450014
rect 340674 414334 341294 449778
rect 340674 414098 340706 414334
rect 340942 414098 341026 414334
rect 341262 414098 341294 414334
rect 340674 414014 341294 414098
rect 340674 413778 340706 414014
rect 340942 413778 341026 414014
rect 341262 413778 341294 414014
rect 340674 378334 341294 413778
rect 340674 378098 340706 378334
rect 340942 378098 341026 378334
rect 341262 378098 341294 378334
rect 340674 378014 341294 378098
rect 340674 377778 340706 378014
rect 340942 377778 341026 378014
rect 341262 377778 341294 378014
rect 340674 342334 341294 377778
rect 340674 342098 340706 342334
rect 340942 342098 341026 342334
rect 341262 342098 341294 342334
rect 340674 342014 341294 342098
rect 340674 341778 340706 342014
rect 340942 341778 341026 342014
rect 341262 341778 341294 342014
rect 340674 306334 341294 341778
rect 340674 306098 340706 306334
rect 340942 306098 341026 306334
rect 341262 306098 341294 306334
rect 340674 306014 341294 306098
rect 340674 305778 340706 306014
rect 340942 305778 341026 306014
rect 341262 305778 341294 306014
rect 340674 270334 341294 305778
rect 340674 270098 340706 270334
rect 340942 270098 341026 270334
rect 341262 270098 341294 270334
rect 340674 270014 341294 270098
rect 340674 269778 340706 270014
rect 340942 269778 341026 270014
rect 341262 269778 341294 270014
rect 340674 234334 341294 269778
rect 340674 234098 340706 234334
rect 340942 234098 341026 234334
rect 341262 234098 341294 234334
rect 340674 234014 341294 234098
rect 340674 233778 340706 234014
rect 340942 233778 341026 234014
rect 341262 233778 341294 234014
rect 340674 198334 341294 233778
rect 340674 198098 340706 198334
rect 340942 198098 341026 198334
rect 341262 198098 341294 198334
rect 340674 198014 341294 198098
rect 340674 197778 340706 198014
rect 340942 197778 341026 198014
rect 341262 197778 341294 198014
rect 340674 162334 341294 197778
rect 340674 162098 340706 162334
rect 340942 162098 341026 162334
rect 341262 162098 341294 162334
rect 340674 162014 341294 162098
rect 340674 161778 340706 162014
rect 340942 161778 341026 162014
rect 341262 161778 341294 162014
rect 340674 126334 341294 161778
rect 340674 126098 340706 126334
rect 340942 126098 341026 126334
rect 341262 126098 341294 126334
rect 340674 126014 341294 126098
rect 340674 125778 340706 126014
rect 340942 125778 341026 126014
rect 341262 125778 341294 126014
rect 340674 90334 341294 125778
rect 340674 90098 340706 90334
rect 340942 90098 341026 90334
rect 341262 90098 341294 90334
rect 340674 90014 341294 90098
rect 340674 89778 340706 90014
rect 340942 89778 341026 90014
rect 341262 89778 341294 90014
rect 340674 54334 341294 89778
rect 340674 54098 340706 54334
rect 340942 54098 341026 54334
rect 341262 54098 341294 54334
rect 340674 54014 341294 54098
rect 340674 53778 340706 54014
rect 340942 53778 341026 54014
rect 341262 53778 341294 54014
rect 340674 18334 341294 53778
rect 340674 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 341294 18334
rect 340674 18014 341294 18098
rect 340674 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 341294 18014
rect 340674 -4186 341294 17778
rect 340674 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 341294 -4186
rect 340674 -4506 341294 -4422
rect 340674 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 341294 -4506
rect 340674 -7654 341294 -4742
rect 344394 709638 345014 711590
rect 344394 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 345014 709638
rect 344394 709318 345014 709402
rect 344394 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 345014 709318
rect 344394 670054 345014 709082
rect 344394 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 345014 670054
rect 344394 669734 345014 669818
rect 344394 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 345014 669734
rect 344394 634054 345014 669498
rect 344394 633818 344426 634054
rect 344662 633818 344746 634054
rect 344982 633818 345014 634054
rect 344394 633734 345014 633818
rect 344394 633498 344426 633734
rect 344662 633498 344746 633734
rect 344982 633498 345014 633734
rect 344394 598054 345014 633498
rect 344394 597818 344426 598054
rect 344662 597818 344746 598054
rect 344982 597818 345014 598054
rect 344394 597734 345014 597818
rect 344394 597498 344426 597734
rect 344662 597498 344746 597734
rect 344982 597498 345014 597734
rect 344394 562054 345014 597498
rect 344394 561818 344426 562054
rect 344662 561818 344746 562054
rect 344982 561818 345014 562054
rect 344394 561734 345014 561818
rect 344394 561498 344426 561734
rect 344662 561498 344746 561734
rect 344982 561498 345014 561734
rect 344394 526054 345014 561498
rect 344394 525818 344426 526054
rect 344662 525818 344746 526054
rect 344982 525818 345014 526054
rect 344394 525734 345014 525818
rect 344394 525498 344426 525734
rect 344662 525498 344746 525734
rect 344982 525498 345014 525734
rect 344394 490054 345014 525498
rect 344394 489818 344426 490054
rect 344662 489818 344746 490054
rect 344982 489818 345014 490054
rect 344394 489734 345014 489818
rect 344394 489498 344426 489734
rect 344662 489498 344746 489734
rect 344982 489498 345014 489734
rect 344394 454054 345014 489498
rect 344394 453818 344426 454054
rect 344662 453818 344746 454054
rect 344982 453818 345014 454054
rect 344394 453734 345014 453818
rect 344394 453498 344426 453734
rect 344662 453498 344746 453734
rect 344982 453498 345014 453734
rect 344394 418054 345014 453498
rect 344394 417818 344426 418054
rect 344662 417818 344746 418054
rect 344982 417818 345014 418054
rect 344394 417734 345014 417818
rect 344394 417498 344426 417734
rect 344662 417498 344746 417734
rect 344982 417498 345014 417734
rect 344394 382054 345014 417498
rect 344394 381818 344426 382054
rect 344662 381818 344746 382054
rect 344982 381818 345014 382054
rect 344394 381734 345014 381818
rect 344394 381498 344426 381734
rect 344662 381498 344746 381734
rect 344982 381498 345014 381734
rect 344394 346054 345014 381498
rect 344394 345818 344426 346054
rect 344662 345818 344746 346054
rect 344982 345818 345014 346054
rect 344394 345734 345014 345818
rect 344394 345498 344426 345734
rect 344662 345498 344746 345734
rect 344982 345498 345014 345734
rect 344394 310054 345014 345498
rect 344394 309818 344426 310054
rect 344662 309818 344746 310054
rect 344982 309818 345014 310054
rect 344394 309734 345014 309818
rect 344394 309498 344426 309734
rect 344662 309498 344746 309734
rect 344982 309498 345014 309734
rect 344394 274054 345014 309498
rect 344394 273818 344426 274054
rect 344662 273818 344746 274054
rect 344982 273818 345014 274054
rect 344394 273734 345014 273818
rect 344394 273498 344426 273734
rect 344662 273498 344746 273734
rect 344982 273498 345014 273734
rect 344394 238054 345014 273498
rect 348114 710598 348734 711590
rect 348114 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 348734 710598
rect 348114 710278 348734 710362
rect 348114 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 348734 710278
rect 348114 673774 348734 710042
rect 348114 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 348734 673774
rect 348114 673454 348734 673538
rect 348114 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 348734 673454
rect 348114 637774 348734 673218
rect 348114 637538 348146 637774
rect 348382 637538 348466 637774
rect 348702 637538 348734 637774
rect 348114 637454 348734 637538
rect 348114 637218 348146 637454
rect 348382 637218 348466 637454
rect 348702 637218 348734 637454
rect 348114 601774 348734 637218
rect 348114 601538 348146 601774
rect 348382 601538 348466 601774
rect 348702 601538 348734 601774
rect 348114 601454 348734 601538
rect 348114 601218 348146 601454
rect 348382 601218 348466 601454
rect 348702 601218 348734 601454
rect 348114 565774 348734 601218
rect 348114 565538 348146 565774
rect 348382 565538 348466 565774
rect 348702 565538 348734 565774
rect 348114 565454 348734 565538
rect 348114 565218 348146 565454
rect 348382 565218 348466 565454
rect 348702 565218 348734 565454
rect 348114 529774 348734 565218
rect 348114 529538 348146 529774
rect 348382 529538 348466 529774
rect 348702 529538 348734 529774
rect 348114 529454 348734 529538
rect 348114 529218 348146 529454
rect 348382 529218 348466 529454
rect 348702 529218 348734 529454
rect 348114 493774 348734 529218
rect 348114 493538 348146 493774
rect 348382 493538 348466 493774
rect 348702 493538 348734 493774
rect 348114 493454 348734 493538
rect 348114 493218 348146 493454
rect 348382 493218 348466 493454
rect 348702 493218 348734 493454
rect 348114 457774 348734 493218
rect 348114 457538 348146 457774
rect 348382 457538 348466 457774
rect 348702 457538 348734 457774
rect 348114 457454 348734 457538
rect 348114 457218 348146 457454
rect 348382 457218 348466 457454
rect 348702 457218 348734 457454
rect 348114 421774 348734 457218
rect 348114 421538 348146 421774
rect 348382 421538 348466 421774
rect 348702 421538 348734 421774
rect 348114 421454 348734 421538
rect 348114 421218 348146 421454
rect 348382 421218 348466 421454
rect 348702 421218 348734 421454
rect 348114 385774 348734 421218
rect 348114 385538 348146 385774
rect 348382 385538 348466 385774
rect 348702 385538 348734 385774
rect 348114 385454 348734 385538
rect 348114 385218 348146 385454
rect 348382 385218 348466 385454
rect 348702 385218 348734 385454
rect 348114 349774 348734 385218
rect 348114 349538 348146 349774
rect 348382 349538 348466 349774
rect 348702 349538 348734 349774
rect 348114 349454 348734 349538
rect 348114 349218 348146 349454
rect 348382 349218 348466 349454
rect 348702 349218 348734 349454
rect 348114 313774 348734 349218
rect 348114 313538 348146 313774
rect 348382 313538 348466 313774
rect 348702 313538 348734 313774
rect 348114 313454 348734 313538
rect 348114 313218 348146 313454
rect 348382 313218 348466 313454
rect 348702 313218 348734 313454
rect 348114 277774 348734 313218
rect 348114 277538 348146 277774
rect 348382 277538 348466 277774
rect 348702 277538 348734 277774
rect 348114 277454 348734 277538
rect 348114 277218 348146 277454
rect 348382 277218 348466 277454
rect 348702 277218 348734 277454
rect 346899 245308 346965 245309
rect 346899 245244 346900 245308
rect 346964 245244 346965 245308
rect 346899 245243 346965 245244
rect 344394 237818 344426 238054
rect 344662 237818 344746 238054
rect 344982 237818 345014 238054
rect 344394 237734 345014 237818
rect 344394 237498 344426 237734
rect 344662 237498 344746 237734
rect 344982 237498 345014 237734
rect 344394 202054 345014 237498
rect 344394 201818 344426 202054
rect 344662 201818 344746 202054
rect 344982 201818 345014 202054
rect 344394 201734 345014 201818
rect 344394 201498 344426 201734
rect 344662 201498 344746 201734
rect 344982 201498 345014 201734
rect 344394 166054 345014 201498
rect 344394 165818 344426 166054
rect 344662 165818 344746 166054
rect 344982 165818 345014 166054
rect 344394 165734 345014 165818
rect 344394 165498 344426 165734
rect 344662 165498 344746 165734
rect 344982 165498 345014 165734
rect 344394 130054 345014 165498
rect 346902 139365 346962 245243
rect 348114 241774 348734 277218
rect 348114 241538 348146 241774
rect 348382 241538 348466 241774
rect 348702 241538 348734 241774
rect 348114 241454 348734 241538
rect 348114 241218 348146 241454
rect 348382 241218 348466 241454
rect 348702 241218 348734 241454
rect 348114 205774 348734 241218
rect 348114 205538 348146 205774
rect 348382 205538 348466 205774
rect 348702 205538 348734 205774
rect 348114 205454 348734 205538
rect 348114 205218 348146 205454
rect 348382 205218 348466 205454
rect 348702 205218 348734 205454
rect 348114 169774 348734 205218
rect 348114 169538 348146 169774
rect 348382 169538 348466 169774
rect 348702 169538 348734 169774
rect 348114 169454 348734 169538
rect 348114 169218 348146 169454
rect 348382 169218 348466 169454
rect 348702 169218 348734 169454
rect 346899 139364 346965 139365
rect 346899 139300 346900 139364
rect 346964 139300 346965 139364
rect 346899 139299 346965 139300
rect 344394 129818 344426 130054
rect 344662 129818 344746 130054
rect 344982 129818 345014 130054
rect 344394 129734 345014 129818
rect 344394 129498 344426 129734
rect 344662 129498 344746 129734
rect 344982 129498 345014 129734
rect 344394 94054 345014 129498
rect 344394 93818 344426 94054
rect 344662 93818 344746 94054
rect 344982 93818 345014 94054
rect 344394 93734 345014 93818
rect 344394 93498 344426 93734
rect 344662 93498 344746 93734
rect 344982 93498 345014 93734
rect 344394 58054 345014 93498
rect 344394 57818 344426 58054
rect 344662 57818 344746 58054
rect 344982 57818 345014 58054
rect 344394 57734 345014 57818
rect 344394 57498 344426 57734
rect 344662 57498 344746 57734
rect 344982 57498 345014 57734
rect 344394 22054 345014 57498
rect 344394 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 345014 22054
rect 344394 21734 345014 21818
rect 344394 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 345014 21734
rect 344394 -5146 345014 21498
rect 344394 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 345014 -5146
rect 344394 -5466 345014 -5382
rect 344394 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 345014 -5466
rect 344394 -7654 345014 -5702
rect 348114 133774 348734 169218
rect 348114 133538 348146 133774
rect 348382 133538 348466 133774
rect 348702 133538 348734 133774
rect 348114 133454 348734 133538
rect 348114 133218 348146 133454
rect 348382 133218 348466 133454
rect 348702 133218 348734 133454
rect 348114 97774 348734 133218
rect 348114 97538 348146 97774
rect 348382 97538 348466 97774
rect 348702 97538 348734 97774
rect 348114 97454 348734 97538
rect 348114 97218 348146 97454
rect 348382 97218 348466 97454
rect 348702 97218 348734 97454
rect 348114 61774 348734 97218
rect 348114 61538 348146 61774
rect 348382 61538 348466 61774
rect 348702 61538 348734 61774
rect 348114 61454 348734 61538
rect 348114 61218 348146 61454
rect 348382 61218 348466 61454
rect 348702 61218 348734 61454
rect 348114 25774 348734 61218
rect 348114 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 348734 25774
rect 348114 25454 348734 25538
rect 348114 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 348734 25454
rect 348114 -6106 348734 25218
rect 348114 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 348734 -6106
rect 348114 -6426 348734 -6342
rect 348114 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 348734 -6426
rect 348114 -7654 348734 -6662
rect 351834 711558 352454 711590
rect 351834 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 352454 711558
rect 351834 711238 352454 711322
rect 351834 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 352454 711238
rect 351834 677494 352454 711002
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 355179 683908 355245 683909
rect 355179 683844 355180 683908
rect 355244 683844 355245 683908
rect 355179 683843 355245 683844
rect 351834 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 352454 677494
rect 351834 677174 352454 677258
rect 351834 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 352454 677174
rect 351834 641494 352454 676938
rect 351834 641258 351866 641494
rect 352102 641258 352186 641494
rect 352422 641258 352454 641494
rect 351834 641174 352454 641258
rect 351834 640938 351866 641174
rect 352102 640938 352186 641174
rect 352422 640938 352454 641174
rect 351834 605494 352454 640938
rect 351834 605258 351866 605494
rect 352102 605258 352186 605494
rect 352422 605258 352454 605494
rect 351834 605174 352454 605258
rect 351834 604938 351866 605174
rect 352102 604938 352186 605174
rect 352422 604938 352454 605174
rect 351834 569494 352454 604938
rect 351834 569258 351866 569494
rect 352102 569258 352186 569494
rect 352422 569258 352454 569494
rect 351834 569174 352454 569258
rect 351834 568938 351866 569174
rect 352102 568938 352186 569174
rect 352422 568938 352454 569174
rect 351834 533494 352454 568938
rect 351834 533258 351866 533494
rect 352102 533258 352186 533494
rect 352422 533258 352454 533494
rect 351834 533174 352454 533258
rect 351834 532938 351866 533174
rect 352102 532938 352186 533174
rect 352422 532938 352454 533174
rect 351834 497494 352454 532938
rect 351834 497258 351866 497494
rect 352102 497258 352186 497494
rect 352422 497258 352454 497494
rect 351834 497174 352454 497258
rect 351834 496938 351866 497174
rect 352102 496938 352186 497174
rect 352422 496938 352454 497174
rect 351834 461494 352454 496938
rect 351834 461258 351866 461494
rect 352102 461258 352186 461494
rect 352422 461258 352454 461494
rect 351834 461174 352454 461258
rect 351834 460938 351866 461174
rect 352102 460938 352186 461174
rect 352422 460938 352454 461174
rect 351834 425494 352454 460938
rect 351834 425258 351866 425494
rect 352102 425258 352186 425494
rect 352422 425258 352454 425494
rect 351834 425174 352454 425258
rect 351834 424938 351866 425174
rect 352102 424938 352186 425174
rect 352422 424938 352454 425174
rect 351834 389494 352454 424938
rect 351834 389258 351866 389494
rect 352102 389258 352186 389494
rect 352422 389258 352454 389494
rect 351834 389174 352454 389258
rect 351834 388938 351866 389174
rect 352102 388938 352186 389174
rect 352422 388938 352454 389174
rect 351834 353494 352454 388938
rect 351834 353258 351866 353494
rect 352102 353258 352186 353494
rect 352422 353258 352454 353494
rect 351834 353174 352454 353258
rect 351834 352938 351866 353174
rect 352102 352938 352186 353174
rect 352422 352938 352454 353174
rect 351834 317494 352454 352938
rect 351834 317258 351866 317494
rect 352102 317258 352186 317494
rect 352422 317258 352454 317494
rect 351834 317174 352454 317258
rect 351834 316938 351866 317174
rect 352102 316938 352186 317174
rect 352422 316938 352454 317174
rect 351834 281494 352454 316938
rect 351834 281258 351866 281494
rect 352102 281258 352186 281494
rect 352422 281258 352454 281494
rect 351834 281174 352454 281258
rect 351834 280938 351866 281174
rect 352102 280938 352186 281174
rect 352422 280938 352454 281174
rect 351834 245494 352454 280938
rect 355182 260269 355242 683843
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 355179 260268 355245 260269
rect 355179 260204 355180 260268
rect 355244 260204 355245 260268
rect 355179 260203 355245 260204
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 355179 248028 355245 248029
rect 355179 247964 355180 248028
rect 355244 247964 355245 248028
rect 355179 247963 355245 247964
rect 353891 246668 353957 246669
rect 353891 246604 353892 246668
rect 353956 246604 353957 246668
rect 353891 246603 353957 246604
rect 351834 245258 351866 245494
rect 352102 245258 352186 245494
rect 352422 245258 352454 245494
rect 351834 245174 352454 245258
rect 351834 244938 351866 245174
rect 352102 244938 352186 245174
rect 352422 244938 352454 245174
rect 351834 209494 352454 244938
rect 351834 209258 351866 209494
rect 352102 209258 352186 209494
rect 352422 209258 352454 209494
rect 351834 209174 352454 209258
rect 351834 208938 351866 209174
rect 352102 208938 352186 209174
rect 352422 208938 352454 209174
rect 351834 173494 352454 208938
rect 353894 179213 353954 246603
rect 355182 219061 355242 247963
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 355179 219060 355245 219061
rect 355179 218996 355180 219060
rect 355244 218996 355245 219060
rect 355179 218995 355245 218996
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 353891 179212 353957 179213
rect 353891 179148 353892 179212
rect 353956 179148 353957 179212
rect 353891 179147 353957 179148
rect 351834 173258 351866 173494
rect 352102 173258 352186 173494
rect 352422 173258 352454 173494
rect 351834 173174 352454 173258
rect 351834 172938 351866 173174
rect 352102 172938 352186 173174
rect 352422 172938 352454 173174
rect 351834 137494 352454 172938
rect 351834 137258 351866 137494
rect 352102 137258 352186 137494
rect 352422 137258 352454 137494
rect 351834 137174 352454 137258
rect 351834 136938 351866 137174
rect 352102 136938 352186 137174
rect 352422 136938 352454 137174
rect 351834 101494 352454 136938
rect 351834 101258 351866 101494
rect 352102 101258 352186 101494
rect 352422 101258 352454 101494
rect 351834 101174 352454 101258
rect 351834 100938 351866 101174
rect 352102 100938 352186 101174
rect 352422 100938 352454 101174
rect 351834 65494 352454 100938
rect 351834 65258 351866 65494
rect 352102 65258 352186 65494
rect 352422 65258 352454 65494
rect 351834 65174 352454 65258
rect 351834 64938 351866 65174
rect 352102 64938 352186 65174
rect 352422 64938 352454 65174
rect 351834 29494 352454 64938
rect 351834 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 352454 29494
rect 351834 29174 352454 29258
rect 351834 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 352454 29174
rect 351834 -7066 352454 28938
rect 351834 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 352454 -7066
rect 351834 -7386 352454 -7302
rect 351834 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 352454 -7386
rect 351834 -7654 352454 -7622
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 365514 705798 366134 711590
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 691174 366134 705242
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -1306 366134 6618
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -7654 366134 -1862
rect 369234 706758 369854 711590
rect 369234 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 369854 706758
rect 369234 706438 369854 706522
rect 369234 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 369854 706438
rect 369234 694894 369854 706202
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -2266 369854 10338
rect 369234 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 369854 -2266
rect 369234 -2586 369854 -2502
rect 369234 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 369854 -2586
rect 369234 -7654 369854 -2822
rect 372954 707718 373574 711590
rect 372954 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 373574 707718
rect 372954 707398 373574 707482
rect 372954 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 373574 707398
rect 372954 698614 373574 707162
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 372954 -3226 373574 14058
rect 372954 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 373574 -3226
rect 372954 -3546 373574 -3462
rect 372954 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 373574 -3546
rect 372954 -7654 373574 -3782
rect 376674 708678 377294 711590
rect 376674 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 377294 708678
rect 376674 708358 377294 708442
rect 376674 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 377294 708358
rect 376674 666334 377294 708122
rect 376674 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 377294 666334
rect 376674 666014 377294 666098
rect 376674 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 377294 666014
rect 376674 630334 377294 665778
rect 376674 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 377294 630334
rect 376674 630014 377294 630098
rect 376674 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 377294 630014
rect 376674 594334 377294 629778
rect 376674 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 377294 594334
rect 376674 594014 377294 594098
rect 376674 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 377294 594014
rect 376674 558334 377294 593778
rect 376674 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 377294 558334
rect 376674 558014 377294 558098
rect 376674 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 377294 558014
rect 376674 522334 377294 557778
rect 376674 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 377294 522334
rect 376674 522014 377294 522098
rect 376674 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 377294 522014
rect 376674 486334 377294 521778
rect 376674 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 377294 486334
rect 376674 486014 377294 486098
rect 376674 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 377294 486014
rect 376674 450334 377294 485778
rect 376674 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 377294 450334
rect 376674 450014 377294 450098
rect 376674 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 377294 450014
rect 376674 414334 377294 449778
rect 376674 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 377294 414334
rect 376674 414014 377294 414098
rect 376674 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 377294 414014
rect 376674 378334 377294 413778
rect 376674 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 377294 378334
rect 376674 378014 377294 378098
rect 376674 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 377294 378014
rect 376674 342334 377294 377778
rect 376674 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 377294 342334
rect 376674 342014 377294 342098
rect 376674 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 377294 342014
rect 376674 306334 377294 341778
rect 376674 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 377294 306334
rect 376674 306014 377294 306098
rect 376674 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 377294 306014
rect 376674 270334 377294 305778
rect 376674 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 377294 270334
rect 376674 270014 377294 270098
rect 376674 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 377294 270014
rect 376674 234334 377294 269778
rect 376674 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 377294 234334
rect 376674 234014 377294 234098
rect 376674 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 377294 234014
rect 376674 198334 377294 233778
rect 376674 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 377294 198334
rect 376674 198014 377294 198098
rect 376674 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 377294 198014
rect 376674 162334 377294 197778
rect 376674 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 377294 162334
rect 376674 162014 377294 162098
rect 376674 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 377294 162014
rect 376674 126334 377294 161778
rect 376674 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 377294 126334
rect 376674 126014 377294 126098
rect 376674 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 377294 126014
rect 376674 90334 377294 125778
rect 376674 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 377294 90334
rect 376674 90014 377294 90098
rect 376674 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 377294 90014
rect 376674 54334 377294 89778
rect 376674 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 377294 54334
rect 376674 54014 377294 54098
rect 376674 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 377294 54014
rect 376674 18334 377294 53778
rect 376674 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 377294 18334
rect 376674 18014 377294 18098
rect 376674 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 377294 18014
rect 376674 -4186 377294 17778
rect 376674 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 377294 -4186
rect 376674 -4506 377294 -4422
rect 376674 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 377294 -4506
rect 376674 -7654 377294 -4742
rect 380394 709638 381014 711590
rect 380394 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 381014 709638
rect 380394 709318 381014 709402
rect 380394 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 381014 709318
rect 380394 670054 381014 709082
rect 380394 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 381014 670054
rect 380394 669734 381014 669818
rect 380394 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 381014 669734
rect 380394 634054 381014 669498
rect 380394 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 381014 634054
rect 380394 633734 381014 633818
rect 380394 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 381014 633734
rect 380394 598054 381014 633498
rect 380394 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 381014 598054
rect 380394 597734 381014 597818
rect 380394 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 381014 597734
rect 380394 562054 381014 597498
rect 380394 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 381014 562054
rect 380394 561734 381014 561818
rect 380394 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 381014 561734
rect 380394 526054 381014 561498
rect 380394 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 381014 526054
rect 380394 525734 381014 525818
rect 380394 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 381014 525734
rect 380394 490054 381014 525498
rect 380394 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 381014 490054
rect 380394 489734 381014 489818
rect 380394 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 381014 489734
rect 380394 454054 381014 489498
rect 380394 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 381014 454054
rect 380394 453734 381014 453818
rect 380394 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 381014 453734
rect 380394 418054 381014 453498
rect 380394 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 381014 418054
rect 380394 417734 381014 417818
rect 380394 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 381014 417734
rect 380394 382054 381014 417498
rect 380394 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 381014 382054
rect 380394 381734 381014 381818
rect 380394 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 381014 381734
rect 380394 346054 381014 381498
rect 380394 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 381014 346054
rect 380394 345734 381014 345818
rect 380394 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 381014 345734
rect 380394 310054 381014 345498
rect 380394 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 381014 310054
rect 380394 309734 381014 309818
rect 380394 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 381014 309734
rect 380394 274054 381014 309498
rect 380394 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 381014 274054
rect 380394 273734 381014 273818
rect 380394 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 381014 273734
rect 380394 238054 381014 273498
rect 380394 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 381014 238054
rect 380394 237734 381014 237818
rect 380394 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 381014 237734
rect 380394 202054 381014 237498
rect 380394 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 381014 202054
rect 380394 201734 381014 201818
rect 380394 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 381014 201734
rect 380394 166054 381014 201498
rect 380394 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 381014 166054
rect 380394 165734 381014 165818
rect 380394 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 381014 165734
rect 380394 130054 381014 165498
rect 380394 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 381014 130054
rect 380394 129734 381014 129818
rect 380394 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 381014 129734
rect 380394 94054 381014 129498
rect 380394 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 381014 94054
rect 380394 93734 381014 93818
rect 380394 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 381014 93734
rect 380394 58054 381014 93498
rect 380394 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 381014 58054
rect 380394 57734 381014 57818
rect 380394 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 381014 57734
rect 380394 22054 381014 57498
rect 380394 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 381014 22054
rect 380394 21734 381014 21818
rect 380394 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 381014 21734
rect 380394 -5146 381014 21498
rect 380394 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 381014 -5146
rect 380394 -5466 381014 -5382
rect 380394 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 381014 -5466
rect 380394 -7654 381014 -5702
rect 384114 710598 384734 711590
rect 384114 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 384734 710598
rect 384114 710278 384734 710362
rect 384114 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 384734 710278
rect 384114 673774 384734 710042
rect 384114 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 384734 673774
rect 384114 673454 384734 673538
rect 384114 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 384734 673454
rect 384114 637774 384734 673218
rect 384114 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 384734 637774
rect 384114 637454 384734 637538
rect 384114 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 384734 637454
rect 384114 601774 384734 637218
rect 384114 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 384734 601774
rect 384114 601454 384734 601538
rect 384114 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 384734 601454
rect 384114 565774 384734 601218
rect 384114 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 384734 565774
rect 384114 565454 384734 565538
rect 384114 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 384734 565454
rect 384114 529774 384734 565218
rect 384114 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 384734 529774
rect 384114 529454 384734 529538
rect 384114 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 384734 529454
rect 384114 493774 384734 529218
rect 384114 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 384734 493774
rect 384114 493454 384734 493538
rect 384114 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 384734 493454
rect 384114 457774 384734 493218
rect 384114 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 384734 457774
rect 384114 457454 384734 457538
rect 384114 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 384734 457454
rect 384114 421774 384734 457218
rect 384114 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 384734 421774
rect 384114 421454 384734 421538
rect 384114 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 384734 421454
rect 384114 385774 384734 421218
rect 384114 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 384734 385774
rect 384114 385454 384734 385538
rect 384114 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 384734 385454
rect 384114 349774 384734 385218
rect 384114 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 384734 349774
rect 384114 349454 384734 349538
rect 384114 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 384734 349454
rect 384114 313774 384734 349218
rect 384114 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 384734 313774
rect 384114 313454 384734 313538
rect 384114 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 384734 313454
rect 384114 277774 384734 313218
rect 384114 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 384734 277774
rect 384114 277454 384734 277538
rect 384114 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 384734 277454
rect 384114 241774 384734 277218
rect 384114 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 384734 241774
rect 384114 241454 384734 241538
rect 384114 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 384734 241454
rect 384114 205774 384734 241218
rect 384114 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 384734 205774
rect 384114 205454 384734 205538
rect 384114 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 384734 205454
rect 384114 169774 384734 205218
rect 384114 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 384734 169774
rect 384114 169454 384734 169538
rect 384114 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 384734 169454
rect 384114 133774 384734 169218
rect 384114 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 384734 133774
rect 384114 133454 384734 133538
rect 384114 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 384734 133454
rect 384114 97774 384734 133218
rect 384114 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 384734 97774
rect 384114 97454 384734 97538
rect 384114 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 384734 97454
rect 384114 61774 384734 97218
rect 384114 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 384734 61774
rect 384114 61454 384734 61538
rect 384114 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 384734 61454
rect 384114 25774 384734 61218
rect 384114 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 384734 25774
rect 384114 25454 384734 25538
rect 384114 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 384734 25454
rect 384114 -6106 384734 25218
rect 384114 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 384734 -6106
rect 384114 -6426 384734 -6342
rect 384114 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 384734 -6426
rect 384114 -7654 384734 -6662
rect 387834 711558 388454 711590
rect 387834 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 388454 711558
rect 387834 711238 388454 711322
rect 387834 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 388454 711238
rect 387834 677494 388454 711002
rect 387834 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 388454 677494
rect 387834 677174 388454 677258
rect 387834 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 388454 677174
rect 387834 641494 388454 676938
rect 387834 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 388454 641494
rect 387834 641174 388454 641258
rect 387834 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 388454 641174
rect 387834 605494 388454 640938
rect 387834 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 388454 605494
rect 387834 605174 388454 605258
rect 387834 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 388454 605174
rect 387834 569494 388454 604938
rect 387834 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 388454 569494
rect 387834 569174 388454 569258
rect 387834 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 388454 569174
rect 387834 533494 388454 568938
rect 387834 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 388454 533494
rect 387834 533174 388454 533258
rect 387834 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 388454 533174
rect 387834 497494 388454 532938
rect 387834 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 388454 497494
rect 387834 497174 388454 497258
rect 387834 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 388454 497174
rect 387834 461494 388454 496938
rect 387834 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 388454 461494
rect 387834 461174 388454 461258
rect 387834 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 388454 461174
rect 387834 425494 388454 460938
rect 387834 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 388454 425494
rect 387834 425174 388454 425258
rect 387834 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 388454 425174
rect 387834 389494 388454 424938
rect 387834 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 388454 389494
rect 387834 389174 388454 389258
rect 387834 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 388454 389174
rect 387834 353494 388454 388938
rect 387834 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 388454 353494
rect 387834 353174 388454 353258
rect 387834 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 388454 353174
rect 387834 317494 388454 352938
rect 387834 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 388454 317494
rect 387834 317174 388454 317258
rect 387834 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 388454 317174
rect 387834 281494 388454 316938
rect 387834 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 388454 281494
rect 387834 281174 388454 281258
rect 387834 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 388454 281174
rect 387834 245494 388454 280938
rect 387834 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 388454 245494
rect 387834 245174 388454 245258
rect 387834 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 388454 245174
rect 387834 209494 388454 244938
rect 387834 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 388454 209494
rect 387834 209174 388454 209258
rect 387834 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 388454 209174
rect 387834 173494 388454 208938
rect 387834 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 388454 173494
rect 387834 173174 388454 173258
rect 387834 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 388454 173174
rect 387834 137494 388454 172938
rect 387834 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 388454 137494
rect 387834 137174 388454 137258
rect 387834 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 388454 137174
rect 387834 101494 388454 136938
rect 387834 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 388454 101494
rect 387834 101174 388454 101258
rect 387834 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 388454 101174
rect 387834 65494 388454 100938
rect 387834 65258 387866 65494
rect 388102 65258 388186 65494
rect 388422 65258 388454 65494
rect 387834 65174 388454 65258
rect 387834 64938 387866 65174
rect 388102 64938 388186 65174
rect 388422 64938 388454 65174
rect 387834 29494 388454 64938
rect 387834 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 388454 29494
rect 387834 29174 388454 29258
rect 387834 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 388454 29174
rect 387834 -7066 388454 28938
rect 387834 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 388454 -7066
rect 387834 -7386 388454 -7302
rect 387834 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 388454 -7386
rect 387834 -7654 388454 -7622
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 401514 705798 402134 711590
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 401514 691174 402134 705242
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -1306 402134 6618
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -7654 402134 -1862
rect 405234 706758 405854 711590
rect 405234 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 405854 706758
rect 405234 706438 405854 706522
rect 405234 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 405854 706438
rect 405234 694894 405854 706202
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -2266 405854 10338
rect 405234 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 405854 -2266
rect 405234 -2586 405854 -2502
rect 405234 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 405854 -2586
rect 405234 -7654 405854 -2822
rect 408954 707718 409574 711590
rect 408954 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 409574 707718
rect 408954 707398 409574 707482
rect 408954 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 409574 707398
rect 408954 698614 409574 707162
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 408954 -3226 409574 14058
rect 408954 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 409574 -3226
rect 408954 -3546 409574 -3462
rect 408954 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 409574 -3546
rect 408954 -7654 409574 -3782
rect 412674 708678 413294 711590
rect 412674 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 413294 708678
rect 412674 708358 413294 708442
rect 412674 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 413294 708358
rect 412674 666334 413294 708122
rect 412674 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 413294 666334
rect 412674 666014 413294 666098
rect 412674 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 413294 666014
rect 412674 630334 413294 665778
rect 412674 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 413294 630334
rect 412674 630014 413294 630098
rect 412674 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 413294 630014
rect 412674 594334 413294 629778
rect 412674 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 413294 594334
rect 412674 594014 413294 594098
rect 412674 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 413294 594014
rect 412674 558334 413294 593778
rect 412674 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 413294 558334
rect 412674 558014 413294 558098
rect 412674 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 413294 558014
rect 412674 522334 413294 557778
rect 412674 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 413294 522334
rect 412674 522014 413294 522098
rect 412674 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 413294 522014
rect 412674 486334 413294 521778
rect 412674 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 413294 486334
rect 412674 486014 413294 486098
rect 412674 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 413294 486014
rect 412674 450334 413294 485778
rect 412674 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 413294 450334
rect 412674 450014 413294 450098
rect 412674 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 413294 450014
rect 412674 414334 413294 449778
rect 412674 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 413294 414334
rect 412674 414014 413294 414098
rect 412674 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 413294 414014
rect 412674 378334 413294 413778
rect 412674 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 413294 378334
rect 412674 378014 413294 378098
rect 412674 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 413294 378014
rect 412674 342334 413294 377778
rect 412674 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 413294 342334
rect 412674 342014 413294 342098
rect 412674 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 413294 342014
rect 412674 306334 413294 341778
rect 412674 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 413294 306334
rect 412674 306014 413294 306098
rect 412674 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 413294 306014
rect 412674 270334 413294 305778
rect 412674 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 413294 270334
rect 412674 270014 413294 270098
rect 412674 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 413294 270014
rect 412674 234334 413294 269778
rect 412674 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 413294 234334
rect 412674 234014 413294 234098
rect 412674 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 413294 234014
rect 412674 198334 413294 233778
rect 412674 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 413294 198334
rect 412674 198014 413294 198098
rect 412674 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 413294 198014
rect 412674 162334 413294 197778
rect 412674 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 413294 162334
rect 412674 162014 413294 162098
rect 412674 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 413294 162014
rect 412674 126334 413294 161778
rect 412674 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 413294 126334
rect 412674 126014 413294 126098
rect 412674 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 413294 126014
rect 412674 90334 413294 125778
rect 412674 90098 412706 90334
rect 412942 90098 413026 90334
rect 413262 90098 413294 90334
rect 412674 90014 413294 90098
rect 412674 89778 412706 90014
rect 412942 89778 413026 90014
rect 413262 89778 413294 90014
rect 412674 54334 413294 89778
rect 412674 54098 412706 54334
rect 412942 54098 413026 54334
rect 413262 54098 413294 54334
rect 412674 54014 413294 54098
rect 412674 53778 412706 54014
rect 412942 53778 413026 54014
rect 413262 53778 413294 54014
rect 412674 18334 413294 53778
rect 412674 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 413294 18334
rect 412674 18014 413294 18098
rect 412674 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 413294 18014
rect 412674 -4186 413294 17778
rect 412674 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 413294 -4186
rect 412674 -4506 413294 -4422
rect 412674 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 413294 -4506
rect 412674 -7654 413294 -4742
rect 416394 709638 417014 711590
rect 416394 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 417014 709638
rect 416394 709318 417014 709402
rect 416394 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 417014 709318
rect 416394 670054 417014 709082
rect 416394 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 417014 670054
rect 416394 669734 417014 669818
rect 416394 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 417014 669734
rect 416394 634054 417014 669498
rect 416394 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 417014 634054
rect 416394 633734 417014 633818
rect 416394 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 417014 633734
rect 416394 598054 417014 633498
rect 416394 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 417014 598054
rect 416394 597734 417014 597818
rect 416394 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 417014 597734
rect 416394 562054 417014 597498
rect 416394 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 417014 562054
rect 416394 561734 417014 561818
rect 416394 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 417014 561734
rect 416394 526054 417014 561498
rect 416394 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 417014 526054
rect 416394 525734 417014 525818
rect 416394 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 417014 525734
rect 416394 490054 417014 525498
rect 416394 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 417014 490054
rect 416394 489734 417014 489818
rect 416394 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 417014 489734
rect 416394 454054 417014 489498
rect 416394 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 417014 454054
rect 416394 453734 417014 453818
rect 416394 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 417014 453734
rect 416394 418054 417014 453498
rect 416394 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 417014 418054
rect 416394 417734 417014 417818
rect 416394 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 417014 417734
rect 416394 382054 417014 417498
rect 416394 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 417014 382054
rect 416394 381734 417014 381818
rect 416394 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 417014 381734
rect 416394 346054 417014 381498
rect 416394 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 417014 346054
rect 416394 345734 417014 345818
rect 416394 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 417014 345734
rect 416394 310054 417014 345498
rect 416394 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 417014 310054
rect 416394 309734 417014 309818
rect 416394 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 417014 309734
rect 416394 274054 417014 309498
rect 416394 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 417014 274054
rect 416394 273734 417014 273818
rect 416394 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 417014 273734
rect 416394 238054 417014 273498
rect 416394 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 417014 238054
rect 416394 237734 417014 237818
rect 416394 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 417014 237734
rect 416394 202054 417014 237498
rect 416394 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 417014 202054
rect 416394 201734 417014 201818
rect 416394 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 417014 201734
rect 416394 166054 417014 201498
rect 416394 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 417014 166054
rect 416394 165734 417014 165818
rect 416394 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 417014 165734
rect 416394 130054 417014 165498
rect 416394 129818 416426 130054
rect 416662 129818 416746 130054
rect 416982 129818 417014 130054
rect 416394 129734 417014 129818
rect 416394 129498 416426 129734
rect 416662 129498 416746 129734
rect 416982 129498 417014 129734
rect 416394 94054 417014 129498
rect 416394 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 417014 94054
rect 416394 93734 417014 93818
rect 416394 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 417014 93734
rect 416394 58054 417014 93498
rect 416394 57818 416426 58054
rect 416662 57818 416746 58054
rect 416982 57818 417014 58054
rect 416394 57734 417014 57818
rect 416394 57498 416426 57734
rect 416662 57498 416746 57734
rect 416982 57498 417014 57734
rect 416394 22054 417014 57498
rect 416394 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 417014 22054
rect 416394 21734 417014 21818
rect 416394 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 417014 21734
rect 416394 -5146 417014 21498
rect 416394 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 417014 -5146
rect 416394 -5466 417014 -5382
rect 416394 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 417014 -5466
rect 416394 -7654 417014 -5702
rect 420114 710598 420734 711590
rect 420114 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 420734 710598
rect 420114 710278 420734 710362
rect 420114 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 420734 710278
rect 420114 673774 420734 710042
rect 420114 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 420734 673774
rect 420114 673454 420734 673538
rect 420114 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 420734 673454
rect 420114 637774 420734 673218
rect 420114 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 420734 637774
rect 420114 637454 420734 637538
rect 420114 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 420734 637454
rect 420114 601774 420734 637218
rect 420114 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 420734 601774
rect 420114 601454 420734 601538
rect 420114 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 420734 601454
rect 420114 565774 420734 601218
rect 420114 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 420734 565774
rect 420114 565454 420734 565538
rect 420114 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 420734 565454
rect 420114 529774 420734 565218
rect 420114 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 420734 529774
rect 420114 529454 420734 529538
rect 420114 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 420734 529454
rect 420114 493774 420734 529218
rect 420114 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 420734 493774
rect 420114 493454 420734 493538
rect 420114 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 420734 493454
rect 420114 457774 420734 493218
rect 420114 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 420734 457774
rect 420114 457454 420734 457538
rect 420114 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 420734 457454
rect 420114 421774 420734 457218
rect 420114 421538 420146 421774
rect 420382 421538 420466 421774
rect 420702 421538 420734 421774
rect 420114 421454 420734 421538
rect 420114 421218 420146 421454
rect 420382 421218 420466 421454
rect 420702 421218 420734 421454
rect 420114 385774 420734 421218
rect 420114 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 420734 385774
rect 420114 385454 420734 385538
rect 420114 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 420734 385454
rect 420114 349774 420734 385218
rect 420114 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 420734 349774
rect 420114 349454 420734 349538
rect 420114 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 420734 349454
rect 420114 313774 420734 349218
rect 420114 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 420734 313774
rect 420114 313454 420734 313538
rect 420114 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 420734 313454
rect 420114 277774 420734 313218
rect 420114 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 420734 277774
rect 420114 277454 420734 277538
rect 420114 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 420734 277454
rect 420114 241774 420734 277218
rect 420114 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 420734 241774
rect 420114 241454 420734 241538
rect 420114 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 420734 241454
rect 420114 205774 420734 241218
rect 420114 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 420734 205774
rect 420114 205454 420734 205538
rect 420114 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 420734 205454
rect 420114 169774 420734 205218
rect 420114 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 420734 169774
rect 420114 169454 420734 169538
rect 420114 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 420734 169454
rect 420114 133774 420734 169218
rect 420114 133538 420146 133774
rect 420382 133538 420466 133774
rect 420702 133538 420734 133774
rect 420114 133454 420734 133538
rect 420114 133218 420146 133454
rect 420382 133218 420466 133454
rect 420702 133218 420734 133454
rect 420114 97774 420734 133218
rect 420114 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 420734 97774
rect 420114 97454 420734 97538
rect 420114 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 420734 97454
rect 420114 61774 420734 97218
rect 420114 61538 420146 61774
rect 420382 61538 420466 61774
rect 420702 61538 420734 61774
rect 420114 61454 420734 61538
rect 420114 61218 420146 61454
rect 420382 61218 420466 61454
rect 420702 61218 420734 61454
rect 420114 25774 420734 61218
rect 420114 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 420734 25774
rect 420114 25454 420734 25538
rect 420114 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 420734 25454
rect 420114 -6106 420734 25218
rect 420114 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 420734 -6106
rect 420114 -6426 420734 -6342
rect 420114 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 420734 -6426
rect 420114 -7654 420734 -6662
rect 423834 711558 424454 711590
rect 423834 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 424454 711558
rect 423834 711238 424454 711322
rect 423834 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 424454 711238
rect 423834 677494 424454 711002
rect 423834 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 424454 677494
rect 423834 677174 424454 677258
rect 423834 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 424454 677174
rect 423834 641494 424454 676938
rect 423834 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 424454 641494
rect 423834 641174 424454 641258
rect 423834 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 424454 641174
rect 423834 605494 424454 640938
rect 423834 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 424454 605494
rect 423834 605174 424454 605258
rect 423834 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 424454 605174
rect 423834 569494 424454 604938
rect 423834 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 424454 569494
rect 423834 569174 424454 569258
rect 423834 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 424454 569174
rect 423834 533494 424454 568938
rect 423834 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 424454 533494
rect 423834 533174 424454 533258
rect 423834 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 424454 533174
rect 423834 497494 424454 532938
rect 423834 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 424454 497494
rect 423834 497174 424454 497258
rect 423834 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 424454 497174
rect 423834 461494 424454 496938
rect 423834 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 424454 461494
rect 423834 461174 424454 461258
rect 423834 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 424454 461174
rect 423834 425494 424454 460938
rect 423834 425258 423866 425494
rect 424102 425258 424186 425494
rect 424422 425258 424454 425494
rect 423834 425174 424454 425258
rect 423834 424938 423866 425174
rect 424102 424938 424186 425174
rect 424422 424938 424454 425174
rect 423834 389494 424454 424938
rect 423834 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 424454 389494
rect 423834 389174 424454 389258
rect 423834 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 424454 389174
rect 423834 353494 424454 388938
rect 423834 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 424454 353494
rect 423834 353174 424454 353258
rect 423834 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 424454 353174
rect 423834 317494 424454 352938
rect 423834 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 424454 317494
rect 423834 317174 424454 317258
rect 423834 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 424454 317174
rect 423834 281494 424454 316938
rect 423834 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 424454 281494
rect 423834 281174 424454 281258
rect 423834 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 424454 281174
rect 423834 245494 424454 280938
rect 423834 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 424454 245494
rect 423834 245174 424454 245258
rect 423834 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 424454 245174
rect 423834 209494 424454 244938
rect 423834 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 424454 209494
rect 423834 209174 424454 209258
rect 423834 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 424454 209174
rect 423834 173494 424454 208938
rect 423834 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 424454 173494
rect 423834 173174 424454 173258
rect 423834 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 424454 173174
rect 423834 137494 424454 172938
rect 423834 137258 423866 137494
rect 424102 137258 424186 137494
rect 424422 137258 424454 137494
rect 423834 137174 424454 137258
rect 423834 136938 423866 137174
rect 424102 136938 424186 137174
rect 424422 136938 424454 137174
rect 423834 101494 424454 136938
rect 423834 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 424454 101494
rect 423834 101174 424454 101258
rect 423834 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 424454 101174
rect 423834 65494 424454 100938
rect 423834 65258 423866 65494
rect 424102 65258 424186 65494
rect 424422 65258 424454 65494
rect 423834 65174 424454 65258
rect 423834 64938 423866 65174
rect 424102 64938 424186 65174
rect 424422 64938 424454 65174
rect 423834 29494 424454 64938
rect 423834 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 424454 29494
rect 423834 29174 424454 29258
rect 423834 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 424454 29174
rect 423834 -7066 424454 28938
rect 423834 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 424454 -7066
rect 423834 -7386 424454 -7302
rect 423834 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 424454 -7386
rect 423834 -7654 424454 -7622
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 437514 705798 438134 711590
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 691174 438134 705242
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -7654 438134 -1862
rect 441234 706758 441854 711590
rect 441234 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 441854 706758
rect 441234 706438 441854 706522
rect 441234 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 441854 706438
rect 441234 694894 441854 706202
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -2266 441854 10338
rect 441234 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 441854 -2266
rect 441234 -2586 441854 -2502
rect 441234 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 441854 -2586
rect 441234 -7654 441854 -2822
rect 444954 707718 445574 711590
rect 444954 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 445574 707718
rect 444954 707398 445574 707482
rect 444954 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 445574 707398
rect 444954 698614 445574 707162
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 444954 -3226 445574 14058
rect 444954 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 445574 -3226
rect 444954 -3546 445574 -3462
rect 444954 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 445574 -3546
rect 444954 -7654 445574 -3782
rect 448674 708678 449294 711590
rect 448674 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 449294 708678
rect 448674 708358 449294 708442
rect 448674 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 449294 708358
rect 448674 666334 449294 708122
rect 448674 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 449294 666334
rect 448674 666014 449294 666098
rect 448674 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 449294 666014
rect 448674 630334 449294 665778
rect 448674 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 449294 630334
rect 448674 630014 449294 630098
rect 448674 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 449294 630014
rect 448674 594334 449294 629778
rect 448674 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 449294 594334
rect 448674 594014 449294 594098
rect 448674 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 449294 594014
rect 448674 558334 449294 593778
rect 448674 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 449294 558334
rect 448674 558014 449294 558098
rect 448674 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 449294 558014
rect 448674 522334 449294 557778
rect 448674 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 449294 522334
rect 448674 522014 449294 522098
rect 448674 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 449294 522014
rect 448674 486334 449294 521778
rect 448674 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 449294 486334
rect 448674 486014 449294 486098
rect 448674 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 449294 486014
rect 448674 450334 449294 485778
rect 448674 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 449294 450334
rect 448674 450014 449294 450098
rect 448674 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 449294 450014
rect 448674 414334 449294 449778
rect 448674 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 449294 414334
rect 448674 414014 449294 414098
rect 448674 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 449294 414014
rect 448674 378334 449294 413778
rect 448674 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 449294 378334
rect 448674 378014 449294 378098
rect 448674 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 449294 378014
rect 448674 342334 449294 377778
rect 448674 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 449294 342334
rect 448674 342014 449294 342098
rect 448674 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 449294 342014
rect 448674 306334 449294 341778
rect 448674 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 449294 306334
rect 448674 306014 449294 306098
rect 448674 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 449294 306014
rect 448674 270334 449294 305778
rect 448674 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 449294 270334
rect 448674 270014 449294 270098
rect 448674 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 449294 270014
rect 448674 234334 449294 269778
rect 448674 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 449294 234334
rect 448674 234014 449294 234098
rect 448674 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 449294 234014
rect 448674 198334 449294 233778
rect 448674 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 449294 198334
rect 448674 198014 449294 198098
rect 448674 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 449294 198014
rect 448674 162334 449294 197778
rect 448674 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 449294 162334
rect 448674 162014 449294 162098
rect 448674 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 449294 162014
rect 448674 126334 449294 161778
rect 448674 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 449294 126334
rect 448674 126014 449294 126098
rect 448674 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 449294 126014
rect 448674 90334 449294 125778
rect 448674 90098 448706 90334
rect 448942 90098 449026 90334
rect 449262 90098 449294 90334
rect 448674 90014 449294 90098
rect 448674 89778 448706 90014
rect 448942 89778 449026 90014
rect 449262 89778 449294 90014
rect 448674 54334 449294 89778
rect 448674 54098 448706 54334
rect 448942 54098 449026 54334
rect 449262 54098 449294 54334
rect 448674 54014 449294 54098
rect 448674 53778 448706 54014
rect 448942 53778 449026 54014
rect 449262 53778 449294 54014
rect 448674 18334 449294 53778
rect 448674 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 449294 18334
rect 448674 18014 449294 18098
rect 448674 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 449294 18014
rect 448674 -4186 449294 17778
rect 448674 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 449294 -4186
rect 448674 -4506 449294 -4422
rect 448674 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 449294 -4506
rect 448674 -7654 449294 -4742
rect 452394 709638 453014 711590
rect 452394 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 453014 709638
rect 452394 709318 453014 709402
rect 452394 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 453014 709318
rect 452394 670054 453014 709082
rect 452394 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 453014 670054
rect 452394 669734 453014 669818
rect 452394 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 453014 669734
rect 452394 634054 453014 669498
rect 452394 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 453014 634054
rect 452394 633734 453014 633818
rect 452394 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 453014 633734
rect 452394 598054 453014 633498
rect 452394 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 453014 598054
rect 452394 597734 453014 597818
rect 452394 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 453014 597734
rect 452394 562054 453014 597498
rect 452394 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 453014 562054
rect 452394 561734 453014 561818
rect 452394 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 453014 561734
rect 452394 526054 453014 561498
rect 452394 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 453014 526054
rect 452394 525734 453014 525818
rect 452394 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 453014 525734
rect 452394 490054 453014 525498
rect 452394 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 453014 490054
rect 452394 489734 453014 489818
rect 452394 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 453014 489734
rect 452394 454054 453014 489498
rect 452394 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 453818 453014 454054
rect 452394 453734 453014 453818
rect 452394 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 453014 453734
rect 452394 418054 453014 453498
rect 452394 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 453014 418054
rect 452394 417734 453014 417818
rect 452394 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 453014 417734
rect 452394 382054 453014 417498
rect 452394 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 453014 382054
rect 452394 381734 453014 381818
rect 452394 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 453014 381734
rect 452394 346054 453014 381498
rect 452394 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 453014 346054
rect 452394 345734 453014 345818
rect 452394 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 453014 345734
rect 452394 310054 453014 345498
rect 452394 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 453014 310054
rect 452394 309734 453014 309818
rect 452394 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 453014 309734
rect 452394 274054 453014 309498
rect 452394 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 453014 274054
rect 452394 273734 453014 273818
rect 452394 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 453014 273734
rect 452394 238054 453014 273498
rect 452394 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 453014 238054
rect 452394 237734 453014 237818
rect 452394 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 453014 237734
rect 452394 202054 453014 237498
rect 452394 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 453014 202054
rect 452394 201734 453014 201818
rect 452394 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 453014 201734
rect 452394 166054 453014 201498
rect 452394 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 453014 166054
rect 452394 165734 453014 165818
rect 452394 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 453014 165734
rect 452394 130054 453014 165498
rect 452394 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 453014 130054
rect 452394 129734 453014 129818
rect 452394 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 453014 129734
rect 452394 94054 453014 129498
rect 452394 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 453014 94054
rect 452394 93734 453014 93818
rect 452394 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 453014 93734
rect 452394 58054 453014 93498
rect 452394 57818 452426 58054
rect 452662 57818 452746 58054
rect 452982 57818 453014 58054
rect 452394 57734 453014 57818
rect 452394 57498 452426 57734
rect 452662 57498 452746 57734
rect 452982 57498 453014 57734
rect 452394 22054 453014 57498
rect 452394 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 453014 22054
rect 452394 21734 453014 21818
rect 452394 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 453014 21734
rect 452394 -5146 453014 21498
rect 452394 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 453014 -5146
rect 452394 -5466 453014 -5382
rect 452394 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 453014 -5466
rect 452394 -7654 453014 -5702
rect 456114 710598 456734 711590
rect 456114 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 456734 710598
rect 456114 710278 456734 710362
rect 456114 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 456734 710278
rect 456114 673774 456734 710042
rect 456114 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 456734 673774
rect 456114 673454 456734 673538
rect 456114 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 456734 673454
rect 456114 637774 456734 673218
rect 456114 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 456734 637774
rect 456114 637454 456734 637538
rect 456114 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 456734 637454
rect 456114 601774 456734 637218
rect 456114 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 456734 601774
rect 456114 601454 456734 601538
rect 456114 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 456734 601454
rect 456114 565774 456734 601218
rect 456114 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 456734 565774
rect 456114 565454 456734 565538
rect 456114 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 456734 565454
rect 456114 529774 456734 565218
rect 456114 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 456734 529774
rect 456114 529454 456734 529538
rect 456114 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 456734 529454
rect 456114 493774 456734 529218
rect 456114 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 456734 493774
rect 456114 493454 456734 493538
rect 456114 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 456734 493454
rect 456114 457774 456734 493218
rect 456114 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 456734 457774
rect 456114 457454 456734 457538
rect 456114 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 456734 457454
rect 456114 421774 456734 457218
rect 456114 421538 456146 421774
rect 456382 421538 456466 421774
rect 456702 421538 456734 421774
rect 456114 421454 456734 421538
rect 456114 421218 456146 421454
rect 456382 421218 456466 421454
rect 456702 421218 456734 421454
rect 456114 385774 456734 421218
rect 456114 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 456734 385774
rect 456114 385454 456734 385538
rect 456114 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 456734 385454
rect 456114 349774 456734 385218
rect 456114 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 456734 349774
rect 456114 349454 456734 349538
rect 456114 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 456734 349454
rect 456114 313774 456734 349218
rect 456114 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 456734 313774
rect 456114 313454 456734 313538
rect 456114 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 456734 313454
rect 456114 277774 456734 313218
rect 456114 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 456734 277774
rect 456114 277454 456734 277538
rect 456114 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 456734 277454
rect 456114 241774 456734 277218
rect 456114 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 456734 241774
rect 456114 241454 456734 241538
rect 456114 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 456734 241454
rect 459834 711558 460454 711590
rect 459834 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 460454 711558
rect 459834 711238 460454 711322
rect 459834 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 460454 711238
rect 459834 677494 460454 711002
rect 459834 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 460454 677494
rect 459834 677174 460454 677258
rect 459834 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 460454 677174
rect 459834 641494 460454 676938
rect 459834 641258 459866 641494
rect 460102 641258 460186 641494
rect 460422 641258 460454 641494
rect 459834 641174 460454 641258
rect 459834 640938 459866 641174
rect 460102 640938 460186 641174
rect 460422 640938 460454 641174
rect 459834 605494 460454 640938
rect 459834 605258 459866 605494
rect 460102 605258 460186 605494
rect 460422 605258 460454 605494
rect 459834 605174 460454 605258
rect 459834 604938 459866 605174
rect 460102 604938 460186 605174
rect 460422 604938 460454 605174
rect 459834 569494 460454 604938
rect 459834 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 460454 569494
rect 459834 569174 460454 569258
rect 459834 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 460454 569174
rect 459834 533494 460454 568938
rect 459834 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 460454 533494
rect 459834 533174 460454 533258
rect 459834 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 460454 533174
rect 459834 497494 460454 532938
rect 459834 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 460454 497494
rect 459834 497174 460454 497258
rect 459834 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 460454 497174
rect 459834 461494 460454 496938
rect 459834 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 460454 461494
rect 459834 461174 460454 461258
rect 459834 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 460454 461174
rect 459834 425494 460454 460938
rect 459834 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 460454 425494
rect 459834 425174 460454 425258
rect 459834 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 460454 425174
rect 459834 389494 460454 424938
rect 459834 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 460454 389494
rect 459834 389174 460454 389258
rect 459834 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 460454 389174
rect 459834 353494 460454 388938
rect 459834 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 460454 353494
rect 459834 353174 460454 353258
rect 459834 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 460454 353174
rect 459834 317494 460454 352938
rect 459834 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 460454 317494
rect 459834 317174 460454 317258
rect 459834 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 460454 317174
rect 459834 281494 460454 316938
rect 459834 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 460454 281494
rect 459834 281174 460454 281258
rect 459834 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 460454 281174
rect 459834 245494 460454 280938
rect 459834 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 460454 245494
rect 459834 245174 460454 245258
rect 459834 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 460454 245174
rect 456114 205774 456734 241218
rect 457299 241228 457365 241229
rect 457299 241164 457300 241228
rect 457364 241164 457365 241228
rect 457299 241163 457365 241164
rect 456114 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 456734 205774
rect 456114 205454 456734 205538
rect 456114 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 456734 205454
rect 456114 169774 456734 205218
rect 456114 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 456734 169774
rect 456114 169454 456734 169538
rect 456114 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 456734 169454
rect 456114 133774 456734 169218
rect 456114 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 456734 133774
rect 456114 133454 456734 133538
rect 456114 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 456734 133454
rect 456114 97774 456734 133218
rect 456114 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 456734 97774
rect 456114 97454 456734 97538
rect 456114 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 456734 97454
rect 456114 61774 456734 97218
rect 456114 61538 456146 61774
rect 456382 61538 456466 61774
rect 456702 61538 456734 61774
rect 456114 61454 456734 61538
rect 456114 61218 456146 61454
rect 456382 61218 456466 61454
rect 456702 61218 456734 61454
rect 456114 25774 456734 61218
rect 456114 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 456734 25774
rect 456114 25454 456734 25538
rect 456114 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 456734 25454
rect 456114 -6106 456734 25218
rect 457302 19821 457362 241163
rect 459834 209494 460454 244938
rect 459834 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 460454 209494
rect 459834 209174 460454 209258
rect 459834 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 460454 209174
rect 459834 173494 460454 208938
rect 459834 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 460454 173494
rect 459834 173174 460454 173258
rect 459834 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 460454 173174
rect 459834 137494 460454 172938
rect 459834 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 460454 137494
rect 459834 137174 460454 137258
rect 459834 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 460454 137174
rect 459834 101494 460454 136938
rect 459834 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 460454 101494
rect 459834 101174 460454 101258
rect 459834 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 460454 101174
rect 459834 65494 460454 100938
rect 459834 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 460454 65494
rect 459834 65174 460454 65258
rect 459834 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 460454 65174
rect 459834 29494 460454 64938
rect 459834 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 460454 29494
rect 459834 29174 460454 29258
rect 459834 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 460454 29174
rect 457299 19820 457365 19821
rect 457299 19756 457300 19820
rect 457364 19756 457365 19820
rect 457299 19755 457365 19756
rect 456114 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 456734 -6106
rect 456114 -6426 456734 -6342
rect 456114 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 456734 -6426
rect 456114 -7654 456734 -6662
rect 459834 -7066 460454 28938
rect 459834 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 460454 -7066
rect 459834 -7386 460454 -7302
rect 459834 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 460454 -7386
rect 459834 -7654 460454 -7622
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 473514 705798 474134 711590
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 691174 474134 705242
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -7654 474134 -1862
rect 477234 706758 477854 711590
rect 477234 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 477854 706758
rect 477234 706438 477854 706522
rect 477234 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 477854 706438
rect 477234 694894 477854 706202
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -2266 477854 10338
rect 477234 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 477854 -2266
rect 477234 -2586 477854 -2502
rect 477234 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 477854 -2586
rect 477234 -7654 477854 -2822
rect 480954 707718 481574 711590
rect 480954 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 481574 707718
rect 480954 707398 481574 707482
rect 480954 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 481574 707398
rect 480954 698614 481574 707162
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 480954 -3226 481574 14058
rect 480954 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 481574 -3226
rect 480954 -3546 481574 -3462
rect 480954 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 481574 -3546
rect 480954 -7654 481574 -3782
rect 484674 708678 485294 711590
rect 484674 708442 484706 708678
rect 484942 708442 485026 708678
rect 485262 708442 485294 708678
rect 484674 708358 485294 708442
rect 484674 708122 484706 708358
rect 484942 708122 485026 708358
rect 485262 708122 485294 708358
rect 484674 666334 485294 708122
rect 484674 666098 484706 666334
rect 484942 666098 485026 666334
rect 485262 666098 485294 666334
rect 484674 666014 485294 666098
rect 484674 665778 484706 666014
rect 484942 665778 485026 666014
rect 485262 665778 485294 666014
rect 484674 630334 485294 665778
rect 484674 630098 484706 630334
rect 484942 630098 485026 630334
rect 485262 630098 485294 630334
rect 484674 630014 485294 630098
rect 484674 629778 484706 630014
rect 484942 629778 485026 630014
rect 485262 629778 485294 630014
rect 484674 594334 485294 629778
rect 484674 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 485294 594334
rect 484674 594014 485294 594098
rect 484674 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 485294 594014
rect 484674 558334 485294 593778
rect 484674 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 485294 558334
rect 484674 558014 485294 558098
rect 484674 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 485294 558014
rect 484674 522334 485294 557778
rect 484674 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 485294 522334
rect 484674 522014 485294 522098
rect 484674 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 485294 522014
rect 484674 486334 485294 521778
rect 484674 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 485294 486334
rect 484674 486014 485294 486098
rect 484674 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 485294 486014
rect 484674 450334 485294 485778
rect 484674 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 485294 450334
rect 484674 450014 485294 450098
rect 484674 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 485294 450014
rect 484674 414334 485294 449778
rect 484674 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 485294 414334
rect 484674 414014 485294 414098
rect 484674 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 485294 414014
rect 484674 378334 485294 413778
rect 484674 378098 484706 378334
rect 484942 378098 485026 378334
rect 485262 378098 485294 378334
rect 484674 378014 485294 378098
rect 484674 377778 484706 378014
rect 484942 377778 485026 378014
rect 485262 377778 485294 378014
rect 484674 342334 485294 377778
rect 484674 342098 484706 342334
rect 484942 342098 485026 342334
rect 485262 342098 485294 342334
rect 484674 342014 485294 342098
rect 484674 341778 484706 342014
rect 484942 341778 485026 342014
rect 485262 341778 485294 342014
rect 484674 306334 485294 341778
rect 484674 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 485294 306334
rect 484674 306014 485294 306098
rect 484674 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 485294 306014
rect 484674 270334 485294 305778
rect 484674 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 485294 270334
rect 484674 270014 485294 270098
rect 484674 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 485294 270014
rect 484674 234334 485294 269778
rect 484674 234098 484706 234334
rect 484942 234098 485026 234334
rect 485262 234098 485294 234334
rect 484674 234014 485294 234098
rect 484674 233778 484706 234014
rect 484942 233778 485026 234014
rect 485262 233778 485294 234014
rect 484674 198334 485294 233778
rect 484674 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 485294 198334
rect 484674 198014 485294 198098
rect 484674 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 485294 198014
rect 484674 162334 485294 197778
rect 484674 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 485294 162334
rect 484674 162014 485294 162098
rect 484674 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 485294 162014
rect 484674 126334 485294 161778
rect 484674 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 485294 126334
rect 484674 126014 485294 126098
rect 484674 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 485294 126014
rect 484674 90334 485294 125778
rect 484674 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 485294 90334
rect 484674 90014 485294 90098
rect 484674 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 485294 90014
rect 484674 54334 485294 89778
rect 484674 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 485294 54334
rect 484674 54014 485294 54098
rect 484674 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 485294 54014
rect 484674 18334 485294 53778
rect 484674 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 485294 18334
rect 484674 18014 485294 18098
rect 484674 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 485294 18014
rect 484674 -4186 485294 17778
rect 484674 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 485294 -4186
rect 484674 -4506 485294 -4422
rect 484674 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 485294 -4506
rect 484674 -7654 485294 -4742
rect 488394 709638 489014 711590
rect 488394 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 489014 709638
rect 488394 709318 489014 709402
rect 488394 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 489014 709318
rect 488394 670054 489014 709082
rect 488394 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 489014 670054
rect 488394 669734 489014 669818
rect 488394 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 489014 669734
rect 488394 634054 489014 669498
rect 488394 633818 488426 634054
rect 488662 633818 488746 634054
rect 488982 633818 489014 634054
rect 488394 633734 489014 633818
rect 488394 633498 488426 633734
rect 488662 633498 488746 633734
rect 488982 633498 489014 633734
rect 488394 598054 489014 633498
rect 488394 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 489014 598054
rect 488394 597734 489014 597818
rect 488394 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 489014 597734
rect 488394 562054 489014 597498
rect 488394 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 489014 562054
rect 488394 561734 489014 561818
rect 488394 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 489014 561734
rect 488394 526054 489014 561498
rect 488394 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 489014 526054
rect 488394 525734 489014 525818
rect 488394 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 489014 525734
rect 488394 490054 489014 525498
rect 488394 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 489014 490054
rect 488394 489734 489014 489818
rect 488394 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 489014 489734
rect 488394 454054 489014 489498
rect 488394 453818 488426 454054
rect 488662 453818 488746 454054
rect 488982 453818 489014 454054
rect 488394 453734 489014 453818
rect 488394 453498 488426 453734
rect 488662 453498 488746 453734
rect 488982 453498 489014 453734
rect 488394 418054 489014 453498
rect 488394 417818 488426 418054
rect 488662 417818 488746 418054
rect 488982 417818 489014 418054
rect 488394 417734 489014 417818
rect 488394 417498 488426 417734
rect 488662 417498 488746 417734
rect 488982 417498 489014 417734
rect 488394 382054 489014 417498
rect 488394 381818 488426 382054
rect 488662 381818 488746 382054
rect 488982 381818 489014 382054
rect 488394 381734 489014 381818
rect 488394 381498 488426 381734
rect 488662 381498 488746 381734
rect 488982 381498 489014 381734
rect 488394 346054 489014 381498
rect 488394 345818 488426 346054
rect 488662 345818 488746 346054
rect 488982 345818 489014 346054
rect 488394 345734 489014 345818
rect 488394 345498 488426 345734
rect 488662 345498 488746 345734
rect 488982 345498 489014 345734
rect 488394 310054 489014 345498
rect 488394 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 489014 310054
rect 488394 309734 489014 309818
rect 488394 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 489014 309734
rect 488394 274054 489014 309498
rect 488394 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 489014 274054
rect 488394 273734 489014 273818
rect 488394 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 489014 273734
rect 488394 238054 489014 273498
rect 488394 237818 488426 238054
rect 488662 237818 488746 238054
rect 488982 237818 489014 238054
rect 488394 237734 489014 237818
rect 488394 237498 488426 237734
rect 488662 237498 488746 237734
rect 488982 237498 489014 237734
rect 488394 202054 489014 237498
rect 488394 201818 488426 202054
rect 488662 201818 488746 202054
rect 488982 201818 489014 202054
rect 488394 201734 489014 201818
rect 488394 201498 488426 201734
rect 488662 201498 488746 201734
rect 488982 201498 489014 201734
rect 488394 166054 489014 201498
rect 488394 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 489014 166054
rect 488394 165734 489014 165818
rect 488394 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 489014 165734
rect 488394 130054 489014 165498
rect 488394 129818 488426 130054
rect 488662 129818 488746 130054
rect 488982 129818 489014 130054
rect 488394 129734 489014 129818
rect 488394 129498 488426 129734
rect 488662 129498 488746 129734
rect 488982 129498 489014 129734
rect 488394 94054 489014 129498
rect 488394 93818 488426 94054
rect 488662 93818 488746 94054
rect 488982 93818 489014 94054
rect 488394 93734 489014 93818
rect 488394 93498 488426 93734
rect 488662 93498 488746 93734
rect 488982 93498 489014 93734
rect 488394 58054 489014 93498
rect 488394 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 489014 58054
rect 488394 57734 489014 57818
rect 488394 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 489014 57734
rect 488394 22054 489014 57498
rect 488394 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 489014 22054
rect 488394 21734 489014 21818
rect 488394 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 489014 21734
rect 488394 -5146 489014 21498
rect 488394 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 489014 -5146
rect 488394 -5466 489014 -5382
rect 488394 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 489014 -5466
rect 488394 -7654 489014 -5702
rect 492114 710598 492734 711590
rect 492114 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 492734 710598
rect 492114 710278 492734 710362
rect 492114 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 492734 710278
rect 492114 673774 492734 710042
rect 492114 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 492734 673774
rect 492114 673454 492734 673538
rect 492114 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 492734 673454
rect 492114 637774 492734 673218
rect 495834 711558 496454 711590
rect 495834 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 496454 711558
rect 495834 711238 496454 711322
rect 495834 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 496454 711238
rect 495834 677494 496454 711002
rect 495834 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 496454 677494
rect 495834 677174 496454 677258
rect 495834 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 496454 677174
rect 495834 654737 496454 676938
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 501643 655620 501709 655621
rect 501643 655556 501644 655620
rect 501708 655556 501709 655620
rect 501643 655555 501709 655556
rect 500355 654940 500421 654941
rect 500355 654876 500356 654940
rect 500420 654876 500421 654940
rect 500355 654875 500421 654876
rect 500358 653445 500418 654875
rect 501646 654397 501706 655555
rect 505794 654737 506414 686898
rect 509514 705798 510134 711590
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 691174 510134 705242
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 654956 510134 690618
rect 513234 706758 513854 711590
rect 513234 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 513854 706758
rect 513234 706438 513854 706522
rect 513234 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 513854 706438
rect 513234 694894 513854 706202
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 654737 513854 658338
rect 516954 707718 517574 711590
rect 516954 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 517574 707718
rect 516954 707398 517574 707482
rect 516954 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 517574 707398
rect 516954 698614 517574 707162
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 654737 517574 662058
rect 520674 708678 521294 711590
rect 520674 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 521294 708678
rect 520674 708358 521294 708442
rect 520674 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 521294 708358
rect 520674 666334 521294 708122
rect 520674 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 521294 666334
rect 520674 666014 521294 666098
rect 520674 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 521294 666014
rect 520674 654737 521294 665778
rect 524394 709638 525014 711590
rect 524394 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 525014 709638
rect 524394 709318 525014 709402
rect 524394 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 525014 709318
rect 524394 670054 525014 709082
rect 524394 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 525014 670054
rect 524394 669734 525014 669818
rect 524394 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 525014 669734
rect 524394 654956 525014 669498
rect 528114 710598 528734 711590
rect 528114 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 528734 710598
rect 528114 710278 528734 710362
rect 528114 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 528734 710278
rect 528114 673774 528734 710042
rect 528114 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 528734 673774
rect 528114 673454 528734 673538
rect 528114 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 528734 673454
rect 528114 654737 528734 673218
rect 531834 711558 532454 711590
rect 531834 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 532454 711558
rect 531834 711238 532454 711322
rect 531834 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 532454 711238
rect 531834 677494 532454 711002
rect 531834 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 532454 677494
rect 531834 677174 532454 677258
rect 531834 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 532454 677174
rect 531834 654737 532454 676938
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 501643 654396 501709 654397
rect 501643 654332 501644 654396
rect 501708 654332 501709 654396
rect 501643 654331 501709 654332
rect 500355 653444 500421 653445
rect 500355 653380 500356 653444
rect 500420 653380 500421 653444
rect 500355 653379 500421 653380
rect 494208 651454 494528 651486
rect 494208 651218 494250 651454
rect 494486 651218 494528 651454
rect 494208 651134 494528 651218
rect 494208 650898 494250 651134
rect 494486 650898 494528 651134
rect 494208 650866 494528 650898
rect 524928 651454 525248 651486
rect 524928 651218 524970 651454
rect 525206 651218 525248 651454
rect 524928 651134 525248 651218
rect 524928 650898 524970 651134
rect 525206 650898 525248 651134
rect 524928 650866 525248 650898
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 492114 637538 492146 637774
rect 492382 637538 492466 637774
rect 492702 637538 492734 637774
rect 492114 637454 492734 637538
rect 492114 637218 492146 637454
rect 492382 637218 492466 637454
rect 492702 637218 492734 637454
rect 492114 601774 492734 637218
rect 509568 619174 509888 619206
rect 509568 618938 509610 619174
rect 509846 618938 509888 619174
rect 509568 618854 509888 618938
rect 509568 618618 509610 618854
rect 509846 618618 509888 618854
rect 509568 618586 509888 618618
rect 541019 618628 541085 618629
rect 541019 618564 541020 618628
rect 541084 618564 541085 618628
rect 541019 618563 541085 618564
rect 494208 615454 494528 615486
rect 494208 615218 494250 615454
rect 494486 615218 494528 615454
rect 494208 615134 494528 615218
rect 494208 614898 494250 615134
rect 494486 614898 494528 615134
rect 494208 614866 494528 614898
rect 524928 615454 525248 615486
rect 524928 615218 524970 615454
rect 525206 615218 525248 615454
rect 524928 615134 525248 615218
rect 524928 614898 524970 615134
rect 525206 614898 525248 615134
rect 524928 614866 525248 614898
rect 539363 603668 539429 603669
rect 539363 603604 539364 603668
rect 539428 603604 539429 603668
rect 539363 603603 539429 603604
rect 492114 601538 492146 601774
rect 492382 601538 492466 601774
rect 492702 601538 492734 601774
rect 492114 601454 492734 601538
rect 492114 601218 492146 601454
rect 492382 601218 492466 601454
rect 492702 601218 492734 601454
rect 492114 565774 492734 601218
rect 492114 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 492734 565774
rect 492114 565454 492734 565538
rect 492114 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 492734 565454
rect 492114 529774 492734 565218
rect 492114 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 492734 529774
rect 492114 529454 492734 529538
rect 492114 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 492734 529454
rect 492114 493774 492734 529218
rect 492114 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 492734 493774
rect 492114 493454 492734 493538
rect 492114 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 492734 493454
rect 492114 457774 492734 493218
rect 492114 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 492734 457774
rect 492114 457454 492734 457538
rect 492114 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 492734 457454
rect 492114 421774 492734 457218
rect 492114 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 492734 421774
rect 492114 421454 492734 421538
rect 492114 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 492734 421454
rect 492114 385774 492734 421218
rect 492114 385538 492146 385774
rect 492382 385538 492466 385774
rect 492702 385538 492734 385774
rect 492114 385454 492734 385538
rect 492114 385218 492146 385454
rect 492382 385218 492466 385454
rect 492702 385218 492734 385454
rect 492114 349774 492734 385218
rect 492114 349538 492146 349774
rect 492382 349538 492466 349774
rect 492702 349538 492734 349774
rect 492114 349454 492734 349538
rect 492114 349218 492146 349454
rect 492382 349218 492466 349454
rect 492702 349218 492734 349454
rect 492114 313774 492734 349218
rect 492114 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 492734 313774
rect 492114 313454 492734 313538
rect 492114 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 492734 313454
rect 492114 277774 492734 313218
rect 492114 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 492734 277774
rect 492114 277454 492734 277538
rect 492114 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 492734 277454
rect 492114 241774 492734 277218
rect 492114 241538 492146 241774
rect 492382 241538 492466 241774
rect 492702 241538 492734 241774
rect 492114 241454 492734 241538
rect 492114 241218 492146 241454
rect 492382 241218 492466 241454
rect 492702 241218 492734 241454
rect 492114 205774 492734 241218
rect 492114 205538 492146 205774
rect 492382 205538 492466 205774
rect 492702 205538 492734 205774
rect 492114 205454 492734 205538
rect 492114 205218 492146 205454
rect 492382 205218 492466 205454
rect 492702 205218 492734 205454
rect 492114 169774 492734 205218
rect 492114 169538 492146 169774
rect 492382 169538 492466 169774
rect 492702 169538 492734 169774
rect 492114 169454 492734 169538
rect 492114 169218 492146 169454
rect 492382 169218 492466 169454
rect 492702 169218 492734 169454
rect 492114 133774 492734 169218
rect 492114 133538 492146 133774
rect 492382 133538 492466 133774
rect 492702 133538 492734 133774
rect 492114 133454 492734 133538
rect 492114 133218 492146 133454
rect 492382 133218 492466 133454
rect 492702 133218 492734 133454
rect 492114 97774 492734 133218
rect 492114 97538 492146 97774
rect 492382 97538 492466 97774
rect 492702 97538 492734 97774
rect 492114 97454 492734 97538
rect 492114 97218 492146 97454
rect 492382 97218 492466 97454
rect 492702 97218 492734 97454
rect 492114 61774 492734 97218
rect 492114 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 492734 61774
rect 492114 61454 492734 61538
rect 492114 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 492734 61454
rect 492114 25774 492734 61218
rect 492114 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 492734 25774
rect 492114 25454 492734 25538
rect 492114 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 492734 25454
rect 492114 -6106 492734 25218
rect 492114 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 492734 -6106
rect 492114 -6426 492734 -6342
rect 492114 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 492734 -6426
rect 492114 -7654 492734 -6662
rect 495834 569494 496454 600207
rect 495834 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 496454 569494
rect 495834 569174 496454 569258
rect 495834 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 496454 569174
rect 495834 533494 496454 568938
rect 495834 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 496454 533494
rect 495834 533174 496454 533258
rect 495834 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 496454 533174
rect 495834 497494 496454 532938
rect 495834 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 496454 497494
rect 495834 497174 496454 497258
rect 495834 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 496454 497174
rect 495834 461494 496454 496938
rect 495834 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 496454 461494
rect 495834 461174 496454 461258
rect 495834 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 496454 461174
rect 495834 425494 496454 460938
rect 495834 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 496454 425494
rect 495834 425174 496454 425258
rect 495834 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 496454 425174
rect 495834 389494 496454 424938
rect 505794 579454 506414 600207
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 500171 418300 500237 418301
rect 500171 418236 500172 418300
rect 500236 418236 500237 418300
rect 500171 418235 500237 418236
rect 495834 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 496454 389494
rect 495834 389174 496454 389258
rect 495834 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 496454 389174
rect 495834 353494 496454 388938
rect 495834 353258 495866 353494
rect 496102 353258 496186 353494
rect 496422 353258 496454 353494
rect 495834 353174 496454 353258
rect 495834 352938 495866 353174
rect 496102 352938 496186 353174
rect 496422 352938 496454 353174
rect 495834 317494 496454 352938
rect 495834 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 496454 317494
rect 495834 317174 496454 317258
rect 495834 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 496454 317174
rect 495834 281494 496454 316938
rect 495834 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 496454 281494
rect 495834 281174 496454 281258
rect 495834 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 496454 281174
rect 495834 245494 496454 280938
rect 500174 253469 500234 418235
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 500171 253468 500237 253469
rect 500171 253404 500172 253468
rect 500236 253404 500237 253468
rect 500171 253403 500237 253404
rect 495834 245258 495866 245494
rect 496102 245258 496186 245494
rect 496422 245258 496454 245494
rect 495834 245174 496454 245258
rect 495834 244938 495866 245174
rect 496102 244938 496186 245174
rect 496422 244938 496454 245174
rect 495834 209494 496454 244938
rect 500171 243948 500237 243949
rect 500171 243884 500172 243948
rect 500236 243884 500237 243948
rect 500171 243883 500237 243884
rect 495834 209258 495866 209494
rect 496102 209258 496186 209494
rect 496422 209258 496454 209494
rect 495834 209174 496454 209258
rect 495834 208938 495866 209174
rect 496102 208938 496186 209174
rect 496422 208938 496454 209174
rect 495834 173494 496454 208938
rect 495834 173258 495866 173494
rect 496102 173258 496186 173494
rect 496422 173258 496454 173494
rect 495834 173174 496454 173258
rect 495834 172938 495866 173174
rect 496102 172938 496186 173174
rect 496422 172938 496454 173174
rect 495834 137494 496454 172938
rect 495834 137258 495866 137494
rect 496102 137258 496186 137494
rect 496422 137258 496454 137494
rect 495834 137174 496454 137258
rect 495834 136938 495866 137174
rect 496102 136938 496186 137174
rect 496422 136938 496454 137174
rect 495834 101494 496454 136938
rect 495834 101258 495866 101494
rect 496102 101258 496186 101494
rect 496422 101258 496454 101494
rect 495834 101174 496454 101258
rect 495834 100938 495866 101174
rect 496102 100938 496186 101174
rect 496422 100938 496454 101174
rect 495834 65494 496454 100938
rect 500174 99517 500234 243883
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 500171 99516 500237 99517
rect 500171 99452 500172 99516
rect 500236 99452 500237 99516
rect 500171 99451 500237 99452
rect 495834 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 496454 65494
rect 495834 65174 496454 65258
rect 495834 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 496454 65174
rect 495834 29494 496454 64938
rect 495834 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 496454 29494
rect 495834 29174 496454 29258
rect 495834 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 496454 29174
rect 495834 -7066 496454 28938
rect 495834 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 496454 -7066
rect 495834 -7386 496454 -7302
rect 495834 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 496454 -7386
rect 495834 -7654 496454 -7622
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 509514 583174 510134 599988
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -7654 510134 -1862
rect 513234 586894 513854 600207
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -2266 513854 10338
rect 513234 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 513854 -2266
rect 513234 -2586 513854 -2502
rect 513234 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 513854 -2586
rect 513234 -7654 513854 -2822
rect 516954 590614 517574 600207
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 516954 -3226 517574 14058
rect 516954 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 517574 -3226
rect 516954 -3546 517574 -3462
rect 516954 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 517574 -3546
rect 516954 -7654 517574 -3782
rect 520674 594334 521294 600207
rect 520674 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 521294 594334
rect 520674 594014 521294 594098
rect 520674 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 521294 594014
rect 520674 558334 521294 593778
rect 520674 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 521294 558334
rect 520674 558014 521294 558098
rect 520674 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 521294 558014
rect 520674 522334 521294 557778
rect 520674 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 521294 522334
rect 520674 522014 521294 522098
rect 520674 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 521294 522014
rect 520674 486334 521294 521778
rect 520674 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 521294 486334
rect 520674 486014 521294 486098
rect 520674 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 521294 486014
rect 520674 450334 521294 485778
rect 520674 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 521294 450334
rect 520674 450014 521294 450098
rect 520674 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 521294 450014
rect 520674 414334 521294 449778
rect 520674 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 521294 414334
rect 520674 414014 521294 414098
rect 520674 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 521294 414014
rect 520674 378334 521294 413778
rect 520674 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 521294 378334
rect 520674 378014 521294 378098
rect 520674 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 521294 378014
rect 520674 342334 521294 377778
rect 520674 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 521294 342334
rect 520674 342014 521294 342098
rect 520674 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 521294 342014
rect 520674 306334 521294 341778
rect 520674 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 521294 306334
rect 520674 306014 521294 306098
rect 520674 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 521294 306014
rect 520674 270334 521294 305778
rect 520674 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 521294 270334
rect 520674 270014 521294 270098
rect 520674 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 521294 270014
rect 520674 234334 521294 269778
rect 520674 234098 520706 234334
rect 520942 234098 521026 234334
rect 521262 234098 521294 234334
rect 520674 234014 521294 234098
rect 520674 233778 520706 234014
rect 520942 233778 521026 234014
rect 521262 233778 521294 234014
rect 520674 198334 521294 233778
rect 520674 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 521294 198334
rect 520674 198014 521294 198098
rect 520674 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 521294 198014
rect 520674 162334 521294 197778
rect 520674 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 521294 162334
rect 520674 162014 521294 162098
rect 520674 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 521294 162014
rect 520674 126334 521294 161778
rect 520674 126098 520706 126334
rect 520942 126098 521026 126334
rect 521262 126098 521294 126334
rect 520674 126014 521294 126098
rect 520674 125778 520706 126014
rect 520942 125778 521026 126014
rect 521262 125778 521294 126014
rect 520674 90334 521294 125778
rect 520674 90098 520706 90334
rect 520942 90098 521026 90334
rect 521262 90098 521294 90334
rect 520674 90014 521294 90098
rect 520674 89778 520706 90014
rect 520942 89778 521026 90014
rect 521262 89778 521294 90014
rect 520674 54334 521294 89778
rect 520674 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 521294 54334
rect 520674 54014 521294 54098
rect 520674 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 521294 54014
rect 520674 18334 521294 53778
rect 520674 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 521294 18334
rect 520674 18014 521294 18098
rect 520674 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 521294 18014
rect 520674 -4186 521294 17778
rect 520674 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 521294 -4186
rect 520674 -4506 521294 -4422
rect 520674 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 521294 -4506
rect 520674 -7654 521294 -4742
rect 524394 598054 525014 599988
rect 524394 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 525014 598054
rect 524394 597734 525014 597818
rect 524394 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 525014 597734
rect 524394 562054 525014 597498
rect 524394 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 525014 562054
rect 524394 561734 525014 561818
rect 524394 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 525014 561734
rect 524394 526054 525014 561498
rect 524394 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 525014 526054
rect 524394 525734 525014 525818
rect 524394 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 525014 525734
rect 524394 490054 525014 525498
rect 524394 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 525014 490054
rect 524394 489734 525014 489818
rect 524394 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 525014 489734
rect 524394 454054 525014 489498
rect 524394 453818 524426 454054
rect 524662 453818 524746 454054
rect 524982 453818 525014 454054
rect 524394 453734 525014 453818
rect 524394 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 525014 453734
rect 524394 418054 525014 453498
rect 524394 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 525014 418054
rect 524394 417734 525014 417818
rect 524394 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 525014 417734
rect 524394 382054 525014 417498
rect 524394 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 525014 382054
rect 524394 381734 525014 381818
rect 524394 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 525014 381734
rect 524394 346054 525014 381498
rect 524394 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 525014 346054
rect 524394 345734 525014 345818
rect 524394 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 525014 345734
rect 524394 310054 525014 345498
rect 524394 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 525014 310054
rect 524394 309734 525014 309818
rect 524394 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 525014 309734
rect 524394 274054 525014 309498
rect 524394 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 525014 274054
rect 524394 273734 525014 273818
rect 524394 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 525014 273734
rect 524394 238054 525014 273498
rect 524394 237818 524426 238054
rect 524662 237818 524746 238054
rect 524982 237818 525014 238054
rect 524394 237734 525014 237818
rect 524394 237498 524426 237734
rect 524662 237498 524746 237734
rect 524982 237498 525014 237734
rect 524394 202054 525014 237498
rect 524394 201818 524426 202054
rect 524662 201818 524746 202054
rect 524982 201818 525014 202054
rect 524394 201734 525014 201818
rect 524394 201498 524426 201734
rect 524662 201498 524746 201734
rect 524982 201498 525014 201734
rect 524394 166054 525014 201498
rect 524394 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 525014 166054
rect 524394 165734 525014 165818
rect 524394 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 525014 165734
rect 524394 130054 525014 165498
rect 524394 129818 524426 130054
rect 524662 129818 524746 130054
rect 524982 129818 525014 130054
rect 524394 129734 525014 129818
rect 524394 129498 524426 129734
rect 524662 129498 524746 129734
rect 524982 129498 525014 129734
rect 524394 94054 525014 129498
rect 524394 93818 524426 94054
rect 524662 93818 524746 94054
rect 524982 93818 525014 94054
rect 524394 93734 525014 93818
rect 524394 93498 524426 93734
rect 524662 93498 524746 93734
rect 524982 93498 525014 93734
rect 524394 58054 525014 93498
rect 524394 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 525014 58054
rect 524394 57734 525014 57818
rect 524394 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 525014 57734
rect 524394 22054 525014 57498
rect 524394 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 525014 22054
rect 524394 21734 525014 21818
rect 524394 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 525014 21734
rect 524394 -5146 525014 21498
rect 524394 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 525014 -5146
rect 524394 -5466 525014 -5382
rect 524394 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 525014 -5466
rect 524394 -7654 525014 -5702
rect 528114 565774 528734 600207
rect 528114 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 528734 565774
rect 528114 565454 528734 565538
rect 528114 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 528734 565454
rect 528114 529774 528734 565218
rect 528114 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 528734 529774
rect 528114 529454 528734 529538
rect 528114 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 528734 529454
rect 528114 493774 528734 529218
rect 528114 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 528734 493774
rect 528114 493454 528734 493538
rect 528114 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 528734 493454
rect 528114 457774 528734 493218
rect 528114 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 528734 457774
rect 528114 457454 528734 457538
rect 528114 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 528734 457454
rect 528114 421774 528734 457218
rect 528114 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 528734 421774
rect 528114 421454 528734 421538
rect 528114 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 528734 421454
rect 528114 385774 528734 421218
rect 528114 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 528734 385774
rect 528114 385454 528734 385538
rect 528114 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 528734 385454
rect 528114 349774 528734 385218
rect 528114 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 528734 349774
rect 528114 349454 528734 349538
rect 528114 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 528734 349454
rect 528114 313774 528734 349218
rect 528114 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 528734 313774
rect 528114 313454 528734 313538
rect 528114 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 528734 313454
rect 528114 277774 528734 313218
rect 528114 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 528734 277774
rect 528114 277454 528734 277538
rect 528114 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 528734 277454
rect 528114 241774 528734 277218
rect 528114 241538 528146 241774
rect 528382 241538 528466 241774
rect 528702 241538 528734 241774
rect 528114 241454 528734 241538
rect 528114 241218 528146 241454
rect 528382 241218 528466 241454
rect 528702 241218 528734 241454
rect 528114 205774 528734 241218
rect 528114 205538 528146 205774
rect 528382 205538 528466 205774
rect 528702 205538 528734 205774
rect 528114 205454 528734 205538
rect 528114 205218 528146 205454
rect 528382 205218 528466 205454
rect 528702 205218 528734 205454
rect 528114 169774 528734 205218
rect 528114 169538 528146 169774
rect 528382 169538 528466 169774
rect 528702 169538 528734 169774
rect 528114 169454 528734 169538
rect 528114 169218 528146 169454
rect 528382 169218 528466 169454
rect 528702 169218 528734 169454
rect 528114 133774 528734 169218
rect 528114 133538 528146 133774
rect 528382 133538 528466 133774
rect 528702 133538 528734 133774
rect 528114 133454 528734 133538
rect 528114 133218 528146 133454
rect 528382 133218 528466 133454
rect 528702 133218 528734 133454
rect 528114 97774 528734 133218
rect 528114 97538 528146 97774
rect 528382 97538 528466 97774
rect 528702 97538 528734 97774
rect 528114 97454 528734 97538
rect 528114 97218 528146 97454
rect 528382 97218 528466 97454
rect 528702 97218 528734 97454
rect 528114 61774 528734 97218
rect 528114 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 528734 61774
rect 528114 61454 528734 61538
rect 528114 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 528734 61454
rect 528114 25774 528734 61218
rect 528114 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 528734 25774
rect 528114 25454 528734 25538
rect 528114 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 528734 25454
rect 528114 -6106 528734 25218
rect 528114 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 528734 -6106
rect 528114 -6426 528734 -6342
rect 528114 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 528734 -6426
rect 528114 -7654 528734 -6662
rect 531834 569494 532454 600207
rect 531834 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 532454 569494
rect 531834 569174 532454 569258
rect 531834 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 532454 569174
rect 531834 533494 532454 568938
rect 531834 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 532454 533494
rect 531834 533174 532454 533258
rect 531834 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 532454 533174
rect 531834 497494 532454 532938
rect 531834 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 532454 497494
rect 531834 497174 532454 497258
rect 531834 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 532454 497174
rect 531834 461494 532454 496938
rect 539366 468485 539426 603603
rect 539363 468484 539429 468485
rect 539363 468420 539364 468484
rect 539428 468420 539429 468484
rect 539363 468419 539429 468420
rect 531834 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 532454 461494
rect 531834 461174 532454 461258
rect 531834 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 532454 461174
rect 531834 425494 532454 460938
rect 541022 456109 541082 618563
rect 541794 615454 542414 650898
rect 545514 705798 546134 711590
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 542675 636308 542741 636309
rect 542675 636244 542676 636308
rect 542740 636244 542741 636308
rect 542675 636243 542741 636244
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 542678 476781 542738 636243
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 542859 607748 542925 607749
rect 542859 607684 542860 607748
rect 542924 607684 542925 607748
rect 542859 607683 542925 607684
rect 542675 476780 542741 476781
rect 542675 476716 542676 476780
rect 542740 476716 542741 476780
rect 542675 476715 542741 476716
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541019 456108 541085 456109
rect 541019 456044 541020 456108
rect 541084 456044 541085 456108
rect 541019 456043 541085 456044
rect 531834 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 532454 425494
rect 531834 425174 532454 425258
rect 531834 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 532454 425174
rect 531834 389494 532454 424938
rect 531834 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 532454 389494
rect 531834 389174 532454 389258
rect 531834 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 532454 389174
rect 531834 353494 532454 388938
rect 531834 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 532454 353494
rect 531834 353174 532454 353258
rect 531834 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 532454 353174
rect 531834 317494 532454 352938
rect 531834 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 532454 317494
rect 531834 317174 532454 317258
rect 531834 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 532454 317174
rect 531834 281494 532454 316938
rect 531834 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 532454 281494
rect 531834 281174 532454 281258
rect 531834 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 532454 281174
rect 531834 245494 532454 280938
rect 531834 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 532454 245494
rect 531834 245174 532454 245258
rect 531834 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 532454 245174
rect 531834 209494 532454 244938
rect 531834 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 532454 209494
rect 531834 209174 532454 209258
rect 531834 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 532454 209174
rect 531834 173494 532454 208938
rect 531834 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 532454 173494
rect 531834 173174 532454 173258
rect 531834 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 532454 173174
rect 531834 137494 532454 172938
rect 531834 137258 531866 137494
rect 532102 137258 532186 137494
rect 532422 137258 532454 137494
rect 531834 137174 532454 137258
rect 531834 136938 531866 137174
rect 532102 136938 532186 137174
rect 532422 136938 532454 137174
rect 531834 101494 532454 136938
rect 531834 101258 531866 101494
rect 532102 101258 532186 101494
rect 532422 101258 532454 101494
rect 531834 101174 532454 101258
rect 531834 100938 531866 101174
rect 532102 100938 532186 101174
rect 532422 100938 532454 101174
rect 531834 65494 532454 100938
rect 531834 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 532454 65494
rect 531834 65174 532454 65258
rect 531834 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 532454 65174
rect 531834 29494 532454 64938
rect 531834 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 532454 29494
rect 531834 29174 532454 29258
rect 531834 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 532454 29174
rect 531834 -7066 532454 28938
rect 531834 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 532454 -7066
rect 531834 -7386 532454 -7302
rect 531834 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 532454 -7386
rect 531834 -7654 532454 -7622
rect 541794 435454 542414 470898
rect 542862 450533 542922 607683
rect 543043 606388 543109 606389
rect 543043 606324 543044 606388
rect 543108 606324 543109 606388
rect 543043 606323 543109 606324
rect 543046 474061 543106 606323
rect 543227 605028 543293 605029
rect 543227 604964 543228 605028
rect 543292 604964 543293 605028
rect 543227 604963 543293 604964
rect 543230 479501 543290 604963
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 543227 479500 543293 479501
rect 543227 479436 543228 479500
rect 543292 479436 543293 479500
rect 543227 479435 543293 479436
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 543043 474060 543109 474061
rect 543043 473996 543044 474060
rect 543108 473996 543109 474060
rect 543043 473995 543109 473996
rect 542859 450532 542925 450533
rect 542859 450468 542860 450532
rect 542924 450468 542925 450532
rect 542859 450467 542925 450468
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 544331 312084 544397 312085
rect 544331 312020 544332 312084
rect 544396 312020 544397 312084
rect 544331 312019 544397 312020
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 544334 250749 544394 312019
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 544331 250748 544397 250749
rect 544331 250684 544332 250748
rect 544396 250684 544397 250748
rect 544331 250683 544397 250684
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -7654 546134 -1862
rect 549234 706758 549854 711590
rect 549234 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 549854 706758
rect 549234 706438 549854 706522
rect 549234 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 549854 706438
rect 549234 694894 549854 706202
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -2266 549854 10338
rect 549234 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 549854 -2266
rect 549234 -2586 549854 -2502
rect 549234 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 549854 -2586
rect 549234 -7654 549854 -2822
rect 552954 707718 553574 711590
rect 552954 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 553574 707718
rect 552954 707398 553574 707482
rect 552954 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 553574 707398
rect 552954 698614 553574 707162
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 552954 -3226 553574 14058
rect 552954 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 553574 -3226
rect 552954 -3546 553574 -3462
rect 552954 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 553574 -3546
rect 552954 -7654 553574 -3782
rect 556674 708678 557294 711590
rect 556674 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 557294 708678
rect 556674 708358 557294 708442
rect 556674 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 557294 708358
rect 556674 666334 557294 708122
rect 556674 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 557294 666334
rect 556674 666014 557294 666098
rect 556674 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 557294 666014
rect 556674 630334 557294 665778
rect 556674 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 557294 630334
rect 556674 630014 557294 630098
rect 556674 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 557294 630014
rect 556674 594334 557294 629778
rect 556674 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 557294 594334
rect 556674 594014 557294 594098
rect 556674 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 557294 594014
rect 556674 558334 557294 593778
rect 556674 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 557294 558334
rect 556674 558014 557294 558098
rect 556674 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 557294 558014
rect 556674 522334 557294 557778
rect 556674 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 557294 522334
rect 556674 522014 557294 522098
rect 556674 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 557294 522014
rect 556674 486334 557294 521778
rect 556674 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 557294 486334
rect 556674 486014 557294 486098
rect 556674 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 557294 486014
rect 556674 450334 557294 485778
rect 556674 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 557294 450334
rect 556674 450014 557294 450098
rect 556674 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 557294 450014
rect 556674 414334 557294 449778
rect 556674 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 557294 414334
rect 556674 414014 557294 414098
rect 556674 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 557294 414014
rect 556674 378334 557294 413778
rect 556674 378098 556706 378334
rect 556942 378098 557026 378334
rect 557262 378098 557294 378334
rect 556674 378014 557294 378098
rect 556674 377778 556706 378014
rect 556942 377778 557026 378014
rect 557262 377778 557294 378014
rect 556674 342334 557294 377778
rect 556674 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 557294 342334
rect 556674 342014 557294 342098
rect 556674 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 557294 342014
rect 556674 306334 557294 341778
rect 556674 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 557294 306334
rect 556674 306014 557294 306098
rect 556674 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 557294 306014
rect 556674 270334 557294 305778
rect 556674 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 557294 270334
rect 556674 270014 557294 270098
rect 556674 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 557294 270014
rect 556674 234334 557294 269778
rect 560394 709638 561014 711590
rect 560394 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 561014 709638
rect 560394 709318 561014 709402
rect 560394 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 561014 709318
rect 560394 670054 561014 709082
rect 560394 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 561014 670054
rect 560394 669734 561014 669818
rect 560394 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 561014 669734
rect 560394 634054 561014 669498
rect 560394 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 561014 634054
rect 560394 633734 561014 633818
rect 560394 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 561014 633734
rect 560394 598054 561014 633498
rect 560394 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 561014 598054
rect 560394 597734 561014 597818
rect 560394 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 561014 597734
rect 560394 562054 561014 597498
rect 560394 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 561014 562054
rect 560394 561734 561014 561818
rect 560394 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 561014 561734
rect 560394 526054 561014 561498
rect 560394 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 561014 526054
rect 560394 525734 561014 525818
rect 560394 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 561014 525734
rect 560394 490054 561014 525498
rect 560394 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 561014 490054
rect 560394 489734 561014 489818
rect 560394 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 561014 489734
rect 560394 454054 561014 489498
rect 560394 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 561014 454054
rect 560394 453734 561014 453818
rect 560394 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 561014 453734
rect 560394 418054 561014 453498
rect 560394 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 561014 418054
rect 560394 417734 561014 417818
rect 560394 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 561014 417734
rect 560394 382054 561014 417498
rect 560394 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 561014 382054
rect 560394 381734 561014 381818
rect 560394 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 561014 381734
rect 560394 346054 561014 381498
rect 560394 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 561014 346054
rect 560394 345734 561014 345818
rect 560394 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 561014 345734
rect 560394 310054 561014 345498
rect 560394 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 561014 310054
rect 560394 309734 561014 309818
rect 560394 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 561014 309734
rect 560394 274054 561014 309498
rect 560394 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 561014 274054
rect 560394 273734 561014 273818
rect 560394 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 561014 273734
rect 559419 242588 559485 242589
rect 559419 242524 559420 242588
rect 559484 242524 559485 242588
rect 559419 242523 559485 242524
rect 556674 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 557294 234334
rect 556674 234014 557294 234098
rect 556674 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 557294 234014
rect 556674 198334 557294 233778
rect 556674 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 557294 198334
rect 556674 198014 557294 198098
rect 556674 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 557294 198014
rect 556674 162334 557294 197778
rect 556674 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 557294 162334
rect 556674 162014 557294 162098
rect 556674 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 557294 162014
rect 556674 126334 557294 161778
rect 556674 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 557294 126334
rect 556674 126014 557294 126098
rect 556674 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 557294 126014
rect 556674 90334 557294 125778
rect 556674 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 557294 90334
rect 556674 90014 557294 90098
rect 556674 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 557294 90014
rect 556674 54334 557294 89778
rect 559422 59669 559482 242523
rect 560394 238054 561014 273498
rect 560394 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 561014 238054
rect 560394 237734 561014 237818
rect 560394 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 561014 237734
rect 560394 202054 561014 237498
rect 560394 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 561014 202054
rect 560394 201734 561014 201818
rect 560394 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 561014 201734
rect 560394 166054 561014 201498
rect 560394 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 561014 166054
rect 560394 165734 561014 165818
rect 560394 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 561014 165734
rect 560394 130054 561014 165498
rect 560394 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 561014 130054
rect 560394 129734 561014 129818
rect 560394 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 561014 129734
rect 560394 94054 561014 129498
rect 560394 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 561014 94054
rect 560394 93734 561014 93818
rect 560394 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 561014 93734
rect 559419 59668 559485 59669
rect 559419 59604 559420 59668
rect 559484 59604 559485 59668
rect 559419 59603 559485 59604
rect 556674 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 557294 54334
rect 556674 54014 557294 54098
rect 556674 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 557294 54014
rect 556674 18334 557294 53778
rect 556674 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 557294 18334
rect 556674 18014 557294 18098
rect 556674 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 557294 18014
rect 556674 -4186 557294 17778
rect 556674 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 557294 -4186
rect 556674 -4506 557294 -4422
rect 556674 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 557294 -4506
rect 556674 -7654 557294 -4742
rect 560394 58054 561014 93498
rect 560394 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 561014 58054
rect 560394 57734 561014 57818
rect 560394 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 561014 57734
rect 560394 22054 561014 57498
rect 560394 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 561014 22054
rect 560394 21734 561014 21818
rect 560394 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 561014 21734
rect 560394 -5146 561014 21498
rect 560394 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 561014 -5146
rect 560394 -5466 561014 -5382
rect 560394 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 561014 -5466
rect 560394 -7654 561014 -5702
rect 564114 710598 564734 711590
rect 564114 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 564734 710598
rect 564114 710278 564734 710362
rect 564114 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 564734 710278
rect 564114 673774 564734 710042
rect 564114 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 564734 673774
rect 564114 673454 564734 673538
rect 564114 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 564734 673454
rect 564114 637774 564734 673218
rect 564114 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 564734 637774
rect 564114 637454 564734 637538
rect 564114 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 564734 637454
rect 564114 601774 564734 637218
rect 564114 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 564734 601774
rect 564114 601454 564734 601538
rect 564114 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 564734 601454
rect 564114 565774 564734 601218
rect 564114 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 564734 565774
rect 564114 565454 564734 565538
rect 564114 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 564734 565454
rect 564114 529774 564734 565218
rect 564114 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 564734 529774
rect 564114 529454 564734 529538
rect 564114 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 564734 529454
rect 564114 493774 564734 529218
rect 564114 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 564734 493774
rect 564114 493454 564734 493538
rect 564114 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 564734 493454
rect 564114 457774 564734 493218
rect 564114 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 564734 457774
rect 564114 457454 564734 457538
rect 564114 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 564734 457454
rect 564114 421774 564734 457218
rect 564114 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 564734 421774
rect 564114 421454 564734 421538
rect 564114 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 564734 421454
rect 564114 385774 564734 421218
rect 564114 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 564734 385774
rect 564114 385454 564734 385538
rect 564114 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 564734 385454
rect 564114 349774 564734 385218
rect 564114 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 564734 349774
rect 564114 349454 564734 349538
rect 564114 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 564734 349454
rect 564114 313774 564734 349218
rect 564114 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 564734 313774
rect 564114 313454 564734 313538
rect 564114 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 564734 313454
rect 564114 277774 564734 313218
rect 564114 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 564734 277774
rect 564114 277454 564734 277538
rect 564114 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 564734 277454
rect 564114 241774 564734 277218
rect 564114 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 564734 241774
rect 564114 241454 564734 241538
rect 564114 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 564734 241454
rect 564114 205774 564734 241218
rect 564114 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 564734 205774
rect 564114 205454 564734 205538
rect 564114 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 564734 205454
rect 564114 169774 564734 205218
rect 564114 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 564734 169774
rect 564114 169454 564734 169538
rect 564114 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 564734 169454
rect 564114 133774 564734 169218
rect 564114 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 564734 133774
rect 564114 133454 564734 133538
rect 564114 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 564734 133454
rect 564114 97774 564734 133218
rect 564114 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 564734 97774
rect 564114 97454 564734 97538
rect 564114 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 564734 97454
rect 564114 61774 564734 97218
rect 564114 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 564734 61774
rect 564114 61454 564734 61538
rect 564114 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 564734 61454
rect 564114 25774 564734 61218
rect 564114 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 564734 25774
rect 564114 25454 564734 25538
rect 564114 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 564734 25454
rect 564114 -6106 564734 25218
rect 564114 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 564734 -6106
rect 564114 -6426 564734 -6342
rect 564114 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 564734 -6426
rect 564114 -7654 564734 -6662
rect 567834 711558 568454 711590
rect 567834 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 568454 711558
rect 567834 711238 568454 711322
rect 567834 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 568454 711238
rect 567834 677494 568454 711002
rect 567834 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 568454 677494
rect 567834 677174 568454 677258
rect 567834 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 568454 677174
rect 567834 641494 568454 676938
rect 567834 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 568454 641494
rect 567834 641174 568454 641258
rect 567834 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 568454 641174
rect 567834 605494 568454 640938
rect 567834 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 568454 605494
rect 567834 605174 568454 605258
rect 567834 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 568454 605174
rect 567834 569494 568454 604938
rect 567834 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 568454 569494
rect 567834 569174 568454 569258
rect 567834 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 568454 569174
rect 567834 533494 568454 568938
rect 567834 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 568454 533494
rect 567834 533174 568454 533258
rect 567834 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 568454 533174
rect 567834 497494 568454 532938
rect 567834 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 568454 497494
rect 567834 497174 568454 497258
rect 567834 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 568454 497174
rect 567834 461494 568454 496938
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 580211 630868 580277 630869
rect 580211 630804 580212 630868
rect 580276 630804 580277 630868
rect 580211 630803 580277 630804
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 580214 591293 580274 630803
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 580211 591292 580277 591293
rect 580211 591228 580212 591292
rect 580276 591228 580277 591292
rect 580211 591227 580277 591228
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 574691 471476 574757 471477
rect 574691 471412 574692 471476
rect 574756 471412 574757 471476
rect 574691 471411 574757 471412
rect 577794 471454 578414 506898
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 580211 484668 580277 484669
rect 580211 484604 580212 484668
rect 580276 484604 580277 484668
rect 580211 484603 580277 484604
rect 580214 478141 580274 484603
rect 580211 478140 580277 478141
rect 580211 478076 580212 478140
rect 580276 478076 580277 478140
rect 580211 478075 580277 478076
rect 567834 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 568454 461494
rect 567834 461174 568454 461258
rect 567834 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 568454 461174
rect 567834 425494 568454 460938
rect 567834 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 568454 425494
rect 567834 425174 568454 425258
rect 567834 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 568454 425174
rect 567834 389494 568454 424938
rect 567834 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 568454 389494
rect 567834 389174 568454 389258
rect 567834 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 568454 389174
rect 567834 353494 568454 388938
rect 567834 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 568454 353494
rect 567834 353174 568454 353258
rect 567834 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 568454 353174
rect 567834 317494 568454 352938
rect 567834 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 568454 317494
rect 567834 317174 568454 317258
rect 567834 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 568454 317174
rect 567834 281494 568454 316938
rect 567834 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 568454 281494
rect 567834 281174 568454 281258
rect 567834 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 568454 281174
rect 567834 245494 568454 280938
rect 574694 254829 574754 471411
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 580211 365124 580277 365125
rect 580211 365060 580212 365124
rect 580276 365060 580277 365124
rect 580211 365059 580277 365060
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 580214 329085 580274 365059
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 580211 329084 580277 329085
rect 580211 329020 580212 329084
rect 580276 329020 580277 329084
rect 580211 329019 580277 329020
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 580211 325276 580277 325277
rect 580211 325212 580212 325276
rect 580276 325212 580277 325276
rect 580211 325211 580277 325212
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 574691 254828 574757 254829
rect 574691 254764 574692 254828
rect 574756 254764 574757 254828
rect 574691 254763 574757 254764
rect 567834 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 568454 245494
rect 567834 245174 568454 245258
rect 567834 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 568454 245174
rect 567834 209494 568454 244938
rect 567834 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 568454 209494
rect 567834 209174 568454 209258
rect 567834 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 568454 209174
rect 567834 173494 568454 208938
rect 567834 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 568454 173494
rect 567834 173174 568454 173258
rect 567834 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 568454 173174
rect 567834 137494 568454 172938
rect 567834 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 568454 137494
rect 567834 137174 568454 137258
rect 567834 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 568454 137174
rect 567834 101494 568454 136938
rect 567834 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 568454 101494
rect 567834 101174 568454 101258
rect 567834 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 568454 101174
rect 567834 65494 568454 100938
rect 567834 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 568454 65494
rect 567834 65174 568454 65258
rect 567834 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 568454 65174
rect 567834 29494 568454 64938
rect 567834 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 568454 29494
rect 567834 29174 568454 29258
rect 567834 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 568454 29174
rect 567834 -7066 568454 28938
rect 567834 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 568454 -7066
rect 567834 -7386 568454 -7302
rect 567834 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 568454 -7386
rect 567834 -7654 568454 -7622
rect 577794 219454 578414 254898
rect 580214 240005 580274 325211
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 580395 272236 580461 272237
rect 580395 272172 580396 272236
rect 580460 272172 580461 272236
rect 580395 272171 580461 272172
rect 580211 240004 580277 240005
rect 580211 239940 580212 240004
rect 580276 239940 580277 240004
rect 580211 239939 580277 239940
rect 580398 239053 580458 272171
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 580395 239052 580461 239053
rect 580395 238988 580396 239052
rect 580460 238988 580461 239052
rect 580395 238987 580461 238988
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 587850 694894
rect 587230 694574 587850 694658
rect 587230 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 587850 694574
rect 587230 658894 587850 694338
rect 587230 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 587850 658894
rect 587230 658574 587850 658658
rect 587230 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 587850 658574
rect 587230 622894 587850 658338
rect 587230 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 587850 622894
rect 587230 622574 587850 622658
rect 587230 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 587850 622574
rect 587230 586894 587850 622338
rect 587230 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 587850 586894
rect 587230 586574 587850 586658
rect 587230 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 587850 586574
rect 587230 550894 587850 586338
rect 587230 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 587850 550894
rect 587230 550574 587850 550658
rect 587230 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 587850 550574
rect 587230 514894 587850 550338
rect 587230 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 587850 514894
rect 587230 514574 587850 514658
rect 587230 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 587850 514574
rect 587230 478894 587850 514338
rect 587230 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 587850 478894
rect 587230 478574 587850 478658
rect 587230 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 587850 478574
rect 587230 442894 587850 478338
rect 587230 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 587850 442894
rect 587230 442574 587850 442658
rect 587230 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 587850 442574
rect 587230 406894 587850 442338
rect 587230 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 587850 406894
rect 587230 406574 587850 406658
rect 587230 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 587850 406574
rect 587230 370894 587850 406338
rect 587230 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 587850 370894
rect 587230 370574 587850 370658
rect 587230 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 587850 370574
rect 587230 334894 587850 370338
rect 587230 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 587850 334894
rect 587230 334574 587850 334658
rect 587230 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 587850 334574
rect 587230 298894 587850 334338
rect 587230 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 587850 298894
rect 587230 298574 587850 298658
rect 587230 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 587850 298574
rect 587230 262894 587850 298338
rect 587230 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 587850 262894
rect 587230 262574 587850 262658
rect 587230 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 587850 262574
rect 587230 226894 587850 262338
rect 587230 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 587850 226894
rect 587230 226574 587850 226658
rect 587230 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 587850 226574
rect 587230 190894 587850 226338
rect 587230 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 587850 190894
rect 587230 190574 587850 190658
rect 587230 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 587850 190574
rect 587230 154894 587850 190338
rect 587230 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 587850 154894
rect 587230 154574 587850 154658
rect 587230 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 587850 154574
rect 587230 118894 587850 154338
rect 587230 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 587850 118894
rect 587230 118574 587850 118658
rect 587230 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 587850 118574
rect 587230 82894 587850 118338
rect 587230 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 587850 82894
rect 587230 82574 587850 82658
rect 587230 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 587850 82574
rect 587230 46894 587850 82338
rect 587230 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 587850 46894
rect 587230 46574 587850 46658
rect 587230 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 587850 46574
rect 587230 10894 587850 46338
rect 587230 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 587850 10894
rect 587230 10574 587850 10658
rect 587230 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 587850 10574
rect 587230 -2266 587850 10338
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 588810 698614
rect 588190 698294 588810 698378
rect 588190 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 588810 698294
rect 588190 662614 588810 698058
rect 588190 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 588810 662614
rect 588190 662294 588810 662378
rect 588190 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 588810 662294
rect 588190 626614 588810 662058
rect 588190 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 588810 626614
rect 588190 626294 588810 626378
rect 588190 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 588810 626294
rect 588190 590614 588810 626058
rect 588190 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 588810 590614
rect 588190 590294 588810 590378
rect 588190 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 588810 590294
rect 588190 554614 588810 590058
rect 588190 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 588810 554614
rect 588190 554294 588810 554378
rect 588190 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 588810 554294
rect 588190 518614 588810 554058
rect 588190 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 588810 518614
rect 588190 518294 588810 518378
rect 588190 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 588810 518294
rect 588190 482614 588810 518058
rect 588190 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 588810 482614
rect 588190 482294 588810 482378
rect 588190 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 588810 482294
rect 588190 446614 588810 482058
rect 588190 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 588810 446614
rect 588190 446294 588810 446378
rect 588190 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 588810 446294
rect 588190 410614 588810 446058
rect 588190 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 588810 410614
rect 588190 410294 588810 410378
rect 588190 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 588810 410294
rect 588190 374614 588810 410058
rect 588190 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 588810 374614
rect 588190 374294 588810 374378
rect 588190 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 588810 374294
rect 588190 338614 588810 374058
rect 588190 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 588810 338614
rect 588190 338294 588810 338378
rect 588190 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 588810 338294
rect 588190 302614 588810 338058
rect 588190 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 588810 302614
rect 588190 302294 588810 302378
rect 588190 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 588810 302294
rect 588190 266614 588810 302058
rect 588190 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 588810 266614
rect 588190 266294 588810 266378
rect 588190 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 588810 266294
rect 588190 230614 588810 266058
rect 588190 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 588810 230614
rect 588190 230294 588810 230378
rect 588190 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 588810 230294
rect 588190 194614 588810 230058
rect 588190 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 588810 194614
rect 588190 194294 588810 194378
rect 588190 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 588810 194294
rect 588190 158614 588810 194058
rect 588190 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 588810 158614
rect 588190 158294 588810 158378
rect 588190 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 588810 158294
rect 588190 122614 588810 158058
rect 588190 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 588810 122614
rect 588190 122294 588810 122378
rect 588190 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 588810 122294
rect 588190 86614 588810 122058
rect 588190 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 588810 86614
rect 588190 86294 588810 86378
rect 588190 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 588810 86294
rect 588190 50614 588810 86058
rect 588190 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 588810 50614
rect 588190 50294 588810 50378
rect 588190 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 588810 50294
rect 588190 14614 588810 50058
rect 588190 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 588810 14614
rect 588190 14294 588810 14378
rect 588190 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 588810 14294
rect 588190 -3226 588810 14058
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 589770 666334
rect 589150 666014 589770 666098
rect 589150 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 589770 666014
rect 589150 630334 589770 665778
rect 589150 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 589770 630334
rect 589150 630014 589770 630098
rect 589150 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 589770 630014
rect 589150 594334 589770 629778
rect 589150 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 589770 594334
rect 589150 594014 589770 594098
rect 589150 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 589770 594014
rect 589150 558334 589770 593778
rect 589150 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 589770 558334
rect 589150 558014 589770 558098
rect 589150 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 589770 558014
rect 589150 522334 589770 557778
rect 589150 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 589770 522334
rect 589150 522014 589770 522098
rect 589150 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 589770 522014
rect 589150 486334 589770 521778
rect 589150 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 589770 486334
rect 589150 486014 589770 486098
rect 589150 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 589770 486014
rect 589150 450334 589770 485778
rect 589150 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 589770 450334
rect 589150 450014 589770 450098
rect 589150 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 589770 450014
rect 589150 414334 589770 449778
rect 589150 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 589770 414334
rect 589150 414014 589770 414098
rect 589150 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 589770 414014
rect 589150 378334 589770 413778
rect 589150 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 589770 378334
rect 589150 378014 589770 378098
rect 589150 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 589770 378014
rect 589150 342334 589770 377778
rect 589150 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 589770 342334
rect 589150 342014 589770 342098
rect 589150 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 589770 342014
rect 589150 306334 589770 341778
rect 589150 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 589770 306334
rect 589150 306014 589770 306098
rect 589150 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 589770 306014
rect 589150 270334 589770 305778
rect 589150 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 589770 270334
rect 589150 270014 589770 270098
rect 589150 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 589770 270014
rect 589150 234334 589770 269778
rect 589150 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 589770 234334
rect 589150 234014 589770 234098
rect 589150 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 589770 234014
rect 589150 198334 589770 233778
rect 589150 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 589770 198334
rect 589150 198014 589770 198098
rect 589150 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 589770 198014
rect 589150 162334 589770 197778
rect 589150 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 589770 162334
rect 589150 162014 589770 162098
rect 589150 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 589770 162014
rect 589150 126334 589770 161778
rect 589150 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 589770 126334
rect 589150 126014 589770 126098
rect 589150 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 589770 126014
rect 589150 90334 589770 125778
rect 589150 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 589770 90334
rect 589150 90014 589770 90098
rect 589150 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 589770 90014
rect 589150 54334 589770 89778
rect 589150 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 589770 54334
rect 589150 54014 589770 54098
rect 589150 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 589770 54014
rect 589150 18334 589770 53778
rect 589150 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 589770 18334
rect 589150 18014 589770 18098
rect 589150 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 589770 18014
rect 589150 -4186 589770 17778
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 590730 670054
rect 590110 669734 590730 669818
rect 590110 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 590730 669734
rect 590110 634054 590730 669498
rect 590110 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 590730 634054
rect 590110 633734 590730 633818
rect 590110 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 590730 633734
rect 590110 598054 590730 633498
rect 590110 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 590730 598054
rect 590110 597734 590730 597818
rect 590110 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 590730 597734
rect 590110 562054 590730 597498
rect 590110 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 590730 562054
rect 590110 561734 590730 561818
rect 590110 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 590730 561734
rect 590110 526054 590730 561498
rect 590110 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 590730 526054
rect 590110 525734 590730 525818
rect 590110 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 590730 525734
rect 590110 490054 590730 525498
rect 590110 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 590730 490054
rect 590110 489734 590730 489818
rect 590110 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 590730 489734
rect 590110 454054 590730 489498
rect 590110 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 590730 454054
rect 590110 453734 590730 453818
rect 590110 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 590730 453734
rect 590110 418054 590730 453498
rect 590110 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 590730 418054
rect 590110 417734 590730 417818
rect 590110 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 590730 417734
rect 590110 382054 590730 417498
rect 590110 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 590730 382054
rect 590110 381734 590730 381818
rect 590110 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 590730 381734
rect 590110 346054 590730 381498
rect 590110 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 590730 346054
rect 590110 345734 590730 345818
rect 590110 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 590730 345734
rect 590110 310054 590730 345498
rect 590110 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 590730 310054
rect 590110 309734 590730 309818
rect 590110 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 590730 309734
rect 590110 274054 590730 309498
rect 590110 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 590730 274054
rect 590110 273734 590730 273818
rect 590110 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 590730 273734
rect 590110 238054 590730 273498
rect 590110 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 590730 238054
rect 590110 237734 590730 237818
rect 590110 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 590730 237734
rect 590110 202054 590730 237498
rect 590110 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 590730 202054
rect 590110 201734 590730 201818
rect 590110 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 590730 201734
rect 590110 166054 590730 201498
rect 590110 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 590730 166054
rect 590110 165734 590730 165818
rect 590110 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 590730 165734
rect 590110 130054 590730 165498
rect 590110 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 590730 130054
rect 590110 129734 590730 129818
rect 590110 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 590730 129734
rect 590110 94054 590730 129498
rect 590110 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 590730 94054
rect 590110 93734 590730 93818
rect 590110 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 590730 93734
rect 590110 58054 590730 93498
rect 590110 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 590730 58054
rect 590110 57734 590730 57818
rect 590110 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 590730 57734
rect 590110 22054 590730 57498
rect 590110 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 590730 22054
rect 590110 21734 590730 21818
rect 590110 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 590730 21734
rect 590110 -5146 590730 21498
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 591690 673774
rect 591070 673454 591690 673538
rect 591070 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 591690 673454
rect 591070 637774 591690 673218
rect 591070 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 591690 637774
rect 591070 637454 591690 637538
rect 591070 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 591690 637454
rect 591070 601774 591690 637218
rect 591070 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 591690 601774
rect 591070 601454 591690 601538
rect 591070 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 591690 601454
rect 591070 565774 591690 601218
rect 591070 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 591690 565774
rect 591070 565454 591690 565538
rect 591070 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 591690 565454
rect 591070 529774 591690 565218
rect 591070 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 591690 529774
rect 591070 529454 591690 529538
rect 591070 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 591690 529454
rect 591070 493774 591690 529218
rect 591070 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 591690 493774
rect 591070 493454 591690 493538
rect 591070 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 591690 493454
rect 591070 457774 591690 493218
rect 591070 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 591690 457774
rect 591070 457454 591690 457538
rect 591070 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 591690 457454
rect 591070 421774 591690 457218
rect 591070 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 591690 421774
rect 591070 421454 591690 421538
rect 591070 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 591690 421454
rect 591070 385774 591690 421218
rect 591070 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 591690 385774
rect 591070 385454 591690 385538
rect 591070 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 591690 385454
rect 591070 349774 591690 385218
rect 591070 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 591690 349774
rect 591070 349454 591690 349538
rect 591070 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 591690 349454
rect 591070 313774 591690 349218
rect 591070 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 591690 313774
rect 591070 313454 591690 313538
rect 591070 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 591690 313454
rect 591070 277774 591690 313218
rect 591070 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 591690 277774
rect 591070 277454 591690 277538
rect 591070 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 591690 277454
rect 591070 241774 591690 277218
rect 591070 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 591690 241774
rect 591070 241454 591690 241538
rect 591070 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 591690 241454
rect 591070 205774 591690 241218
rect 591070 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 591690 205774
rect 591070 205454 591690 205538
rect 591070 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 591690 205454
rect 591070 169774 591690 205218
rect 591070 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 591690 169774
rect 591070 169454 591690 169538
rect 591070 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 591690 169454
rect 591070 133774 591690 169218
rect 591070 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 591690 133774
rect 591070 133454 591690 133538
rect 591070 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 591690 133454
rect 591070 97774 591690 133218
rect 591070 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 591690 97774
rect 591070 97454 591690 97538
rect 591070 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 591690 97454
rect 591070 61774 591690 97218
rect 591070 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 591690 61774
rect 591070 61454 591690 61538
rect 591070 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 591690 61454
rect 591070 25774 591690 61218
rect 591070 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 591690 25774
rect 591070 25454 591690 25538
rect 591070 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 591690 25454
rect 591070 -6106 591690 25218
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect 592030 677174 592650 677258
rect 592030 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect 592030 641494 592650 676938
rect 592030 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect 592030 641174 592650 641258
rect 592030 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect 592030 605494 592650 640938
rect 592030 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect 592030 605174 592650 605258
rect 592030 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect 592030 569494 592650 604938
rect 592030 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect 592030 569174 592650 569258
rect 592030 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect 592030 533494 592650 568938
rect 592030 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect 592030 533174 592650 533258
rect 592030 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect 592030 497494 592650 532938
rect 592030 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect 592030 497174 592650 497258
rect 592030 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect 592030 461494 592650 496938
rect 592030 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect 592030 461174 592650 461258
rect 592030 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect 592030 425494 592650 460938
rect 592030 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect 592030 425174 592650 425258
rect 592030 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect 592030 389494 592650 424938
rect 592030 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect 592030 389174 592650 389258
rect 592030 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect 592030 353494 592650 388938
rect 592030 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect 592030 353174 592650 353258
rect 592030 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect 592030 317494 592650 352938
rect 592030 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect 592030 317174 592650 317258
rect 592030 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect 592030 281494 592650 316938
rect 592030 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect 592030 281174 592650 281258
rect 592030 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect 592030 245494 592650 280938
rect 592030 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect 592030 245174 592650 245258
rect 592030 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect 592030 209494 592650 244938
rect 592030 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect 592030 209174 592650 209258
rect 592030 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect 592030 173494 592650 208938
rect 592030 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect 592030 173174 592650 173258
rect 592030 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect 592030 137494 592650 172938
rect 592030 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect 592030 137174 592650 137258
rect 592030 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect 592030 101494 592650 136938
rect 592030 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect 592030 101174 592650 101258
rect 592030 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect 592030 65494 592650 100938
rect 592030 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect 592030 65174 592650 65258
rect 592030 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect 592030 29494 592650 64938
rect 592030 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect 592030 29174 592650 29258
rect 592030 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect 592030 -7066 592650 28938
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 677258 -8458 677494
rect -8374 677258 -8138 677494
rect -8694 676938 -8458 677174
rect -8374 676938 -8138 677174
rect -8694 641258 -8458 641494
rect -8374 641258 -8138 641494
rect -8694 640938 -8458 641174
rect -8374 640938 -8138 641174
rect -8694 605258 -8458 605494
rect -8374 605258 -8138 605494
rect -8694 604938 -8458 605174
rect -8374 604938 -8138 605174
rect -8694 569258 -8458 569494
rect -8374 569258 -8138 569494
rect -8694 568938 -8458 569174
rect -8374 568938 -8138 569174
rect -8694 533258 -8458 533494
rect -8374 533258 -8138 533494
rect -8694 532938 -8458 533174
rect -8374 532938 -8138 533174
rect -8694 497258 -8458 497494
rect -8374 497258 -8138 497494
rect -8694 496938 -8458 497174
rect -8374 496938 -8138 497174
rect -8694 461258 -8458 461494
rect -8374 461258 -8138 461494
rect -8694 460938 -8458 461174
rect -8374 460938 -8138 461174
rect -8694 425258 -8458 425494
rect -8374 425258 -8138 425494
rect -8694 424938 -8458 425174
rect -8374 424938 -8138 425174
rect -8694 389258 -8458 389494
rect -8374 389258 -8138 389494
rect -8694 388938 -8458 389174
rect -8374 388938 -8138 389174
rect -8694 353258 -8458 353494
rect -8374 353258 -8138 353494
rect -8694 352938 -8458 353174
rect -8374 352938 -8138 353174
rect -8694 317258 -8458 317494
rect -8374 317258 -8138 317494
rect -8694 316938 -8458 317174
rect -8374 316938 -8138 317174
rect -8694 281258 -8458 281494
rect -8374 281258 -8138 281494
rect -8694 280938 -8458 281174
rect -8374 280938 -8138 281174
rect -8694 245258 -8458 245494
rect -8374 245258 -8138 245494
rect -8694 244938 -8458 245174
rect -8374 244938 -8138 245174
rect -8694 209258 -8458 209494
rect -8374 209258 -8138 209494
rect -8694 208938 -8458 209174
rect -8374 208938 -8138 209174
rect -8694 173258 -8458 173494
rect -8374 173258 -8138 173494
rect -8694 172938 -8458 173174
rect -8374 172938 -8138 173174
rect -8694 137258 -8458 137494
rect -8374 137258 -8138 137494
rect -8694 136938 -8458 137174
rect -8374 136938 -8138 137174
rect -8694 101258 -8458 101494
rect -8374 101258 -8138 101494
rect -8694 100938 -8458 101174
rect -8374 100938 -8138 101174
rect -8694 65258 -8458 65494
rect -8374 65258 -8138 65494
rect -8694 64938 -8458 65174
rect -8374 64938 -8138 65174
rect -8694 29258 -8458 29494
rect -8374 29258 -8138 29494
rect -8694 28938 -8458 29174
rect -8374 28938 -8138 29174
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 673538 -7498 673774
rect -7414 673538 -7178 673774
rect -7734 673218 -7498 673454
rect -7414 673218 -7178 673454
rect -7734 637538 -7498 637774
rect -7414 637538 -7178 637774
rect -7734 637218 -7498 637454
rect -7414 637218 -7178 637454
rect -7734 601538 -7498 601774
rect -7414 601538 -7178 601774
rect -7734 601218 -7498 601454
rect -7414 601218 -7178 601454
rect -7734 565538 -7498 565774
rect -7414 565538 -7178 565774
rect -7734 565218 -7498 565454
rect -7414 565218 -7178 565454
rect -7734 529538 -7498 529774
rect -7414 529538 -7178 529774
rect -7734 529218 -7498 529454
rect -7414 529218 -7178 529454
rect -7734 493538 -7498 493774
rect -7414 493538 -7178 493774
rect -7734 493218 -7498 493454
rect -7414 493218 -7178 493454
rect -7734 457538 -7498 457774
rect -7414 457538 -7178 457774
rect -7734 457218 -7498 457454
rect -7414 457218 -7178 457454
rect -7734 421538 -7498 421774
rect -7414 421538 -7178 421774
rect -7734 421218 -7498 421454
rect -7414 421218 -7178 421454
rect -7734 385538 -7498 385774
rect -7414 385538 -7178 385774
rect -7734 385218 -7498 385454
rect -7414 385218 -7178 385454
rect -7734 349538 -7498 349774
rect -7414 349538 -7178 349774
rect -7734 349218 -7498 349454
rect -7414 349218 -7178 349454
rect -7734 313538 -7498 313774
rect -7414 313538 -7178 313774
rect -7734 313218 -7498 313454
rect -7414 313218 -7178 313454
rect -7734 277538 -7498 277774
rect -7414 277538 -7178 277774
rect -7734 277218 -7498 277454
rect -7414 277218 -7178 277454
rect -7734 241538 -7498 241774
rect -7414 241538 -7178 241774
rect -7734 241218 -7498 241454
rect -7414 241218 -7178 241454
rect -7734 205538 -7498 205774
rect -7414 205538 -7178 205774
rect -7734 205218 -7498 205454
rect -7414 205218 -7178 205454
rect -7734 169538 -7498 169774
rect -7414 169538 -7178 169774
rect -7734 169218 -7498 169454
rect -7414 169218 -7178 169454
rect -7734 133538 -7498 133774
rect -7414 133538 -7178 133774
rect -7734 133218 -7498 133454
rect -7414 133218 -7178 133454
rect -7734 97538 -7498 97774
rect -7414 97538 -7178 97774
rect -7734 97218 -7498 97454
rect -7414 97218 -7178 97454
rect -7734 61538 -7498 61774
rect -7414 61538 -7178 61774
rect -7734 61218 -7498 61454
rect -7414 61218 -7178 61454
rect -7734 25538 -7498 25774
rect -7414 25538 -7178 25774
rect -7734 25218 -7498 25454
rect -7414 25218 -7178 25454
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 669818 -6538 670054
rect -6454 669818 -6218 670054
rect -6774 669498 -6538 669734
rect -6454 669498 -6218 669734
rect -6774 633818 -6538 634054
rect -6454 633818 -6218 634054
rect -6774 633498 -6538 633734
rect -6454 633498 -6218 633734
rect -6774 597818 -6538 598054
rect -6454 597818 -6218 598054
rect -6774 597498 -6538 597734
rect -6454 597498 -6218 597734
rect -6774 561818 -6538 562054
rect -6454 561818 -6218 562054
rect -6774 561498 -6538 561734
rect -6454 561498 -6218 561734
rect -6774 525818 -6538 526054
rect -6454 525818 -6218 526054
rect -6774 525498 -6538 525734
rect -6454 525498 -6218 525734
rect -6774 489818 -6538 490054
rect -6454 489818 -6218 490054
rect -6774 489498 -6538 489734
rect -6454 489498 -6218 489734
rect -6774 453818 -6538 454054
rect -6454 453818 -6218 454054
rect -6774 453498 -6538 453734
rect -6454 453498 -6218 453734
rect -6774 417818 -6538 418054
rect -6454 417818 -6218 418054
rect -6774 417498 -6538 417734
rect -6454 417498 -6218 417734
rect -6774 381818 -6538 382054
rect -6454 381818 -6218 382054
rect -6774 381498 -6538 381734
rect -6454 381498 -6218 381734
rect -6774 345818 -6538 346054
rect -6454 345818 -6218 346054
rect -6774 345498 -6538 345734
rect -6454 345498 -6218 345734
rect -6774 309818 -6538 310054
rect -6454 309818 -6218 310054
rect -6774 309498 -6538 309734
rect -6454 309498 -6218 309734
rect -6774 273818 -6538 274054
rect -6454 273818 -6218 274054
rect -6774 273498 -6538 273734
rect -6454 273498 -6218 273734
rect -6774 237818 -6538 238054
rect -6454 237818 -6218 238054
rect -6774 237498 -6538 237734
rect -6454 237498 -6218 237734
rect -6774 201818 -6538 202054
rect -6454 201818 -6218 202054
rect -6774 201498 -6538 201734
rect -6454 201498 -6218 201734
rect -6774 165818 -6538 166054
rect -6454 165818 -6218 166054
rect -6774 165498 -6538 165734
rect -6454 165498 -6218 165734
rect -6774 129818 -6538 130054
rect -6454 129818 -6218 130054
rect -6774 129498 -6538 129734
rect -6454 129498 -6218 129734
rect -6774 93818 -6538 94054
rect -6454 93818 -6218 94054
rect -6774 93498 -6538 93734
rect -6454 93498 -6218 93734
rect -6774 57818 -6538 58054
rect -6454 57818 -6218 58054
rect -6774 57498 -6538 57734
rect -6454 57498 -6218 57734
rect -6774 21818 -6538 22054
rect -6454 21818 -6218 22054
rect -6774 21498 -6538 21734
rect -6454 21498 -6218 21734
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 666098 -5578 666334
rect -5494 666098 -5258 666334
rect -5814 665778 -5578 666014
rect -5494 665778 -5258 666014
rect -5814 630098 -5578 630334
rect -5494 630098 -5258 630334
rect -5814 629778 -5578 630014
rect -5494 629778 -5258 630014
rect -5814 594098 -5578 594334
rect -5494 594098 -5258 594334
rect -5814 593778 -5578 594014
rect -5494 593778 -5258 594014
rect -5814 558098 -5578 558334
rect -5494 558098 -5258 558334
rect -5814 557778 -5578 558014
rect -5494 557778 -5258 558014
rect -5814 522098 -5578 522334
rect -5494 522098 -5258 522334
rect -5814 521778 -5578 522014
rect -5494 521778 -5258 522014
rect -5814 486098 -5578 486334
rect -5494 486098 -5258 486334
rect -5814 485778 -5578 486014
rect -5494 485778 -5258 486014
rect -5814 450098 -5578 450334
rect -5494 450098 -5258 450334
rect -5814 449778 -5578 450014
rect -5494 449778 -5258 450014
rect -5814 414098 -5578 414334
rect -5494 414098 -5258 414334
rect -5814 413778 -5578 414014
rect -5494 413778 -5258 414014
rect -5814 378098 -5578 378334
rect -5494 378098 -5258 378334
rect -5814 377778 -5578 378014
rect -5494 377778 -5258 378014
rect -5814 342098 -5578 342334
rect -5494 342098 -5258 342334
rect -5814 341778 -5578 342014
rect -5494 341778 -5258 342014
rect -5814 306098 -5578 306334
rect -5494 306098 -5258 306334
rect -5814 305778 -5578 306014
rect -5494 305778 -5258 306014
rect -5814 270098 -5578 270334
rect -5494 270098 -5258 270334
rect -5814 269778 -5578 270014
rect -5494 269778 -5258 270014
rect -5814 234098 -5578 234334
rect -5494 234098 -5258 234334
rect -5814 233778 -5578 234014
rect -5494 233778 -5258 234014
rect -5814 198098 -5578 198334
rect -5494 198098 -5258 198334
rect -5814 197778 -5578 198014
rect -5494 197778 -5258 198014
rect -5814 162098 -5578 162334
rect -5494 162098 -5258 162334
rect -5814 161778 -5578 162014
rect -5494 161778 -5258 162014
rect -5814 126098 -5578 126334
rect -5494 126098 -5258 126334
rect -5814 125778 -5578 126014
rect -5494 125778 -5258 126014
rect -5814 90098 -5578 90334
rect -5494 90098 -5258 90334
rect -5814 89778 -5578 90014
rect -5494 89778 -5258 90014
rect -5814 54098 -5578 54334
rect -5494 54098 -5258 54334
rect -5814 53778 -5578 54014
rect -5494 53778 -5258 54014
rect -5814 18098 -5578 18334
rect -5494 18098 -5258 18334
rect -5814 17778 -5578 18014
rect -5494 17778 -5258 18014
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 698378 -4618 698614
rect -4534 698378 -4298 698614
rect -4854 698058 -4618 698294
rect -4534 698058 -4298 698294
rect -4854 662378 -4618 662614
rect -4534 662378 -4298 662614
rect -4854 662058 -4618 662294
rect -4534 662058 -4298 662294
rect -4854 626378 -4618 626614
rect -4534 626378 -4298 626614
rect -4854 626058 -4618 626294
rect -4534 626058 -4298 626294
rect -4854 590378 -4618 590614
rect -4534 590378 -4298 590614
rect -4854 590058 -4618 590294
rect -4534 590058 -4298 590294
rect -4854 554378 -4618 554614
rect -4534 554378 -4298 554614
rect -4854 554058 -4618 554294
rect -4534 554058 -4298 554294
rect -4854 518378 -4618 518614
rect -4534 518378 -4298 518614
rect -4854 518058 -4618 518294
rect -4534 518058 -4298 518294
rect -4854 482378 -4618 482614
rect -4534 482378 -4298 482614
rect -4854 482058 -4618 482294
rect -4534 482058 -4298 482294
rect -4854 446378 -4618 446614
rect -4534 446378 -4298 446614
rect -4854 446058 -4618 446294
rect -4534 446058 -4298 446294
rect -4854 410378 -4618 410614
rect -4534 410378 -4298 410614
rect -4854 410058 -4618 410294
rect -4534 410058 -4298 410294
rect -4854 374378 -4618 374614
rect -4534 374378 -4298 374614
rect -4854 374058 -4618 374294
rect -4534 374058 -4298 374294
rect -4854 338378 -4618 338614
rect -4534 338378 -4298 338614
rect -4854 338058 -4618 338294
rect -4534 338058 -4298 338294
rect -4854 302378 -4618 302614
rect -4534 302378 -4298 302614
rect -4854 302058 -4618 302294
rect -4534 302058 -4298 302294
rect -4854 266378 -4618 266614
rect -4534 266378 -4298 266614
rect -4854 266058 -4618 266294
rect -4534 266058 -4298 266294
rect -4854 230378 -4618 230614
rect -4534 230378 -4298 230614
rect -4854 230058 -4618 230294
rect -4534 230058 -4298 230294
rect -4854 194378 -4618 194614
rect -4534 194378 -4298 194614
rect -4854 194058 -4618 194294
rect -4534 194058 -4298 194294
rect -4854 158378 -4618 158614
rect -4534 158378 -4298 158614
rect -4854 158058 -4618 158294
rect -4534 158058 -4298 158294
rect -4854 122378 -4618 122614
rect -4534 122378 -4298 122614
rect -4854 122058 -4618 122294
rect -4534 122058 -4298 122294
rect -4854 86378 -4618 86614
rect -4534 86378 -4298 86614
rect -4854 86058 -4618 86294
rect -4534 86058 -4298 86294
rect -4854 50378 -4618 50614
rect -4534 50378 -4298 50614
rect -4854 50058 -4618 50294
rect -4534 50058 -4298 50294
rect -4854 14378 -4618 14614
rect -4534 14378 -4298 14614
rect -4854 14058 -4618 14294
rect -4534 14058 -4298 14294
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 694658 -3658 694894
rect -3574 694658 -3338 694894
rect -3894 694338 -3658 694574
rect -3574 694338 -3338 694574
rect -3894 658658 -3658 658894
rect -3574 658658 -3338 658894
rect -3894 658338 -3658 658574
rect -3574 658338 -3338 658574
rect -3894 622658 -3658 622894
rect -3574 622658 -3338 622894
rect -3894 622338 -3658 622574
rect -3574 622338 -3338 622574
rect -3894 586658 -3658 586894
rect -3574 586658 -3338 586894
rect -3894 586338 -3658 586574
rect -3574 586338 -3338 586574
rect -3894 550658 -3658 550894
rect -3574 550658 -3338 550894
rect -3894 550338 -3658 550574
rect -3574 550338 -3338 550574
rect -3894 514658 -3658 514894
rect -3574 514658 -3338 514894
rect -3894 514338 -3658 514574
rect -3574 514338 -3338 514574
rect -3894 478658 -3658 478894
rect -3574 478658 -3338 478894
rect -3894 478338 -3658 478574
rect -3574 478338 -3338 478574
rect -3894 442658 -3658 442894
rect -3574 442658 -3338 442894
rect -3894 442338 -3658 442574
rect -3574 442338 -3338 442574
rect -3894 406658 -3658 406894
rect -3574 406658 -3338 406894
rect -3894 406338 -3658 406574
rect -3574 406338 -3338 406574
rect -3894 370658 -3658 370894
rect -3574 370658 -3338 370894
rect -3894 370338 -3658 370574
rect -3574 370338 -3338 370574
rect -3894 334658 -3658 334894
rect -3574 334658 -3338 334894
rect -3894 334338 -3658 334574
rect -3574 334338 -3338 334574
rect -3894 298658 -3658 298894
rect -3574 298658 -3338 298894
rect -3894 298338 -3658 298574
rect -3574 298338 -3338 298574
rect -3894 262658 -3658 262894
rect -3574 262658 -3338 262894
rect -3894 262338 -3658 262574
rect -3574 262338 -3338 262574
rect -3894 226658 -3658 226894
rect -3574 226658 -3338 226894
rect -3894 226338 -3658 226574
rect -3574 226338 -3338 226574
rect -3894 190658 -3658 190894
rect -3574 190658 -3338 190894
rect -3894 190338 -3658 190574
rect -3574 190338 -3338 190574
rect -3894 154658 -3658 154894
rect -3574 154658 -3338 154894
rect -3894 154338 -3658 154574
rect -3574 154338 -3338 154574
rect -3894 118658 -3658 118894
rect -3574 118658 -3338 118894
rect -3894 118338 -3658 118574
rect -3574 118338 -3338 118574
rect -3894 82658 -3658 82894
rect -3574 82658 -3338 82894
rect -3894 82338 -3658 82574
rect -3574 82338 -3338 82574
rect -3894 46658 -3658 46894
rect -3574 46658 -3338 46894
rect -3894 46338 -3658 46574
rect -3574 46338 -3338 46574
rect -3894 10658 -3658 10894
rect -3574 10658 -3338 10894
rect -3894 10338 -3658 10574
rect -3574 10338 -3338 10574
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 9266 706522 9502 706758
rect 9586 706522 9822 706758
rect 9266 706202 9502 706438
rect 9586 706202 9822 706438
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 9266 -2502 9502 -2266
rect 9586 -2502 9822 -2266
rect 9266 -2822 9502 -2586
rect 9586 -2822 9822 -2586
rect 12986 707482 13222 707718
rect 13306 707482 13542 707718
rect 12986 707162 13222 707398
rect 13306 707162 13542 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect 12986 -3462 13222 -3226
rect 13306 -3462 13542 -3226
rect 12986 -3782 13222 -3546
rect 13306 -3782 13542 -3546
rect 16706 708442 16942 708678
rect 17026 708442 17262 708678
rect 16706 708122 16942 708358
rect 17026 708122 17262 708358
rect 16706 666098 16942 666334
rect 17026 666098 17262 666334
rect 16706 665778 16942 666014
rect 17026 665778 17262 666014
rect 16706 630098 16942 630334
rect 17026 630098 17262 630334
rect 16706 629778 16942 630014
rect 17026 629778 17262 630014
rect 16706 594098 16942 594334
rect 17026 594098 17262 594334
rect 16706 593778 16942 594014
rect 17026 593778 17262 594014
rect 16706 558098 16942 558334
rect 17026 558098 17262 558334
rect 16706 557778 16942 558014
rect 17026 557778 17262 558014
rect 16706 522098 16942 522334
rect 17026 522098 17262 522334
rect 16706 521778 16942 522014
rect 17026 521778 17262 522014
rect 16706 486098 16942 486334
rect 17026 486098 17262 486334
rect 16706 485778 16942 486014
rect 17026 485778 17262 486014
rect 16706 450098 16942 450334
rect 17026 450098 17262 450334
rect 16706 449778 16942 450014
rect 17026 449778 17262 450014
rect 16706 414098 16942 414334
rect 17026 414098 17262 414334
rect 16706 413778 16942 414014
rect 17026 413778 17262 414014
rect 16706 378098 16942 378334
rect 17026 378098 17262 378334
rect 16706 377778 16942 378014
rect 17026 377778 17262 378014
rect 16706 342098 16942 342334
rect 17026 342098 17262 342334
rect 16706 341778 16942 342014
rect 17026 341778 17262 342014
rect 16706 306098 16942 306334
rect 17026 306098 17262 306334
rect 16706 305778 16942 306014
rect 17026 305778 17262 306014
rect 16706 270098 16942 270334
rect 17026 270098 17262 270334
rect 16706 269778 16942 270014
rect 17026 269778 17262 270014
rect 16706 234098 16942 234334
rect 17026 234098 17262 234334
rect 16706 233778 16942 234014
rect 17026 233778 17262 234014
rect 16706 198098 16942 198334
rect 17026 198098 17262 198334
rect 16706 197778 16942 198014
rect 17026 197778 17262 198014
rect 16706 162098 16942 162334
rect 17026 162098 17262 162334
rect 16706 161778 16942 162014
rect 17026 161778 17262 162014
rect 16706 126098 16942 126334
rect 17026 126098 17262 126334
rect 16706 125778 16942 126014
rect 17026 125778 17262 126014
rect 16706 90098 16942 90334
rect 17026 90098 17262 90334
rect 16706 89778 16942 90014
rect 17026 89778 17262 90014
rect 16706 54098 16942 54334
rect 17026 54098 17262 54334
rect 16706 53778 16942 54014
rect 17026 53778 17262 54014
rect 16706 18098 16942 18334
rect 17026 18098 17262 18334
rect 16706 17778 16942 18014
rect 17026 17778 17262 18014
rect 16706 -4422 16942 -4186
rect 17026 -4422 17262 -4186
rect 16706 -4742 16942 -4506
rect 17026 -4742 17262 -4506
rect 20426 709402 20662 709638
rect 20746 709402 20982 709638
rect 20426 709082 20662 709318
rect 20746 709082 20982 709318
rect 20426 669818 20662 670054
rect 20746 669818 20982 670054
rect 20426 669498 20662 669734
rect 20746 669498 20982 669734
rect 20426 633818 20662 634054
rect 20746 633818 20982 634054
rect 20426 633498 20662 633734
rect 20746 633498 20982 633734
rect 20426 597818 20662 598054
rect 20746 597818 20982 598054
rect 20426 597498 20662 597734
rect 20746 597498 20982 597734
rect 20426 561818 20662 562054
rect 20746 561818 20982 562054
rect 20426 561498 20662 561734
rect 20746 561498 20982 561734
rect 20426 525818 20662 526054
rect 20746 525818 20982 526054
rect 20426 525498 20662 525734
rect 20746 525498 20982 525734
rect 20426 489818 20662 490054
rect 20746 489818 20982 490054
rect 20426 489498 20662 489734
rect 20746 489498 20982 489734
rect 20426 453818 20662 454054
rect 20746 453818 20982 454054
rect 20426 453498 20662 453734
rect 20746 453498 20982 453734
rect 20426 417818 20662 418054
rect 20746 417818 20982 418054
rect 20426 417498 20662 417734
rect 20746 417498 20982 417734
rect 20426 381818 20662 382054
rect 20746 381818 20982 382054
rect 20426 381498 20662 381734
rect 20746 381498 20982 381734
rect 20426 345818 20662 346054
rect 20746 345818 20982 346054
rect 20426 345498 20662 345734
rect 20746 345498 20982 345734
rect 20426 309818 20662 310054
rect 20746 309818 20982 310054
rect 20426 309498 20662 309734
rect 20746 309498 20982 309734
rect 20426 273818 20662 274054
rect 20746 273818 20982 274054
rect 20426 273498 20662 273734
rect 20746 273498 20982 273734
rect 20426 237818 20662 238054
rect 20746 237818 20982 238054
rect 20426 237498 20662 237734
rect 20746 237498 20982 237734
rect 20426 201818 20662 202054
rect 20746 201818 20982 202054
rect 20426 201498 20662 201734
rect 20746 201498 20982 201734
rect 20426 165818 20662 166054
rect 20746 165818 20982 166054
rect 20426 165498 20662 165734
rect 20746 165498 20982 165734
rect 20426 129818 20662 130054
rect 20746 129818 20982 130054
rect 20426 129498 20662 129734
rect 20746 129498 20982 129734
rect 20426 93818 20662 94054
rect 20746 93818 20982 94054
rect 20426 93498 20662 93734
rect 20746 93498 20982 93734
rect 20426 57818 20662 58054
rect 20746 57818 20982 58054
rect 20426 57498 20662 57734
rect 20746 57498 20982 57734
rect 20426 21818 20662 22054
rect 20746 21818 20982 22054
rect 20426 21498 20662 21734
rect 20746 21498 20982 21734
rect 20426 -5382 20662 -5146
rect 20746 -5382 20982 -5146
rect 20426 -5702 20662 -5466
rect 20746 -5702 20982 -5466
rect 24146 710362 24382 710598
rect 24466 710362 24702 710598
rect 24146 710042 24382 710278
rect 24466 710042 24702 710278
rect 24146 673538 24382 673774
rect 24466 673538 24702 673774
rect 24146 673218 24382 673454
rect 24466 673218 24702 673454
rect 24146 637538 24382 637774
rect 24466 637538 24702 637774
rect 24146 637218 24382 637454
rect 24466 637218 24702 637454
rect 24146 601538 24382 601774
rect 24466 601538 24702 601774
rect 24146 601218 24382 601454
rect 24466 601218 24702 601454
rect 24146 565538 24382 565774
rect 24466 565538 24702 565774
rect 24146 565218 24382 565454
rect 24466 565218 24702 565454
rect 24146 529538 24382 529774
rect 24466 529538 24702 529774
rect 24146 529218 24382 529454
rect 24466 529218 24702 529454
rect 24146 493538 24382 493774
rect 24466 493538 24702 493774
rect 24146 493218 24382 493454
rect 24466 493218 24702 493454
rect 24146 457538 24382 457774
rect 24466 457538 24702 457774
rect 24146 457218 24382 457454
rect 24466 457218 24702 457454
rect 24146 421538 24382 421774
rect 24466 421538 24702 421774
rect 24146 421218 24382 421454
rect 24466 421218 24702 421454
rect 24146 385538 24382 385774
rect 24466 385538 24702 385774
rect 24146 385218 24382 385454
rect 24466 385218 24702 385454
rect 24146 349538 24382 349774
rect 24466 349538 24702 349774
rect 24146 349218 24382 349454
rect 24466 349218 24702 349454
rect 24146 313538 24382 313774
rect 24466 313538 24702 313774
rect 24146 313218 24382 313454
rect 24466 313218 24702 313454
rect 24146 277538 24382 277774
rect 24466 277538 24702 277774
rect 24146 277218 24382 277454
rect 24466 277218 24702 277454
rect 24146 241538 24382 241774
rect 24466 241538 24702 241774
rect 24146 241218 24382 241454
rect 24466 241218 24702 241454
rect 24146 205538 24382 205774
rect 24466 205538 24702 205774
rect 24146 205218 24382 205454
rect 24466 205218 24702 205454
rect 24146 169538 24382 169774
rect 24466 169538 24702 169774
rect 24146 169218 24382 169454
rect 24466 169218 24702 169454
rect 24146 133538 24382 133774
rect 24466 133538 24702 133774
rect 24146 133218 24382 133454
rect 24466 133218 24702 133454
rect 24146 97538 24382 97774
rect 24466 97538 24702 97774
rect 24146 97218 24382 97454
rect 24466 97218 24702 97454
rect 24146 61538 24382 61774
rect 24466 61538 24702 61774
rect 24146 61218 24382 61454
rect 24466 61218 24702 61454
rect 24146 25538 24382 25774
rect 24466 25538 24702 25774
rect 24146 25218 24382 25454
rect 24466 25218 24702 25454
rect 24146 -6342 24382 -6106
rect 24466 -6342 24702 -6106
rect 24146 -6662 24382 -6426
rect 24466 -6662 24702 -6426
rect 27866 711322 28102 711558
rect 28186 711322 28422 711558
rect 27866 711002 28102 711238
rect 28186 711002 28422 711238
rect 27866 677258 28102 677494
rect 28186 677258 28422 677494
rect 27866 676938 28102 677174
rect 28186 676938 28422 677174
rect 27866 641258 28102 641494
rect 28186 641258 28422 641494
rect 27866 640938 28102 641174
rect 28186 640938 28422 641174
rect 27866 605258 28102 605494
rect 28186 605258 28422 605494
rect 27866 604938 28102 605174
rect 28186 604938 28422 605174
rect 27866 569258 28102 569494
rect 28186 569258 28422 569494
rect 27866 568938 28102 569174
rect 28186 568938 28422 569174
rect 27866 533258 28102 533494
rect 28186 533258 28422 533494
rect 27866 532938 28102 533174
rect 28186 532938 28422 533174
rect 27866 497258 28102 497494
rect 28186 497258 28422 497494
rect 27866 496938 28102 497174
rect 28186 496938 28422 497174
rect 27866 461258 28102 461494
rect 28186 461258 28422 461494
rect 27866 460938 28102 461174
rect 28186 460938 28422 461174
rect 27866 425258 28102 425494
rect 28186 425258 28422 425494
rect 27866 424938 28102 425174
rect 28186 424938 28422 425174
rect 27866 389258 28102 389494
rect 28186 389258 28422 389494
rect 27866 388938 28102 389174
rect 28186 388938 28422 389174
rect 27866 353258 28102 353494
rect 28186 353258 28422 353494
rect 27866 352938 28102 353174
rect 28186 352938 28422 353174
rect 27866 317258 28102 317494
rect 28186 317258 28422 317494
rect 27866 316938 28102 317174
rect 28186 316938 28422 317174
rect 27866 281258 28102 281494
rect 28186 281258 28422 281494
rect 27866 280938 28102 281174
rect 28186 280938 28422 281174
rect 27866 245258 28102 245494
rect 28186 245258 28422 245494
rect 27866 244938 28102 245174
rect 28186 244938 28422 245174
rect 27866 209258 28102 209494
rect 28186 209258 28422 209494
rect 27866 208938 28102 209174
rect 28186 208938 28422 209174
rect 27866 173258 28102 173494
rect 28186 173258 28422 173494
rect 27866 172938 28102 173174
rect 28186 172938 28422 173174
rect 27866 137258 28102 137494
rect 28186 137258 28422 137494
rect 27866 136938 28102 137174
rect 28186 136938 28422 137174
rect 27866 101258 28102 101494
rect 28186 101258 28422 101494
rect 27866 100938 28102 101174
rect 28186 100938 28422 101174
rect 27866 65258 28102 65494
rect 28186 65258 28422 65494
rect 27866 64938 28102 65174
rect 28186 64938 28422 65174
rect 27866 29258 28102 29494
rect 28186 29258 28422 29494
rect 27866 28938 28102 29174
rect 28186 28938 28422 29174
rect 27866 -7302 28102 -7066
rect 28186 -7302 28422 -7066
rect 27866 -7622 28102 -7386
rect 28186 -7622 28422 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 45266 706522 45502 706758
rect 45586 706522 45822 706758
rect 45266 706202 45502 706438
rect 45586 706202 45822 706438
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 48986 707482 49222 707718
rect 49306 707482 49542 707718
rect 48986 707162 49222 707398
rect 49306 707162 49542 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -2502 45502 -2266
rect 45586 -2502 45822 -2266
rect 45266 -2822 45502 -2586
rect 45586 -2822 45822 -2586
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 48986 -3462 49222 -3226
rect 49306 -3462 49542 -3226
rect 48986 -3782 49222 -3546
rect 49306 -3782 49542 -3546
rect 52706 708442 52942 708678
rect 53026 708442 53262 708678
rect 52706 708122 52942 708358
rect 53026 708122 53262 708358
rect 52706 666098 52942 666334
rect 53026 666098 53262 666334
rect 52706 665778 52942 666014
rect 53026 665778 53262 666014
rect 52706 630098 52942 630334
rect 53026 630098 53262 630334
rect 52706 629778 52942 630014
rect 53026 629778 53262 630014
rect 52706 594098 52942 594334
rect 53026 594098 53262 594334
rect 52706 593778 52942 594014
rect 53026 593778 53262 594014
rect 52706 558098 52942 558334
rect 53026 558098 53262 558334
rect 52706 557778 52942 558014
rect 53026 557778 53262 558014
rect 52706 522098 52942 522334
rect 53026 522098 53262 522334
rect 52706 521778 52942 522014
rect 53026 521778 53262 522014
rect 52706 486098 52942 486334
rect 53026 486098 53262 486334
rect 52706 485778 52942 486014
rect 53026 485778 53262 486014
rect 52706 450098 52942 450334
rect 53026 450098 53262 450334
rect 52706 449778 52942 450014
rect 53026 449778 53262 450014
rect 52706 414098 52942 414334
rect 53026 414098 53262 414334
rect 52706 413778 52942 414014
rect 53026 413778 53262 414014
rect 52706 378098 52942 378334
rect 53026 378098 53262 378334
rect 52706 377778 52942 378014
rect 53026 377778 53262 378014
rect 52706 342098 52942 342334
rect 53026 342098 53262 342334
rect 52706 341778 52942 342014
rect 53026 341778 53262 342014
rect 56426 709402 56662 709638
rect 56746 709402 56982 709638
rect 56426 709082 56662 709318
rect 56746 709082 56982 709318
rect 60146 710362 60382 710598
rect 60466 710362 60702 710598
rect 60146 710042 60382 710278
rect 60466 710042 60702 710278
rect 60146 673538 60382 673774
rect 60466 673538 60702 673774
rect 60146 673218 60382 673454
rect 60466 673218 60702 673454
rect 56426 669818 56662 670054
rect 56746 669818 56982 670054
rect 56426 669498 56662 669734
rect 56746 669498 56982 669734
rect 56426 633818 56662 634054
rect 56746 633818 56982 634054
rect 56426 633498 56662 633734
rect 56746 633498 56982 633734
rect 56426 597818 56662 598054
rect 56746 597818 56982 598054
rect 56426 597498 56662 597734
rect 56746 597498 56982 597734
rect 56426 561818 56662 562054
rect 56746 561818 56982 562054
rect 56426 561498 56662 561734
rect 56746 561498 56982 561734
rect 56426 525818 56662 526054
rect 56746 525818 56982 526054
rect 56426 525498 56662 525734
rect 56746 525498 56982 525734
rect 56426 489818 56662 490054
rect 56746 489818 56982 490054
rect 56426 489498 56662 489734
rect 56746 489498 56982 489734
rect 56426 453818 56662 454054
rect 56746 453818 56982 454054
rect 56426 453498 56662 453734
rect 56746 453498 56982 453734
rect 60146 637538 60382 637774
rect 60466 637538 60702 637774
rect 60146 637218 60382 637454
rect 60466 637218 60702 637454
rect 60146 601538 60382 601774
rect 60466 601538 60702 601774
rect 60146 601218 60382 601454
rect 60466 601218 60702 601454
rect 63866 711322 64102 711558
rect 64186 711322 64422 711558
rect 63866 711002 64102 711238
rect 64186 711002 64422 711238
rect 63866 677258 64102 677494
rect 64186 677258 64422 677494
rect 63866 676938 64102 677174
rect 64186 676938 64422 677174
rect 63866 641258 64102 641494
rect 64186 641258 64422 641494
rect 63866 640938 64102 641174
rect 64186 640938 64422 641174
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 81266 706522 81502 706758
rect 81586 706522 81822 706758
rect 81266 706202 81502 706438
rect 81586 706202 81822 706438
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 84986 707482 85222 707718
rect 85306 707482 85542 707718
rect 84986 707162 85222 707398
rect 85306 707162 85542 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 88706 708442 88942 708678
rect 89026 708442 89262 708678
rect 88706 708122 88942 708358
rect 89026 708122 89262 708358
rect 88706 666098 88942 666334
rect 89026 666098 89262 666334
rect 88706 665778 88942 666014
rect 89026 665778 89262 666014
rect 88706 630098 88942 630334
rect 89026 630098 89262 630334
rect 88706 629778 88942 630014
rect 89026 629778 89262 630014
rect 92426 709402 92662 709638
rect 92746 709402 92982 709638
rect 92426 709082 92662 709318
rect 92746 709082 92982 709318
rect 92426 669818 92662 670054
rect 92746 669818 92982 670054
rect 92426 669498 92662 669734
rect 92746 669498 92982 669734
rect 92426 633818 92662 634054
rect 92746 633818 92982 634054
rect 92426 633498 92662 633734
rect 92746 633498 92982 633734
rect 96146 710362 96382 710598
rect 96466 710362 96702 710598
rect 96146 710042 96382 710278
rect 96466 710042 96702 710278
rect 96146 673538 96382 673774
rect 96466 673538 96702 673774
rect 96146 673218 96382 673454
rect 96466 673218 96702 673454
rect 96146 637538 96382 637774
rect 96466 637538 96702 637774
rect 96146 637218 96382 637454
rect 96466 637218 96702 637454
rect 99866 711322 100102 711558
rect 100186 711322 100422 711558
rect 99866 711002 100102 711238
rect 100186 711002 100422 711238
rect 99866 677258 100102 677494
rect 100186 677258 100422 677494
rect 99866 676938 100102 677174
rect 100186 676938 100422 677174
rect 99866 641258 100102 641494
rect 100186 641258 100422 641494
rect 99866 640938 100102 641174
rect 100186 640938 100422 641174
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 117266 706522 117502 706758
rect 117586 706522 117822 706758
rect 117266 706202 117502 706438
rect 117586 706202 117822 706438
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 120986 707482 121222 707718
rect 121306 707482 121542 707718
rect 120986 707162 121222 707398
rect 121306 707162 121542 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 124706 708442 124942 708678
rect 125026 708442 125262 708678
rect 124706 708122 124942 708358
rect 125026 708122 125262 708358
rect 124706 666098 124942 666334
rect 125026 666098 125262 666334
rect 124706 665778 124942 666014
rect 125026 665778 125262 666014
rect 124706 630098 124942 630334
rect 125026 630098 125262 630334
rect 124706 629778 124942 630014
rect 125026 629778 125262 630014
rect 128426 709402 128662 709638
rect 128746 709402 128982 709638
rect 128426 709082 128662 709318
rect 128746 709082 128982 709318
rect 128426 669818 128662 670054
rect 128746 669818 128982 670054
rect 128426 669498 128662 669734
rect 128746 669498 128982 669734
rect 128426 633818 128662 634054
rect 128746 633818 128982 634054
rect 128426 633498 128662 633734
rect 128746 633498 128982 633734
rect 132146 710362 132382 710598
rect 132466 710362 132702 710598
rect 132146 710042 132382 710278
rect 132466 710042 132702 710278
rect 132146 673538 132382 673774
rect 132466 673538 132702 673774
rect 132146 673218 132382 673454
rect 132466 673218 132702 673454
rect 132146 637538 132382 637774
rect 132466 637538 132702 637774
rect 132146 637218 132382 637454
rect 132466 637218 132702 637454
rect 135866 711322 136102 711558
rect 136186 711322 136422 711558
rect 135866 711002 136102 711238
rect 136186 711002 136422 711238
rect 135866 677258 136102 677494
rect 136186 677258 136422 677494
rect 135866 676938 136102 677174
rect 136186 676938 136422 677174
rect 135866 641258 136102 641494
rect 136186 641258 136422 641494
rect 135866 640938 136102 641174
rect 136186 640938 136422 641174
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 153266 706522 153502 706758
rect 153586 706522 153822 706758
rect 153266 706202 153502 706438
rect 153586 706202 153822 706438
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 156986 707482 157222 707718
rect 157306 707482 157542 707718
rect 156986 707162 157222 707398
rect 157306 707162 157542 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 160706 708442 160942 708678
rect 161026 708442 161262 708678
rect 160706 708122 160942 708358
rect 161026 708122 161262 708358
rect 160706 666098 160942 666334
rect 161026 666098 161262 666334
rect 160706 665778 160942 666014
rect 161026 665778 161262 666014
rect 160706 630098 160942 630334
rect 161026 630098 161262 630334
rect 160706 629778 160942 630014
rect 161026 629778 161262 630014
rect 164426 709402 164662 709638
rect 164746 709402 164982 709638
rect 164426 709082 164662 709318
rect 164746 709082 164982 709318
rect 164426 669818 164662 670054
rect 164746 669818 164982 670054
rect 164426 669498 164662 669734
rect 164746 669498 164982 669734
rect 164426 633818 164662 634054
rect 164746 633818 164982 634054
rect 164426 633498 164662 633734
rect 164746 633498 164982 633734
rect 168146 710362 168382 710598
rect 168466 710362 168702 710598
rect 168146 710042 168382 710278
rect 168466 710042 168702 710278
rect 168146 673538 168382 673774
rect 168466 673538 168702 673774
rect 168146 673218 168382 673454
rect 168466 673218 168702 673454
rect 168146 637538 168382 637774
rect 168466 637538 168702 637774
rect 168146 637218 168382 637454
rect 168466 637218 168702 637454
rect 171866 711322 172102 711558
rect 172186 711322 172422 711558
rect 171866 711002 172102 711238
rect 172186 711002 172422 711238
rect 171866 677258 172102 677494
rect 172186 677258 172422 677494
rect 171866 676938 172102 677174
rect 172186 676938 172422 677174
rect 171866 641258 172102 641494
rect 172186 641258 172422 641494
rect 171866 640938 172102 641174
rect 172186 640938 172422 641174
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 189266 706522 189502 706758
rect 189586 706522 189822 706758
rect 189266 706202 189502 706438
rect 189586 706202 189822 706438
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 192986 707482 193222 707718
rect 193306 707482 193542 707718
rect 192986 707162 193222 707398
rect 193306 707162 193542 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 196706 708442 196942 708678
rect 197026 708442 197262 708678
rect 196706 708122 196942 708358
rect 197026 708122 197262 708358
rect 196706 666098 196942 666334
rect 197026 666098 197262 666334
rect 196706 665778 196942 666014
rect 197026 665778 197262 666014
rect 196706 630098 196942 630334
rect 197026 630098 197262 630334
rect 196706 629778 196942 630014
rect 197026 629778 197262 630014
rect 200426 709402 200662 709638
rect 200746 709402 200982 709638
rect 200426 709082 200662 709318
rect 200746 709082 200982 709318
rect 200426 669818 200662 670054
rect 200746 669818 200982 670054
rect 200426 669498 200662 669734
rect 200746 669498 200982 669734
rect 200426 633818 200662 634054
rect 200746 633818 200982 634054
rect 200426 633498 200662 633734
rect 200746 633498 200982 633734
rect 204146 710362 204382 710598
rect 204466 710362 204702 710598
rect 204146 710042 204382 710278
rect 204466 710042 204702 710278
rect 204146 673538 204382 673774
rect 204466 673538 204702 673774
rect 204146 673218 204382 673454
rect 204466 673218 204702 673454
rect 204146 637538 204382 637774
rect 204466 637538 204702 637774
rect 204146 637218 204382 637454
rect 204466 637218 204702 637454
rect 207866 711322 208102 711558
rect 208186 711322 208422 711558
rect 207866 711002 208102 711238
rect 208186 711002 208422 711238
rect 207866 677258 208102 677494
rect 208186 677258 208422 677494
rect 207866 676938 208102 677174
rect 208186 676938 208422 677174
rect 207866 641258 208102 641494
rect 208186 641258 208422 641494
rect 207866 640938 208102 641174
rect 208186 640938 208422 641174
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 225266 706522 225502 706758
rect 225586 706522 225822 706758
rect 225266 706202 225502 706438
rect 225586 706202 225822 706438
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 228986 707482 229222 707718
rect 229306 707482 229542 707718
rect 228986 707162 229222 707398
rect 229306 707162 229542 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 232706 708442 232942 708678
rect 233026 708442 233262 708678
rect 232706 708122 232942 708358
rect 233026 708122 233262 708358
rect 232706 666098 232942 666334
rect 233026 666098 233262 666334
rect 232706 665778 232942 666014
rect 233026 665778 233262 666014
rect 232706 630098 232942 630334
rect 233026 630098 233262 630334
rect 232706 629778 232942 630014
rect 233026 629778 233262 630014
rect 236426 709402 236662 709638
rect 236746 709402 236982 709638
rect 236426 709082 236662 709318
rect 236746 709082 236982 709318
rect 236426 669818 236662 670054
rect 236746 669818 236982 670054
rect 236426 669498 236662 669734
rect 236746 669498 236982 669734
rect 236426 633818 236662 634054
rect 236746 633818 236982 634054
rect 236426 633498 236662 633734
rect 236746 633498 236982 633734
rect 240146 710362 240382 710598
rect 240466 710362 240702 710598
rect 240146 710042 240382 710278
rect 240466 710042 240702 710278
rect 240146 673538 240382 673774
rect 240466 673538 240702 673774
rect 240146 673218 240382 673454
rect 240466 673218 240702 673454
rect 240146 637538 240382 637774
rect 240466 637538 240702 637774
rect 240146 637218 240382 637454
rect 240466 637218 240702 637454
rect 243866 711322 244102 711558
rect 244186 711322 244422 711558
rect 243866 711002 244102 711238
rect 244186 711002 244422 711238
rect 243866 677258 244102 677494
rect 244186 677258 244422 677494
rect 243866 676938 244102 677174
rect 244186 676938 244422 677174
rect 243866 641258 244102 641494
rect 244186 641258 244422 641494
rect 243866 640938 244102 641174
rect 244186 640938 244422 641174
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 261266 706522 261502 706758
rect 261586 706522 261822 706758
rect 261266 706202 261502 706438
rect 261586 706202 261822 706438
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 264986 707482 265222 707718
rect 265306 707482 265542 707718
rect 264986 707162 265222 707398
rect 265306 707162 265542 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 268706 708442 268942 708678
rect 269026 708442 269262 708678
rect 268706 708122 268942 708358
rect 269026 708122 269262 708358
rect 268706 666098 268942 666334
rect 269026 666098 269262 666334
rect 268706 665778 268942 666014
rect 269026 665778 269262 666014
rect 268706 630098 268942 630334
rect 269026 630098 269262 630334
rect 268706 629778 268942 630014
rect 269026 629778 269262 630014
rect 272426 709402 272662 709638
rect 272746 709402 272982 709638
rect 272426 709082 272662 709318
rect 272746 709082 272982 709318
rect 272426 669818 272662 670054
rect 272746 669818 272982 670054
rect 272426 669498 272662 669734
rect 272746 669498 272982 669734
rect 272426 633818 272662 634054
rect 272746 633818 272982 634054
rect 272426 633498 272662 633734
rect 272746 633498 272982 633734
rect 276146 710362 276382 710598
rect 276466 710362 276702 710598
rect 276146 710042 276382 710278
rect 276466 710042 276702 710278
rect 276146 673538 276382 673774
rect 276466 673538 276702 673774
rect 276146 673218 276382 673454
rect 276466 673218 276702 673454
rect 276146 637538 276382 637774
rect 276466 637538 276702 637774
rect 276146 637218 276382 637454
rect 276466 637218 276702 637454
rect 279866 711322 280102 711558
rect 280186 711322 280422 711558
rect 279866 711002 280102 711238
rect 280186 711002 280422 711238
rect 279866 677258 280102 677494
rect 280186 677258 280422 677494
rect 279866 676938 280102 677174
rect 280186 676938 280422 677174
rect 279866 641258 280102 641494
rect 280186 641258 280422 641494
rect 279866 640938 280102 641174
rect 280186 640938 280422 641174
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 63866 605258 64102 605494
rect 64186 605258 64422 605494
rect 63866 604938 64102 605174
rect 64186 604938 64422 605174
rect 60146 565538 60382 565774
rect 60466 565538 60702 565774
rect 60146 565218 60382 565454
rect 60466 565218 60702 565454
rect 60146 529538 60382 529774
rect 60466 529538 60702 529774
rect 60146 529218 60382 529454
rect 60466 529218 60702 529454
rect 60146 493538 60382 493774
rect 60466 493538 60702 493774
rect 60146 493218 60382 493454
rect 60466 493218 60702 493454
rect 60146 457538 60382 457774
rect 60466 457538 60702 457774
rect 60146 457218 60382 457454
rect 60466 457218 60702 457454
rect 56426 417818 56662 418054
rect 56746 417818 56982 418054
rect 56426 417498 56662 417734
rect 56746 417498 56982 417734
rect 56426 381818 56662 382054
rect 56746 381818 56982 382054
rect 56426 381498 56662 381734
rect 56746 381498 56982 381734
rect 56426 345818 56662 346054
rect 56746 345818 56982 346054
rect 56426 345498 56662 345734
rect 56746 345498 56982 345734
rect 54250 327218 54486 327454
rect 54250 326898 54486 327134
rect 52706 306098 52942 306334
rect 53026 306098 53262 306334
rect 52706 305778 52942 306014
rect 53026 305778 53262 306014
rect 60146 421538 60382 421774
rect 60466 421538 60702 421774
rect 60146 421218 60382 421454
rect 60466 421218 60702 421454
rect 60146 385538 60382 385774
rect 60466 385538 60702 385774
rect 60146 385218 60382 385454
rect 60466 385218 60702 385454
rect 60146 349538 60382 349774
rect 60466 349538 60702 349774
rect 60146 349218 60382 349454
rect 60466 349218 60702 349454
rect 63866 569258 64102 569494
rect 64186 569258 64422 569494
rect 63866 568938 64102 569174
rect 64186 568938 64422 569174
rect 63866 533258 64102 533494
rect 64186 533258 64422 533494
rect 63866 532938 64102 533174
rect 64186 532938 64422 533174
rect 63866 497258 64102 497494
rect 64186 497258 64422 497494
rect 63866 496938 64102 497174
rect 64186 496938 64422 497174
rect 63866 461258 64102 461494
rect 64186 461258 64422 461494
rect 63866 460938 64102 461174
rect 64186 460938 64422 461174
rect 63866 425258 64102 425494
rect 64186 425258 64422 425494
rect 63866 424938 64102 425174
rect 64186 424938 64422 425174
rect 63866 389258 64102 389494
rect 64186 389258 64422 389494
rect 63866 388938 64102 389174
rect 64186 388938 64422 389174
rect 63866 353258 64102 353494
rect 64186 353258 64422 353494
rect 63866 352938 64102 353174
rect 64186 352938 64422 353174
rect 89610 618938 89846 619174
rect 89610 618618 89846 618854
rect 120330 618938 120566 619174
rect 120330 618618 120566 618854
rect 151050 618938 151286 619174
rect 151050 618618 151286 618854
rect 181770 618938 182006 619174
rect 181770 618618 182006 618854
rect 212490 618938 212726 619174
rect 212490 618618 212726 618854
rect 243210 618938 243446 619174
rect 243210 618618 243446 618854
rect 273930 618938 274166 619174
rect 273930 618618 274166 618854
rect 74250 615218 74486 615454
rect 74250 614898 74486 615134
rect 104970 615218 105206 615454
rect 104970 614898 105206 615134
rect 135690 615218 135926 615454
rect 135690 614898 135926 615134
rect 166410 615218 166646 615454
rect 166410 614898 166646 615134
rect 197130 615218 197366 615454
rect 197130 614898 197366 615134
rect 227850 615218 228086 615454
rect 227850 614898 228086 615134
rect 258570 615218 258806 615454
rect 258570 614898 258806 615134
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 89610 582938 89846 583174
rect 89610 582618 89846 582854
rect 120330 582938 120566 583174
rect 120330 582618 120566 582854
rect 151050 582938 151286 583174
rect 151050 582618 151286 582854
rect 181770 582938 182006 583174
rect 181770 582618 182006 582854
rect 212490 582938 212726 583174
rect 212490 582618 212726 582854
rect 243210 582938 243446 583174
rect 243210 582618 243446 582854
rect 273930 582938 274166 583174
rect 273930 582618 274166 582854
rect 74250 579218 74486 579454
rect 74250 578898 74486 579134
rect 104970 579218 105206 579454
rect 104970 578898 105206 579134
rect 135690 579218 135926 579454
rect 135690 578898 135926 579134
rect 166410 579218 166646 579454
rect 166410 578898 166646 579134
rect 197130 579218 197366 579454
rect 197130 578898 197366 579134
rect 227850 579218 228086 579454
rect 227850 578898 228086 579134
rect 258570 579218 258806 579454
rect 258570 578898 258806 579134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 89610 546938 89846 547174
rect 89610 546618 89846 546854
rect 120330 546938 120566 547174
rect 120330 546618 120566 546854
rect 151050 546938 151286 547174
rect 151050 546618 151286 546854
rect 181770 546938 182006 547174
rect 181770 546618 182006 546854
rect 212490 546938 212726 547174
rect 212490 546618 212726 546854
rect 243210 546938 243446 547174
rect 243210 546618 243446 546854
rect 273930 546938 274166 547174
rect 273930 546618 274166 546854
rect 74250 543218 74486 543454
rect 74250 542898 74486 543134
rect 104970 543218 105206 543454
rect 104970 542898 105206 543134
rect 135690 543218 135926 543454
rect 135690 542898 135926 543134
rect 166410 543218 166646 543454
rect 166410 542898 166646 543134
rect 197130 543218 197366 543454
rect 197130 542898 197366 543134
rect 227850 543218 228086 543454
rect 227850 542898 228086 543134
rect 258570 543218 258806 543454
rect 258570 542898 258806 543134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 89610 510938 89846 511174
rect 89610 510618 89846 510854
rect 120330 510938 120566 511174
rect 120330 510618 120566 510854
rect 151050 510938 151286 511174
rect 151050 510618 151286 510854
rect 181770 510938 182006 511174
rect 181770 510618 182006 510854
rect 212490 510938 212726 511174
rect 212490 510618 212726 510854
rect 243210 510938 243446 511174
rect 243210 510618 243446 510854
rect 273930 510938 274166 511174
rect 273930 510618 274166 510854
rect 74250 507218 74486 507454
rect 74250 506898 74486 507134
rect 104970 507218 105206 507454
rect 104970 506898 105206 507134
rect 135690 507218 135926 507454
rect 135690 506898 135926 507134
rect 166410 507218 166646 507454
rect 166410 506898 166646 507134
rect 197130 507218 197366 507454
rect 197130 506898 197366 507134
rect 227850 507218 228086 507454
rect 227850 506898 228086 507134
rect 258570 507218 258806 507454
rect 258570 506898 258806 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 88706 450098 88942 450334
rect 89026 450098 89262 450334
rect 88706 449778 88942 450014
rect 89026 449778 89262 450014
rect 88706 414098 88942 414334
rect 89026 414098 89262 414334
rect 88706 413778 88942 414014
rect 89026 413778 89262 414014
rect 88706 378098 88942 378334
rect 89026 378098 89262 378334
rect 88706 377778 88942 378014
rect 89026 377778 89262 378014
rect 88706 342098 88942 342334
rect 89026 342098 89262 342334
rect 88706 341778 88942 342014
rect 89026 341778 89262 342014
rect 92426 453818 92662 454054
rect 92746 453818 92982 454054
rect 92426 453498 92662 453734
rect 92746 453498 92982 453734
rect 92426 417818 92662 418054
rect 92746 417818 92982 418054
rect 92426 417498 92662 417734
rect 92746 417498 92982 417734
rect 92426 381818 92662 382054
rect 92746 381818 92982 382054
rect 92426 381498 92662 381734
rect 92746 381498 92982 381734
rect 92426 345818 92662 346054
rect 92746 345818 92982 346054
rect 92426 345498 92662 345734
rect 92746 345498 92982 345734
rect 96146 457538 96382 457774
rect 96466 457538 96702 457774
rect 96146 457218 96382 457454
rect 96466 457218 96702 457454
rect 96146 421538 96382 421774
rect 96466 421538 96702 421774
rect 96146 421218 96382 421454
rect 96466 421218 96702 421454
rect 96146 385538 96382 385774
rect 96466 385538 96702 385774
rect 96146 385218 96382 385454
rect 96466 385218 96702 385454
rect 96146 349538 96382 349774
rect 96466 349538 96702 349774
rect 96146 349218 96382 349454
rect 96466 349218 96702 349454
rect 99866 461258 100102 461494
rect 100186 461258 100422 461494
rect 99866 460938 100102 461174
rect 100186 460938 100422 461174
rect 99866 425258 100102 425494
rect 100186 425258 100422 425494
rect 99866 424938 100102 425174
rect 100186 424938 100422 425174
rect 99866 389258 100102 389494
rect 100186 389258 100422 389494
rect 99866 388938 100102 389174
rect 100186 388938 100422 389174
rect 99866 353258 100102 353494
rect 100186 353258 100422 353494
rect 99866 352938 100102 353174
rect 100186 352938 100422 353174
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 109826 399218 110062 399454
rect 110146 399218 110382 399454
rect 109826 398898 110062 399134
rect 110146 398898 110382 399134
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 69610 330938 69846 331174
rect 69610 330618 69846 330854
rect 100330 330938 100566 331174
rect 100330 330618 100566 330854
rect 84970 327218 85206 327454
rect 84970 326898 85206 327134
rect 56426 309818 56662 310054
rect 56746 309818 56982 310054
rect 56426 309498 56662 309734
rect 56746 309498 56982 309734
rect 54250 291218 54486 291454
rect 54250 290898 54486 291134
rect 52706 270098 52942 270334
rect 53026 270098 53262 270334
rect 52706 269778 52942 270014
rect 53026 269778 53262 270014
rect 52706 234098 52942 234334
rect 53026 234098 53262 234334
rect 52706 233778 52942 234014
rect 53026 233778 53262 234014
rect 52706 198098 52942 198334
rect 53026 198098 53262 198334
rect 52706 197778 52942 198014
rect 53026 197778 53262 198014
rect 52706 162098 52942 162334
rect 53026 162098 53262 162334
rect 52706 161778 52942 162014
rect 53026 161778 53262 162014
rect 52706 126098 52942 126334
rect 53026 126098 53262 126334
rect 52706 125778 52942 126014
rect 53026 125778 53262 126014
rect 52706 90098 52942 90334
rect 53026 90098 53262 90334
rect 52706 89778 52942 90014
rect 53026 89778 53262 90014
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 69610 294938 69846 295174
rect 69610 294618 69846 294854
rect 100330 294938 100566 295174
rect 100330 294618 100566 294854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 84970 291218 85206 291454
rect 84970 290898 85206 291134
rect 56426 273818 56662 274054
rect 56746 273818 56982 274054
rect 56426 273498 56662 273734
rect 56746 273498 56982 273734
rect 56426 237818 56662 238054
rect 56746 237818 56982 238054
rect 56426 237498 56662 237734
rect 56746 237498 56982 237734
rect 56426 201818 56662 202054
rect 56746 201818 56982 202054
rect 56426 201498 56662 201734
rect 56746 201498 56982 201734
rect 56426 165818 56662 166054
rect 56746 165818 56982 166054
rect 56426 165498 56662 165734
rect 56746 165498 56982 165734
rect 56426 129818 56662 130054
rect 56746 129818 56982 130054
rect 56426 129498 56662 129734
rect 56746 129498 56982 129734
rect 56426 93818 56662 94054
rect 56746 93818 56982 94054
rect 56426 93498 56662 93734
rect 56746 93498 56982 93734
rect 55080 75218 55316 75454
rect 55080 74898 55316 75134
rect 52706 54098 52942 54334
rect 53026 54098 53262 54334
rect 52706 53778 52942 54014
rect 53026 53778 53262 54014
rect 52706 18098 52942 18334
rect 53026 18098 53262 18334
rect 52706 17778 52942 18014
rect 53026 17778 53262 18014
rect 52706 -4422 52942 -4186
rect 53026 -4422 53262 -4186
rect 52706 -4742 52942 -4506
rect 53026 -4742 53262 -4506
rect 60146 277538 60382 277774
rect 60466 277538 60702 277774
rect 60146 277218 60382 277454
rect 60466 277218 60702 277454
rect 60146 241538 60382 241774
rect 60466 241538 60702 241774
rect 60146 241218 60382 241454
rect 60466 241218 60702 241454
rect 60146 205538 60382 205774
rect 60466 205538 60702 205774
rect 60146 205218 60382 205454
rect 60466 205218 60702 205454
rect 60146 169538 60382 169774
rect 60466 169538 60702 169774
rect 60146 169218 60382 169454
rect 60466 169218 60702 169454
rect 60146 133538 60382 133774
rect 60466 133538 60702 133774
rect 60146 133218 60382 133454
rect 60466 133218 60702 133454
rect 60146 97538 60382 97774
rect 60466 97538 60702 97774
rect 60146 97218 60382 97454
rect 60466 97218 60702 97454
rect 59174 78938 59410 79174
rect 59174 78618 59410 78854
rect 56426 57818 56662 58054
rect 56746 57818 56982 58054
rect 56426 57498 56662 57734
rect 56746 57498 56982 57734
rect 56426 21818 56662 22054
rect 56746 21818 56982 22054
rect 56426 21498 56662 21734
rect 56746 21498 56982 21734
rect 56426 -5382 56662 -5146
rect 56746 -5382 56982 -5146
rect 56426 -5702 56662 -5466
rect 56746 -5702 56982 -5466
rect 63866 245258 64102 245494
rect 64186 245258 64422 245494
rect 63866 244938 64102 245174
rect 64186 244938 64422 245174
rect 63866 209258 64102 209494
rect 64186 209258 64422 209494
rect 63866 208938 64102 209174
rect 64186 208938 64422 209174
rect 63866 173258 64102 173494
rect 64186 173258 64422 173494
rect 63866 172938 64102 173174
rect 64186 172938 64422 173174
rect 63866 137258 64102 137494
rect 64186 137258 64422 137494
rect 63866 136938 64102 137174
rect 64186 136938 64422 137174
rect 63866 101258 64102 101494
rect 64186 101258 64422 101494
rect 63866 100938 64102 101174
rect 64186 100938 64422 101174
rect 63268 75218 63504 75454
rect 63268 74898 63504 75134
rect 60146 61538 60382 61774
rect 60466 61538 60702 61774
rect 60146 61218 60382 61454
rect 60466 61218 60702 61454
rect 60146 25538 60382 25774
rect 60466 25538 60702 25774
rect 60146 25218 60382 25454
rect 60466 25218 60702 25454
rect 60146 -6342 60382 -6106
rect 60466 -6342 60702 -6106
rect 60146 -6662 60382 -6426
rect 60466 -6662 60702 -6426
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 67362 78938 67598 79174
rect 67362 78618 67598 78854
rect 71456 75218 71692 75454
rect 71456 74898 71692 75134
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 75550 78938 75786 79174
rect 75550 78618 75786 78854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 63866 65258 64102 65494
rect 64186 65258 64422 65494
rect 63866 64938 64102 65174
rect 64186 64938 64422 65174
rect 63866 29258 64102 29494
rect 64186 29258 64422 29494
rect 63866 28938 64102 29174
rect 64186 28938 64422 29174
rect 63866 -7302 64102 -7066
rect 64186 -7302 64422 -7066
rect 63866 -7622 64102 -7386
rect 64186 -7622 64422 -7386
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 79644 75218 79880 75454
rect 79644 74898 79880 75134
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 83738 78938 83974 79174
rect 83738 78618 83974 78854
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -2502 81502 -2266
rect 81586 -2502 81822 -2266
rect 81266 -2822 81502 -2586
rect 81586 -2822 81822 -2586
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 84986 -3462 85222 -3226
rect 85306 -3462 85542 -3226
rect 84986 -3782 85222 -3546
rect 85306 -3782 85542 -3546
rect 88706 270098 88942 270334
rect 89026 270098 89262 270334
rect 88706 269778 88942 270014
rect 89026 269778 89262 270014
rect 88706 234098 88942 234334
rect 89026 234098 89262 234334
rect 88706 233778 88942 234014
rect 89026 233778 89262 234014
rect 88706 198098 88942 198334
rect 89026 198098 89262 198334
rect 88706 197778 88942 198014
rect 89026 197778 89262 198014
rect 88706 162098 88942 162334
rect 89026 162098 89262 162334
rect 88706 161778 88942 162014
rect 89026 161778 89262 162014
rect 88706 126098 88942 126334
rect 89026 126098 89262 126334
rect 88706 125778 88942 126014
rect 89026 125778 89262 126014
rect 88706 90098 88942 90334
rect 89026 90098 89262 90334
rect 88706 89778 88942 90014
rect 89026 89778 89262 90014
rect 88706 54098 88942 54334
rect 89026 54098 89262 54334
rect 88706 53778 88942 54014
rect 89026 53778 89262 54014
rect 88706 18098 88942 18334
rect 89026 18098 89262 18334
rect 88706 17778 88942 18014
rect 89026 17778 89262 18014
rect 88706 -4422 88942 -4186
rect 89026 -4422 89262 -4186
rect 88706 -4742 88942 -4506
rect 89026 -4742 89262 -4506
rect 92426 273818 92662 274054
rect 92746 273818 92982 274054
rect 92426 273498 92662 273734
rect 92746 273498 92982 273734
rect 92426 237818 92662 238054
rect 92746 237818 92982 238054
rect 92426 237498 92662 237734
rect 92746 237498 92982 237734
rect 92426 201818 92662 202054
rect 92746 201818 92982 202054
rect 92426 201498 92662 201734
rect 92746 201498 92982 201734
rect 92426 165818 92662 166054
rect 92746 165818 92982 166054
rect 92426 165498 92662 165734
rect 92746 165498 92982 165734
rect 92426 129818 92662 130054
rect 92746 129818 92982 130054
rect 92426 129498 92662 129734
rect 92746 129498 92982 129734
rect 92426 93818 92662 94054
rect 92746 93818 92982 94054
rect 92426 93498 92662 93734
rect 92746 93498 92982 93734
rect 92426 57818 92662 58054
rect 92746 57818 92982 58054
rect 92426 57498 92662 57734
rect 92746 57498 92982 57734
rect 92426 21818 92662 22054
rect 92746 21818 92982 22054
rect 92426 21498 92662 21734
rect 92746 21498 92982 21734
rect 92426 -5382 92662 -5146
rect 92746 -5382 92982 -5146
rect 92426 -5702 92662 -5466
rect 92746 -5702 92982 -5466
rect 96146 277538 96382 277774
rect 96466 277538 96702 277774
rect 96146 277218 96382 277454
rect 96466 277218 96702 277454
rect 96146 241538 96382 241774
rect 96466 241538 96702 241774
rect 96146 241218 96382 241454
rect 96466 241218 96702 241454
rect 96146 205538 96382 205774
rect 96466 205538 96702 205774
rect 96146 205218 96382 205454
rect 96466 205218 96702 205454
rect 96146 169538 96382 169774
rect 96466 169538 96702 169774
rect 96146 169218 96382 169454
rect 96466 169218 96702 169454
rect 96146 133538 96382 133774
rect 96466 133538 96702 133774
rect 96146 133218 96382 133454
rect 96466 133218 96702 133454
rect 96146 97538 96382 97774
rect 96466 97538 96702 97774
rect 96146 97218 96382 97454
rect 96466 97218 96702 97454
rect 96146 61538 96382 61774
rect 96466 61538 96702 61774
rect 96146 61218 96382 61454
rect 96466 61218 96702 61454
rect 96146 25538 96382 25774
rect 96466 25538 96702 25774
rect 96146 25218 96382 25454
rect 96466 25218 96702 25454
rect 96146 -6342 96382 -6106
rect 96466 -6342 96702 -6106
rect 96146 -6662 96382 -6426
rect 96466 -6662 96702 -6426
rect 99866 245258 100102 245494
rect 100186 245258 100422 245494
rect 99866 244938 100102 245174
rect 100186 244938 100422 245174
rect 99866 209258 100102 209494
rect 100186 209258 100422 209494
rect 99866 208938 100102 209174
rect 100186 208938 100422 209174
rect 99866 173258 100102 173494
rect 100186 173258 100422 173494
rect 99866 172938 100102 173174
rect 100186 172938 100422 173174
rect 99866 137258 100102 137494
rect 100186 137258 100422 137494
rect 99866 136938 100102 137174
rect 100186 136938 100422 137174
rect 99866 101258 100102 101494
rect 100186 101258 100422 101494
rect 99866 100938 100102 101174
rect 100186 100938 100422 101174
rect 99866 65258 100102 65494
rect 100186 65258 100422 65494
rect 99866 64938 100102 65174
rect 100186 64938 100422 65174
rect 99866 29258 100102 29494
rect 100186 29258 100422 29494
rect 99866 28938 100102 29174
rect 100186 28938 100422 29174
rect 99866 -7302 100102 -7066
rect 100186 -7302 100422 -7066
rect 99866 -7622 100102 -7386
rect 100186 -7622 100422 -7386
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -2502 117502 -2266
rect 117586 -2502 117822 -2266
rect 117266 -2822 117502 -2586
rect 117586 -2822 117822 -2586
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 124706 450098 124942 450334
rect 125026 450098 125262 450334
rect 124706 449778 124942 450014
rect 125026 449778 125262 450014
rect 124706 414098 124942 414334
rect 125026 414098 125262 414334
rect 124706 413778 124942 414014
rect 125026 413778 125262 414014
rect 124706 378098 124942 378334
rect 125026 378098 125262 378334
rect 124706 377778 124942 378014
rect 125026 377778 125262 378014
rect 124706 342098 124942 342334
rect 125026 342098 125262 342334
rect 124706 341778 124942 342014
rect 125026 341778 125262 342014
rect 124706 306098 124942 306334
rect 125026 306098 125262 306334
rect 124706 305778 124942 306014
rect 125026 305778 125262 306014
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 120986 -3462 121222 -3226
rect 121306 -3462 121542 -3226
rect 120986 -3782 121222 -3546
rect 121306 -3782 121542 -3546
rect 124706 270098 124942 270334
rect 125026 270098 125262 270334
rect 124706 269778 124942 270014
rect 125026 269778 125262 270014
rect 124706 234098 124942 234334
rect 125026 234098 125262 234334
rect 124706 233778 124942 234014
rect 125026 233778 125262 234014
rect 124706 198098 124942 198334
rect 125026 198098 125262 198334
rect 124706 197778 124942 198014
rect 125026 197778 125262 198014
rect 124706 162098 124942 162334
rect 125026 162098 125262 162334
rect 124706 161778 124942 162014
rect 125026 161778 125262 162014
rect 124706 126098 124942 126334
rect 125026 126098 125262 126334
rect 124706 125778 124942 126014
rect 125026 125778 125262 126014
rect 124706 90098 124942 90334
rect 125026 90098 125262 90334
rect 124706 89778 124942 90014
rect 125026 89778 125262 90014
rect 124706 54098 124942 54334
rect 125026 54098 125262 54334
rect 124706 53778 124942 54014
rect 125026 53778 125262 54014
rect 124706 18098 124942 18334
rect 125026 18098 125262 18334
rect 124706 17778 124942 18014
rect 125026 17778 125262 18014
rect 124706 -4422 124942 -4186
rect 125026 -4422 125262 -4186
rect 124706 -4742 124942 -4506
rect 125026 -4742 125262 -4506
rect 128426 453818 128662 454054
rect 128746 453818 128982 454054
rect 128426 453498 128662 453734
rect 128746 453498 128982 453734
rect 128426 417818 128662 418054
rect 128746 417818 128982 418054
rect 128426 417498 128662 417734
rect 128746 417498 128982 417734
rect 128426 381818 128662 382054
rect 128746 381818 128982 382054
rect 128426 381498 128662 381734
rect 128746 381498 128982 381734
rect 128426 345818 128662 346054
rect 128746 345818 128982 346054
rect 128426 345498 128662 345734
rect 128746 345498 128982 345734
rect 128426 309818 128662 310054
rect 128746 309818 128982 310054
rect 128426 309498 128662 309734
rect 128746 309498 128982 309734
rect 132146 457538 132382 457774
rect 132466 457538 132702 457774
rect 132146 457218 132382 457454
rect 132466 457218 132702 457454
rect 132146 421538 132382 421774
rect 132466 421538 132702 421774
rect 132146 421218 132382 421454
rect 132466 421218 132702 421454
rect 132146 385538 132382 385774
rect 132466 385538 132702 385774
rect 132146 385218 132382 385454
rect 132466 385218 132702 385454
rect 132146 349538 132382 349774
rect 132466 349538 132702 349774
rect 132146 349218 132382 349454
rect 132466 349218 132702 349454
rect 132146 313538 132382 313774
rect 132466 313538 132702 313774
rect 132146 313218 132382 313454
rect 132466 313218 132702 313454
rect 128426 273818 128662 274054
rect 128746 273818 128982 274054
rect 128426 273498 128662 273734
rect 128746 273498 128982 273734
rect 128426 237818 128662 238054
rect 128746 237818 128982 238054
rect 128426 237498 128662 237734
rect 128746 237498 128982 237734
rect 128426 201818 128662 202054
rect 128746 201818 128982 202054
rect 128426 201498 128662 201734
rect 128746 201498 128982 201734
rect 128426 165818 128662 166054
rect 128746 165818 128982 166054
rect 128426 165498 128662 165734
rect 128746 165498 128982 165734
rect 128426 129818 128662 130054
rect 128746 129818 128982 130054
rect 128426 129498 128662 129734
rect 128746 129498 128982 129734
rect 128426 93818 128662 94054
rect 128746 93818 128982 94054
rect 128426 93498 128662 93734
rect 128746 93498 128982 93734
rect 128426 57818 128662 58054
rect 128746 57818 128982 58054
rect 128426 57498 128662 57734
rect 128746 57498 128982 57734
rect 128426 21818 128662 22054
rect 128746 21818 128982 22054
rect 128426 21498 128662 21734
rect 128746 21498 128982 21734
rect 128426 -5382 128662 -5146
rect 128746 -5382 128982 -5146
rect 128426 -5702 128662 -5466
rect 128746 -5702 128982 -5466
rect 132146 277538 132382 277774
rect 132466 277538 132702 277774
rect 132146 277218 132382 277454
rect 132466 277218 132702 277454
rect 132146 241538 132382 241774
rect 132466 241538 132702 241774
rect 132146 241218 132382 241454
rect 132466 241218 132702 241454
rect 132146 205538 132382 205774
rect 132466 205538 132702 205774
rect 132146 205218 132382 205454
rect 132466 205218 132702 205454
rect 132146 169538 132382 169774
rect 132466 169538 132702 169774
rect 132146 169218 132382 169454
rect 132466 169218 132702 169454
rect 132146 133538 132382 133774
rect 132466 133538 132702 133774
rect 132146 133218 132382 133454
rect 132466 133218 132702 133454
rect 132146 97538 132382 97774
rect 132466 97538 132702 97774
rect 132146 97218 132382 97454
rect 132466 97218 132702 97454
rect 132146 61538 132382 61774
rect 132466 61538 132702 61774
rect 132146 61218 132382 61454
rect 132466 61218 132702 61454
rect 132146 25538 132382 25774
rect 132466 25538 132702 25774
rect 132146 25218 132382 25454
rect 132466 25218 132702 25454
rect 132146 -6342 132382 -6106
rect 132466 -6342 132702 -6106
rect 132146 -6662 132382 -6426
rect 132466 -6662 132702 -6426
rect 135866 461258 136102 461494
rect 136186 461258 136422 461494
rect 135866 460938 136102 461174
rect 136186 460938 136422 461174
rect 135866 425258 136102 425494
rect 136186 425258 136422 425494
rect 135866 424938 136102 425174
rect 136186 424938 136422 425174
rect 135866 389258 136102 389494
rect 136186 389258 136422 389494
rect 135866 388938 136102 389174
rect 136186 388938 136422 389174
rect 135866 353258 136102 353494
rect 136186 353258 136422 353494
rect 135866 352938 136102 353174
rect 136186 352938 136422 353174
rect 135866 317258 136102 317494
rect 136186 317258 136422 317494
rect 135866 316938 136102 317174
rect 136186 316938 136422 317174
rect 135866 281258 136102 281494
rect 136186 281258 136422 281494
rect 135866 280938 136102 281174
rect 136186 280938 136422 281174
rect 135866 245258 136102 245494
rect 136186 245258 136422 245494
rect 135866 244938 136102 245174
rect 136186 244938 136422 245174
rect 135866 209258 136102 209494
rect 136186 209258 136422 209494
rect 135866 208938 136102 209174
rect 136186 208938 136422 209174
rect 135866 173258 136102 173494
rect 136186 173258 136422 173494
rect 135866 172938 136102 173174
rect 136186 172938 136422 173174
rect 135866 137258 136102 137494
rect 136186 137258 136422 137494
rect 135866 136938 136102 137174
rect 136186 136938 136422 137174
rect 135866 101258 136102 101494
rect 136186 101258 136422 101494
rect 135866 100938 136102 101174
rect 136186 100938 136422 101174
rect 135866 65258 136102 65494
rect 136186 65258 136422 65494
rect 135866 64938 136102 65174
rect 136186 64938 136422 65174
rect 135866 29258 136102 29494
rect 136186 29258 136422 29494
rect 135866 28938 136102 29174
rect 136186 28938 136422 29174
rect 135866 -7302 136102 -7066
rect 136186 -7302 136422 -7066
rect 135866 -7622 136102 -7386
rect 136186 -7622 136422 -7386
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -2502 153502 -2266
rect 153586 -2502 153822 -2266
rect 153266 -2822 153502 -2586
rect 153586 -2822 153822 -2586
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 156986 -3462 157222 -3226
rect 157306 -3462 157542 -3226
rect 156986 -3782 157222 -3546
rect 157306 -3782 157542 -3546
rect 160706 450098 160942 450334
rect 161026 450098 161262 450334
rect 160706 449778 160942 450014
rect 161026 449778 161262 450014
rect 160706 414098 160942 414334
rect 161026 414098 161262 414334
rect 160706 413778 160942 414014
rect 161026 413778 161262 414014
rect 160706 378098 160942 378334
rect 161026 378098 161262 378334
rect 160706 377778 160942 378014
rect 161026 377778 161262 378014
rect 160706 342098 160942 342334
rect 161026 342098 161262 342334
rect 160706 341778 160942 342014
rect 161026 341778 161262 342014
rect 160706 306098 160942 306334
rect 161026 306098 161262 306334
rect 160706 305778 160942 306014
rect 161026 305778 161262 306014
rect 164426 453818 164662 454054
rect 164746 453818 164982 454054
rect 164426 453498 164662 453734
rect 164746 453498 164982 453734
rect 164426 417818 164662 418054
rect 164746 417818 164982 418054
rect 164426 417498 164662 417734
rect 164746 417498 164982 417734
rect 164426 381818 164662 382054
rect 164746 381818 164982 382054
rect 164426 381498 164662 381734
rect 164746 381498 164982 381734
rect 164426 345818 164662 346054
rect 164746 345818 164982 346054
rect 164426 345498 164662 345734
rect 164746 345498 164982 345734
rect 164426 309818 164662 310054
rect 164746 309818 164982 310054
rect 164426 309498 164662 309734
rect 164746 309498 164982 309734
rect 160706 270098 160942 270334
rect 161026 270098 161262 270334
rect 160706 269778 160942 270014
rect 161026 269778 161262 270014
rect 160706 234098 160942 234334
rect 161026 234098 161262 234334
rect 160706 233778 160942 234014
rect 161026 233778 161262 234014
rect 160706 198098 160942 198334
rect 161026 198098 161262 198334
rect 160706 197778 160942 198014
rect 161026 197778 161262 198014
rect 160706 162098 160942 162334
rect 161026 162098 161262 162334
rect 160706 161778 160942 162014
rect 161026 161778 161262 162014
rect 160706 126098 160942 126334
rect 161026 126098 161262 126334
rect 160706 125778 160942 126014
rect 161026 125778 161262 126014
rect 160706 90098 160942 90334
rect 161026 90098 161262 90334
rect 160706 89778 160942 90014
rect 161026 89778 161262 90014
rect 160706 54098 160942 54334
rect 161026 54098 161262 54334
rect 160706 53778 160942 54014
rect 161026 53778 161262 54014
rect 160706 18098 160942 18334
rect 161026 18098 161262 18334
rect 160706 17778 160942 18014
rect 161026 17778 161262 18014
rect 160706 -4422 160942 -4186
rect 161026 -4422 161262 -4186
rect 160706 -4742 160942 -4506
rect 161026 -4742 161262 -4506
rect 164426 273818 164662 274054
rect 164746 273818 164982 274054
rect 164426 273498 164662 273734
rect 164746 273498 164982 273734
rect 168146 457538 168382 457774
rect 168466 457538 168702 457774
rect 168146 457218 168382 457454
rect 168466 457218 168702 457454
rect 168146 421538 168382 421774
rect 168466 421538 168702 421774
rect 168146 421218 168382 421454
rect 168466 421218 168702 421454
rect 168146 385538 168382 385774
rect 168466 385538 168702 385774
rect 168146 385218 168382 385454
rect 168466 385218 168702 385454
rect 168146 349538 168382 349774
rect 168466 349538 168702 349774
rect 168146 349218 168382 349454
rect 168466 349218 168702 349454
rect 168146 313538 168382 313774
rect 168466 313538 168702 313774
rect 168146 313218 168382 313454
rect 168466 313218 168702 313454
rect 168146 277538 168382 277774
rect 168466 277538 168702 277774
rect 168146 277218 168382 277454
rect 168466 277218 168702 277454
rect 164426 237818 164662 238054
rect 164746 237818 164982 238054
rect 164426 237498 164662 237734
rect 164746 237498 164982 237734
rect 164426 201818 164662 202054
rect 164746 201818 164982 202054
rect 164426 201498 164662 201734
rect 164746 201498 164982 201734
rect 164426 165818 164662 166054
rect 164746 165818 164982 166054
rect 164426 165498 164662 165734
rect 164746 165498 164982 165734
rect 164426 129818 164662 130054
rect 164746 129818 164982 130054
rect 164426 129498 164662 129734
rect 164746 129498 164982 129734
rect 164426 93818 164662 94054
rect 164746 93818 164982 94054
rect 164426 93498 164662 93734
rect 164746 93498 164982 93734
rect 164426 57818 164662 58054
rect 164746 57818 164982 58054
rect 164426 57498 164662 57734
rect 164746 57498 164982 57734
rect 164426 21818 164662 22054
rect 164746 21818 164982 22054
rect 164426 21498 164662 21734
rect 164746 21498 164982 21734
rect 164426 -5382 164662 -5146
rect 164746 -5382 164982 -5146
rect 164426 -5702 164662 -5466
rect 164746 -5702 164982 -5466
rect 168146 241538 168382 241774
rect 168466 241538 168702 241774
rect 168146 241218 168382 241454
rect 168466 241218 168702 241454
rect 168146 205538 168382 205774
rect 168466 205538 168702 205774
rect 168146 205218 168382 205454
rect 168466 205218 168702 205454
rect 168146 169538 168382 169774
rect 168466 169538 168702 169774
rect 168146 169218 168382 169454
rect 168466 169218 168702 169454
rect 168146 133538 168382 133774
rect 168466 133538 168702 133774
rect 168146 133218 168382 133454
rect 168466 133218 168702 133454
rect 168146 97538 168382 97774
rect 168466 97538 168702 97774
rect 168146 97218 168382 97454
rect 168466 97218 168702 97454
rect 168146 61538 168382 61774
rect 168466 61538 168702 61774
rect 168146 61218 168382 61454
rect 168466 61218 168702 61454
rect 168146 25538 168382 25774
rect 168466 25538 168702 25774
rect 168146 25218 168382 25454
rect 168466 25218 168702 25454
rect 168146 -6342 168382 -6106
rect 168466 -6342 168702 -6106
rect 168146 -6662 168382 -6426
rect 168466 -6662 168702 -6426
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 171866 461258 172102 461494
rect 172186 461258 172422 461494
rect 171866 460938 172102 461174
rect 172186 460938 172422 461174
rect 171866 425258 172102 425494
rect 172186 425258 172422 425494
rect 171866 424938 172102 425174
rect 172186 424938 172422 425174
rect 171866 389258 172102 389494
rect 172186 389258 172422 389494
rect 171866 388938 172102 389174
rect 172186 388938 172422 389174
rect 171866 353258 172102 353494
rect 172186 353258 172422 353494
rect 171866 352938 172102 353174
rect 172186 352938 172422 353174
rect 171866 317258 172102 317494
rect 172186 317258 172422 317494
rect 171866 316938 172102 317174
rect 172186 316938 172422 317174
rect 171866 281258 172102 281494
rect 172186 281258 172422 281494
rect 171866 280938 172102 281174
rect 172186 280938 172422 281174
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 171866 245258 172102 245494
rect 172186 245258 172422 245494
rect 171866 244938 172102 245174
rect 172186 244938 172422 245174
rect 171866 209258 172102 209494
rect 172186 209258 172422 209494
rect 171866 208938 172102 209174
rect 172186 208938 172422 209174
rect 171866 173258 172102 173494
rect 172186 173258 172422 173494
rect 171866 172938 172102 173174
rect 172186 172938 172422 173174
rect 171866 137258 172102 137494
rect 172186 137258 172422 137494
rect 171866 136938 172102 137174
rect 172186 136938 172422 137174
rect 171866 101258 172102 101494
rect 172186 101258 172422 101494
rect 171866 100938 172102 101174
rect 172186 100938 172422 101174
rect 171866 65258 172102 65494
rect 172186 65258 172422 65494
rect 171866 64938 172102 65174
rect 172186 64938 172422 65174
rect 171866 29258 172102 29494
rect 172186 29258 172422 29494
rect 171866 28938 172102 29174
rect 172186 28938 172422 29174
rect 171866 -7302 172102 -7066
rect 172186 -7302 172422 -7066
rect 171866 -7622 172102 -7386
rect 172186 -7622 172422 -7386
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -2502 189502 -2266
rect 189586 -2502 189822 -2266
rect 189266 -2822 189502 -2586
rect 189586 -2822 189822 -2586
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 192986 -3462 193222 -3226
rect 193306 -3462 193542 -3226
rect 192986 -3782 193222 -3546
rect 193306 -3782 193542 -3546
rect 196706 450098 196942 450334
rect 197026 450098 197262 450334
rect 196706 449778 196942 450014
rect 197026 449778 197262 450014
rect 196706 414098 196942 414334
rect 197026 414098 197262 414334
rect 196706 413778 196942 414014
rect 197026 413778 197262 414014
rect 196706 378098 196942 378334
rect 197026 378098 197262 378334
rect 196706 377778 196942 378014
rect 197026 377778 197262 378014
rect 196706 342098 196942 342334
rect 197026 342098 197262 342334
rect 196706 341778 196942 342014
rect 197026 341778 197262 342014
rect 196706 306098 196942 306334
rect 197026 306098 197262 306334
rect 196706 305778 196942 306014
rect 197026 305778 197262 306014
rect 196706 270098 196942 270334
rect 197026 270098 197262 270334
rect 196706 269778 196942 270014
rect 197026 269778 197262 270014
rect 196706 234098 196942 234334
rect 197026 234098 197262 234334
rect 196706 233778 196942 234014
rect 197026 233778 197262 234014
rect 196706 198098 196942 198334
rect 197026 198098 197262 198334
rect 196706 197778 196942 198014
rect 197026 197778 197262 198014
rect 196706 162098 196942 162334
rect 197026 162098 197262 162334
rect 196706 161778 196942 162014
rect 197026 161778 197262 162014
rect 196706 126098 196942 126334
rect 197026 126098 197262 126334
rect 196706 125778 196942 126014
rect 197026 125778 197262 126014
rect 196706 90098 196942 90334
rect 197026 90098 197262 90334
rect 196706 89778 196942 90014
rect 197026 89778 197262 90014
rect 196706 54098 196942 54334
rect 197026 54098 197262 54334
rect 196706 53778 196942 54014
rect 197026 53778 197262 54014
rect 196706 18098 196942 18334
rect 197026 18098 197262 18334
rect 196706 17778 196942 18014
rect 197026 17778 197262 18014
rect 196706 -4422 196942 -4186
rect 197026 -4422 197262 -4186
rect 196706 -4742 196942 -4506
rect 197026 -4742 197262 -4506
rect 200426 453818 200662 454054
rect 200746 453818 200982 454054
rect 200426 453498 200662 453734
rect 200746 453498 200982 453734
rect 200426 417818 200662 418054
rect 200746 417818 200982 418054
rect 200426 417498 200662 417734
rect 200746 417498 200982 417734
rect 200426 381818 200662 382054
rect 200746 381818 200982 382054
rect 200426 381498 200662 381734
rect 200746 381498 200982 381734
rect 200426 345818 200662 346054
rect 200746 345818 200982 346054
rect 200426 345498 200662 345734
rect 200746 345498 200982 345734
rect 200426 309818 200662 310054
rect 200746 309818 200982 310054
rect 200426 309498 200662 309734
rect 200746 309498 200982 309734
rect 200426 273818 200662 274054
rect 200746 273818 200982 274054
rect 200426 273498 200662 273734
rect 200746 273498 200982 273734
rect 204146 457538 204382 457774
rect 204466 457538 204702 457774
rect 204146 457218 204382 457454
rect 204466 457218 204702 457454
rect 204146 421538 204382 421774
rect 204466 421538 204702 421774
rect 204146 421218 204382 421454
rect 204466 421218 204702 421454
rect 204146 385538 204382 385774
rect 204466 385538 204702 385774
rect 204146 385218 204382 385454
rect 204466 385218 204702 385454
rect 204146 349538 204382 349774
rect 204466 349538 204702 349774
rect 204146 349218 204382 349454
rect 204466 349218 204702 349454
rect 204146 313538 204382 313774
rect 204466 313538 204702 313774
rect 204146 313218 204382 313454
rect 204466 313218 204702 313454
rect 204146 277538 204382 277774
rect 204466 277538 204702 277774
rect 204146 277218 204382 277454
rect 204466 277218 204702 277454
rect 200426 237818 200662 238054
rect 200746 237818 200982 238054
rect 200426 237498 200662 237734
rect 200746 237498 200982 237734
rect 200426 201818 200662 202054
rect 200746 201818 200982 202054
rect 200426 201498 200662 201734
rect 200746 201498 200982 201734
rect 200426 165818 200662 166054
rect 200746 165818 200982 166054
rect 200426 165498 200662 165734
rect 200746 165498 200982 165734
rect 200426 129818 200662 130054
rect 200746 129818 200982 130054
rect 200426 129498 200662 129734
rect 200746 129498 200982 129734
rect 200426 93818 200662 94054
rect 200746 93818 200982 94054
rect 200426 93498 200662 93734
rect 200746 93498 200982 93734
rect 200426 57818 200662 58054
rect 200746 57818 200982 58054
rect 200426 57498 200662 57734
rect 200746 57498 200982 57734
rect 200426 21818 200662 22054
rect 200746 21818 200982 22054
rect 200426 21498 200662 21734
rect 200746 21498 200982 21734
rect 200426 -5382 200662 -5146
rect 200746 -5382 200982 -5146
rect 200426 -5702 200662 -5466
rect 200746 -5702 200982 -5466
rect 204146 241538 204382 241774
rect 204466 241538 204702 241774
rect 204146 241218 204382 241454
rect 204466 241218 204702 241454
rect 204146 205538 204382 205774
rect 204466 205538 204702 205774
rect 204146 205218 204382 205454
rect 204466 205218 204702 205454
rect 204146 169538 204382 169774
rect 204466 169538 204702 169774
rect 204146 169218 204382 169454
rect 204466 169218 204702 169454
rect 204146 133538 204382 133774
rect 204466 133538 204702 133774
rect 204146 133218 204382 133454
rect 204466 133218 204702 133454
rect 204146 97538 204382 97774
rect 204466 97538 204702 97774
rect 204146 97218 204382 97454
rect 204466 97218 204702 97454
rect 204146 61538 204382 61774
rect 204466 61538 204702 61774
rect 204146 61218 204382 61454
rect 204466 61218 204702 61454
rect 204146 25538 204382 25774
rect 204466 25538 204702 25774
rect 204146 25218 204382 25454
rect 204466 25218 204702 25454
rect 204146 -6342 204382 -6106
rect 204466 -6342 204702 -6106
rect 204146 -6662 204382 -6426
rect 204466 -6662 204702 -6426
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 207866 461258 208102 461494
rect 208186 461258 208422 461494
rect 207866 460938 208102 461174
rect 208186 460938 208422 461174
rect 207866 425258 208102 425494
rect 208186 425258 208422 425494
rect 207866 424938 208102 425174
rect 208186 424938 208422 425174
rect 207866 389258 208102 389494
rect 208186 389258 208422 389494
rect 207866 388938 208102 389174
rect 208186 388938 208422 389174
rect 207866 353258 208102 353494
rect 208186 353258 208422 353494
rect 207866 352938 208102 353174
rect 208186 352938 208422 353174
rect 207866 317258 208102 317494
rect 208186 317258 208422 317494
rect 207866 316938 208102 317174
rect 208186 316938 208422 317174
rect 207866 281258 208102 281494
rect 208186 281258 208422 281494
rect 207866 280938 208102 281174
rect 208186 280938 208422 281174
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 207866 245258 208102 245494
rect 208186 245258 208422 245494
rect 207866 244938 208102 245174
rect 208186 244938 208422 245174
rect 207866 209258 208102 209494
rect 208186 209258 208422 209494
rect 207866 208938 208102 209174
rect 208186 208938 208422 209174
rect 207866 173258 208102 173494
rect 208186 173258 208422 173494
rect 207866 172938 208102 173174
rect 208186 172938 208422 173174
rect 207866 137258 208102 137494
rect 208186 137258 208422 137494
rect 207866 136938 208102 137174
rect 208186 136938 208422 137174
rect 207866 101258 208102 101494
rect 208186 101258 208422 101494
rect 207866 100938 208102 101174
rect 208186 100938 208422 101174
rect 207866 65258 208102 65494
rect 208186 65258 208422 65494
rect 207866 64938 208102 65174
rect 208186 64938 208422 65174
rect 207866 29258 208102 29494
rect 208186 29258 208422 29494
rect 207866 28938 208102 29174
rect 208186 28938 208422 29174
rect 207866 -7302 208102 -7066
rect 208186 -7302 208422 -7066
rect 207866 -7622 208102 -7386
rect 208186 -7622 208422 -7386
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 225266 -2502 225502 -2266
rect 225586 -2502 225822 -2266
rect 225266 -2822 225502 -2586
rect 225586 -2822 225822 -2586
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 232706 450098 232942 450334
rect 233026 450098 233262 450334
rect 232706 449778 232942 450014
rect 233026 449778 233262 450014
rect 232706 414098 232942 414334
rect 233026 414098 233262 414334
rect 232706 413778 232942 414014
rect 233026 413778 233262 414014
rect 232706 378098 232942 378334
rect 233026 378098 233262 378334
rect 232706 377778 232942 378014
rect 233026 377778 233262 378014
rect 232706 342098 232942 342334
rect 233026 342098 233262 342334
rect 232706 341778 232942 342014
rect 233026 341778 233262 342014
rect 232706 306098 232942 306334
rect 233026 306098 233262 306334
rect 232706 305778 232942 306014
rect 233026 305778 233262 306014
rect 232706 270098 232942 270334
rect 233026 270098 233262 270334
rect 232706 269778 232942 270014
rect 233026 269778 233262 270014
rect 232706 234098 232942 234334
rect 233026 234098 233262 234334
rect 232706 233778 232942 234014
rect 233026 233778 233262 234014
rect 232706 198098 232942 198334
rect 233026 198098 233262 198334
rect 232706 197778 232942 198014
rect 233026 197778 233262 198014
rect 232706 162098 232942 162334
rect 233026 162098 233262 162334
rect 232706 161778 232942 162014
rect 233026 161778 233262 162014
rect 236426 453818 236662 454054
rect 236746 453818 236982 454054
rect 236426 453498 236662 453734
rect 236746 453498 236982 453734
rect 236426 417818 236662 418054
rect 236746 417818 236982 418054
rect 236426 417498 236662 417734
rect 236746 417498 236982 417734
rect 236426 381818 236662 382054
rect 236746 381818 236982 382054
rect 236426 381498 236662 381734
rect 236746 381498 236982 381734
rect 236426 345818 236662 346054
rect 236746 345818 236982 346054
rect 236426 345498 236662 345734
rect 236746 345498 236982 345734
rect 236426 309818 236662 310054
rect 236746 309818 236982 310054
rect 236426 309498 236662 309734
rect 236746 309498 236982 309734
rect 240146 457538 240382 457774
rect 240466 457538 240702 457774
rect 240146 457218 240382 457454
rect 240466 457218 240702 457454
rect 240146 421538 240382 421774
rect 240466 421538 240702 421774
rect 240146 421218 240382 421454
rect 240466 421218 240702 421454
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 244250 435218 244486 435454
rect 244250 434898 244486 435134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 259610 402938 259846 403174
rect 259610 402618 259846 402854
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 268706 450098 268942 450334
rect 269026 450098 269262 450334
rect 268706 449778 268942 450014
rect 269026 449778 269262 450014
rect 268706 414098 268942 414334
rect 269026 414098 269262 414334
rect 268706 413778 268942 414014
rect 269026 413778 269262 414014
rect 272426 453818 272662 454054
rect 272746 453818 272982 454054
rect 272426 453498 272662 453734
rect 272746 453498 272982 453734
rect 276146 457538 276382 457774
rect 276466 457538 276702 457774
rect 276146 457218 276382 457454
rect 276466 457218 276702 457454
rect 274970 435218 275206 435454
rect 274970 434898 275206 435134
rect 272426 417818 272662 418054
rect 272746 417818 272982 418054
rect 272426 417498 272662 417734
rect 272746 417498 272982 417734
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 279866 461258 280102 461494
rect 280186 461258 280422 461494
rect 279866 460938 280102 461174
rect 280186 460938 280422 461174
rect 276146 421538 276382 421774
rect 276466 421538 276702 421774
rect 276146 421218 276382 421454
rect 276466 421218 276702 421454
rect 244250 399218 244486 399454
rect 244250 398898 244486 399134
rect 274970 399218 275206 399454
rect 274970 398898 275206 399134
rect 279866 425258 280102 425494
rect 280186 425258 280422 425494
rect 279866 424938 280102 425174
rect 280186 424938 280422 425174
rect 279866 389258 280102 389494
rect 280186 389258 280422 389494
rect 279866 388938 280102 389174
rect 280186 388938 280422 389174
rect 259610 366938 259846 367174
rect 259610 366618 259846 366854
rect 244250 363218 244486 363454
rect 244250 362898 244486 363134
rect 274970 363218 275206 363454
rect 274970 362898 275206 363134
rect 279866 353258 280102 353494
rect 280186 353258 280422 353494
rect 279866 352938 280102 353174
rect 280186 352938 280422 353174
rect 259610 330938 259846 331174
rect 259610 330618 259846 330854
rect 244250 327218 244486 327454
rect 244250 326898 244486 327134
rect 274970 327218 275206 327454
rect 274970 326898 275206 327134
rect 279866 317258 280102 317494
rect 280186 317258 280422 317494
rect 279866 316938 280102 317174
rect 280186 316938 280422 317174
rect 259610 294938 259846 295174
rect 259610 294618 259846 294854
rect 236426 273818 236662 274054
rect 236746 273818 236982 274054
rect 236426 273498 236662 273734
rect 236746 273498 236982 273734
rect 236426 237818 236662 238054
rect 236746 237818 236982 238054
rect 236426 237498 236662 237734
rect 236746 237498 236982 237734
rect 244250 291218 244486 291454
rect 236426 201818 236662 202054
rect 236746 201818 236982 202054
rect 236426 201498 236662 201734
rect 236746 201498 236982 201734
rect 244250 290898 244486 291134
rect 274970 291218 275206 291454
rect 274970 290898 275206 291134
rect 236426 165818 236662 166054
rect 236746 165818 236982 166054
rect 236426 165498 236662 165734
rect 236746 165498 236982 165734
rect 232706 126098 232942 126334
rect 233026 126098 233262 126334
rect 232706 125778 232942 126014
rect 233026 125778 233262 126014
rect 232706 90098 232942 90334
rect 233026 90098 233262 90334
rect 232706 89778 232942 90014
rect 233026 89778 233262 90014
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 228986 -3462 229222 -3226
rect 229306 -3462 229542 -3226
rect 228986 -3782 229222 -3546
rect 229306 -3782 229542 -3546
rect 232706 54098 232942 54334
rect 233026 54098 233262 54334
rect 232706 53778 232942 54014
rect 233026 53778 233262 54014
rect 232706 18098 232942 18334
rect 233026 18098 233262 18334
rect 232706 17778 232942 18014
rect 233026 17778 233262 18014
rect 232706 -4422 232942 -4186
rect 233026 -4422 233262 -4186
rect 232706 -4742 232942 -4506
rect 233026 -4742 233262 -4506
rect 236426 129818 236662 130054
rect 236746 129818 236982 130054
rect 236426 129498 236662 129734
rect 236746 129498 236982 129734
rect 259610 258938 259846 259174
rect 259610 258618 259846 258854
rect 244250 255218 244486 255454
rect 244250 254898 244486 255134
rect 274970 255218 275206 255454
rect 274970 254898 275206 255134
rect 240146 205538 240382 205774
rect 240466 205538 240702 205774
rect 240146 205218 240382 205454
rect 240466 205218 240702 205454
rect 240146 169538 240382 169774
rect 240466 169538 240702 169774
rect 240146 169218 240382 169454
rect 240466 169218 240702 169454
rect 240146 133538 240382 133774
rect 240466 133538 240702 133774
rect 240146 133218 240382 133454
rect 240466 133218 240702 133454
rect 236426 93818 236662 94054
rect 236746 93818 236982 94054
rect 236426 93498 236662 93734
rect 236746 93498 236982 93734
rect 236426 57818 236662 58054
rect 236746 57818 236982 58054
rect 236426 57498 236662 57734
rect 236746 57498 236982 57734
rect 236426 21818 236662 22054
rect 236746 21818 236982 22054
rect 236426 21498 236662 21734
rect 236746 21498 236982 21734
rect 236426 -5382 236662 -5146
rect 236746 -5382 236982 -5146
rect 236426 -5702 236662 -5466
rect 236746 -5702 236982 -5466
rect 240146 97538 240382 97774
rect 240466 97538 240702 97774
rect 240146 97218 240382 97454
rect 240466 97218 240702 97454
rect 240146 61538 240382 61774
rect 240466 61538 240702 61774
rect 240146 61218 240382 61454
rect 240466 61218 240702 61454
rect 240146 25538 240382 25774
rect 240466 25538 240702 25774
rect 240146 25218 240382 25454
rect 240466 25218 240702 25454
rect 240146 -6342 240382 -6106
rect 240466 -6342 240702 -6106
rect 240146 -6662 240382 -6426
rect 240466 -6662 240702 -6426
rect 243866 209258 244102 209494
rect 244186 209258 244422 209494
rect 243866 208938 244102 209174
rect 244186 208938 244422 209174
rect 243866 173258 244102 173494
rect 244186 173258 244422 173494
rect 243866 172938 244102 173174
rect 244186 172938 244422 173174
rect 243866 137258 244102 137494
rect 244186 137258 244422 137494
rect 243866 136938 244102 137174
rect 244186 136938 244422 137174
rect 243866 101258 244102 101494
rect 244186 101258 244422 101494
rect 243866 100938 244102 101174
rect 244186 100938 244422 101174
rect 243866 65258 244102 65494
rect 244186 65258 244422 65494
rect 243866 64938 244102 65174
rect 244186 64938 244422 65174
rect 243866 29258 244102 29494
rect 244186 29258 244422 29494
rect 243866 28938 244102 29174
rect 244186 28938 244422 29174
rect 243866 -7302 244102 -7066
rect 244186 -7302 244422 -7066
rect 243866 -7622 244102 -7386
rect 244186 -7622 244422 -7386
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -2502 261502 -2266
rect 261586 -2502 261822 -2266
rect 261266 -2822 261502 -2586
rect 261586 -2822 261822 -2586
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 264986 -3462 265222 -3226
rect 265306 -3462 265542 -3226
rect 264986 -3782 265222 -3546
rect 265306 -3782 265542 -3546
rect 268706 234098 268942 234334
rect 269026 234098 269262 234334
rect 268706 233778 268942 234014
rect 269026 233778 269262 234014
rect 268706 198098 268942 198334
rect 269026 198098 269262 198334
rect 268706 197778 268942 198014
rect 269026 197778 269262 198014
rect 268706 162098 268942 162334
rect 269026 162098 269262 162334
rect 268706 161778 268942 162014
rect 269026 161778 269262 162014
rect 268706 126098 268942 126334
rect 269026 126098 269262 126334
rect 268706 125778 268942 126014
rect 269026 125778 269262 126014
rect 268706 90098 268942 90334
rect 269026 90098 269262 90334
rect 268706 89778 268942 90014
rect 269026 89778 269262 90014
rect 268706 54098 268942 54334
rect 269026 54098 269262 54334
rect 268706 53778 268942 54014
rect 269026 53778 269262 54014
rect 268706 18098 268942 18334
rect 269026 18098 269262 18334
rect 268706 17778 268942 18014
rect 269026 17778 269262 18014
rect 268706 -4422 268942 -4186
rect 269026 -4422 269262 -4186
rect 268706 -4742 268942 -4506
rect 269026 -4742 269262 -4506
rect 272426 237818 272662 238054
rect 272746 237818 272982 238054
rect 272426 237498 272662 237734
rect 272746 237498 272982 237734
rect 272426 201818 272662 202054
rect 272746 201818 272982 202054
rect 272426 201498 272662 201734
rect 272746 201498 272982 201734
rect 272426 165818 272662 166054
rect 272746 165818 272982 166054
rect 272426 165498 272662 165734
rect 272746 165498 272982 165734
rect 272426 129818 272662 130054
rect 272746 129818 272982 130054
rect 272426 129498 272662 129734
rect 272746 129498 272982 129734
rect 272426 93818 272662 94054
rect 272746 93818 272982 94054
rect 272426 93498 272662 93734
rect 272746 93498 272982 93734
rect 272426 57818 272662 58054
rect 272746 57818 272982 58054
rect 272426 57498 272662 57734
rect 272746 57498 272982 57734
rect 272426 21818 272662 22054
rect 272746 21818 272982 22054
rect 272426 21498 272662 21734
rect 272746 21498 272982 21734
rect 272426 -5382 272662 -5146
rect 272746 -5382 272982 -5146
rect 272426 -5702 272662 -5466
rect 272746 -5702 272982 -5466
rect 279866 281258 280102 281494
rect 280186 281258 280422 281494
rect 279866 280938 280102 281174
rect 280186 280938 280422 281174
rect 279866 245258 280102 245494
rect 280186 245258 280422 245494
rect 279866 244938 280102 245174
rect 280186 244938 280422 245174
rect 276146 205538 276382 205774
rect 276466 205538 276702 205774
rect 276146 205218 276382 205454
rect 276466 205218 276702 205454
rect 276146 169538 276382 169774
rect 276466 169538 276702 169774
rect 276146 169218 276382 169454
rect 276466 169218 276702 169454
rect 276146 133538 276382 133774
rect 276466 133538 276702 133774
rect 276146 133218 276382 133454
rect 276466 133218 276702 133454
rect 276146 97538 276382 97774
rect 276466 97538 276702 97774
rect 276146 97218 276382 97454
rect 276466 97218 276702 97454
rect 276146 61538 276382 61774
rect 276466 61538 276702 61774
rect 276146 61218 276382 61454
rect 276466 61218 276702 61454
rect 276146 25538 276382 25774
rect 276466 25538 276702 25774
rect 276146 25218 276382 25454
rect 276466 25218 276702 25454
rect 276146 -6342 276382 -6106
rect 276466 -6342 276702 -6106
rect 276146 -6662 276382 -6426
rect 276466 -6662 276702 -6426
rect 279866 209258 280102 209494
rect 280186 209258 280422 209494
rect 279866 208938 280102 209174
rect 280186 208938 280422 209174
rect 279866 173258 280102 173494
rect 280186 173258 280422 173494
rect 279866 172938 280102 173174
rect 280186 172938 280422 173174
rect 279866 137258 280102 137494
rect 280186 137258 280422 137494
rect 279866 136938 280102 137174
rect 280186 136938 280422 137174
rect 279866 101258 280102 101494
rect 280186 101258 280422 101494
rect 279866 100938 280102 101174
rect 280186 100938 280422 101174
rect 279866 65258 280102 65494
rect 280186 65258 280422 65494
rect 279866 64938 280102 65174
rect 280186 64938 280422 65174
rect 279866 29258 280102 29494
rect 280186 29258 280422 29494
rect 279866 28938 280102 29174
rect 280186 28938 280422 29174
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 279866 -7302 280102 -7066
rect 280186 -7302 280422 -7066
rect 279866 -7622 280102 -7386
rect 280186 -7622 280422 -7386
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 297266 706522 297502 706758
rect 297586 706522 297822 706758
rect 297266 706202 297502 706438
rect 297586 706202 297822 706438
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 300986 707482 301222 707718
rect 301306 707482 301542 707718
rect 300986 707162 301222 707398
rect 301306 707162 301542 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -2502 297502 -2266
rect 297586 -2502 297822 -2266
rect 297266 -2822 297502 -2586
rect 297586 -2822 297822 -2586
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 300986 -3462 301222 -3226
rect 301306 -3462 301542 -3226
rect 300986 -3782 301222 -3546
rect 301306 -3782 301542 -3546
rect 304706 708442 304942 708678
rect 305026 708442 305262 708678
rect 304706 708122 304942 708358
rect 305026 708122 305262 708358
rect 304706 666098 304942 666334
rect 305026 666098 305262 666334
rect 304706 665778 304942 666014
rect 305026 665778 305262 666014
rect 304706 630098 304942 630334
rect 305026 630098 305262 630334
rect 304706 629778 304942 630014
rect 305026 629778 305262 630014
rect 304706 594098 304942 594334
rect 305026 594098 305262 594334
rect 304706 593778 304942 594014
rect 305026 593778 305262 594014
rect 308426 709402 308662 709638
rect 308746 709402 308982 709638
rect 308426 709082 308662 709318
rect 308746 709082 308982 709318
rect 308426 669818 308662 670054
rect 308746 669818 308982 670054
rect 308426 669498 308662 669734
rect 308746 669498 308982 669734
rect 308426 633818 308662 634054
rect 308746 633818 308982 634054
rect 308426 633498 308662 633734
rect 308746 633498 308982 633734
rect 308426 597818 308662 598054
rect 308746 597818 308982 598054
rect 308426 597498 308662 597734
rect 308746 597498 308982 597734
rect 304706 558098 304942 558334
rect 305026 558098 305262 558334
rect 304706 557778 304942 558014
rect 305026 557778 305262 558014
rect 304706 522098 304942 522334
rect 305026 522098 305262 522334
rect 304706 521778 304942 522014
rect 305026 521778 305262 522014
rect 304706 486098 304942 486334
rect 305026 486098 305262 486334
rect 304706 485778 304942 486014
rect 305026 485778 305262 486014
rect 304706 450098 304942 450334
rect 305026 450098 305262 450334
rect 304706 449778 304942 450014
rect 305026 449778 305262 450014
rect 304706 414098 304942 414334
rect 305026 414098 305262 414334
rect 304706 413778 304942 414014
rect 305026 413778 305262 414014
rect 304706 378098 304942 378334
rect 305026 378098 305262 378334
rect 304706 377778 304942 378014
rect 305026 377778 305262 378014
rect 304706 342098 304942 342334
rect 305026 342098 305262 342334
rect 304706 341778 304942 342014
rect 305026 341778 305262 342014
rect 304706 306098 304942 306334
rect 305026 306098 305262 306334
rect 304706 305778 304942 306014
rect 305026 305778 305262 306014
rect 304706 270098 304942 270334
rect 305026 270098 305262 270334
rect 304706 269778 304942 270014
rect 305026 269778 305262 270014
rect 308426 561818 308662 562054
rect 308746 561818 308982 562054
rect 308426 561498 308662 561734
rect 308746 561498 308982 561734
rect 308426 525818 308662 526054
rect 308746 525818 308982 526054
rect 308426 525498 308662 525734
rect 308746 525498 308982 525734
rect 312146 710362 312382 710598
rect 312466 710362 312702 710598
rect 312146 710042 312382 710278
rect 312466 710042 312702 710278
rect 312146 673538 312382 673774
rect 312466 673538 312702 673774
rect 312146 673218 312382 673454
rect 312466 673218 312702 673454
rect 312146 637538 312382 637774
rect 312466 637538 312702 637774
rect 312146 637218 312382 637454
rect 312466 637218 312702 637454
rect 312146 601538 312382 601774
rect 312466 601538 312702 601774
rect 312146 601218 312382 601454
rect 312466 601218 312702 601454
rect 315866 711322 316102 711558
rect 316186 711322 316422 711558
rect 315866 711002 316102 711238
rect 316186 711002 316422 711238
rect 315866 677258 316102 677494
rect 316186 677258 316422 677494
rect 315866 676938 316102 677174
rect 316186 676938 316422 677174
rect 315866 641258 316102 641494
rect 316186 641258 316422 641494
rect 315866 640938 316102 641174
rect 316186 640938 316422 641174
rect 315866 605258 316102 605494
rect 316186 605258 316422 605494
rect 315866 604938 316102 605174
rect 316186 604938 316422 605174
rect 312146 565538 312382 565774
rect 312466 565538 312702 565774
rect 312146 565218 312382 565454
rect 312466 565218 312702 565454
rect 312146 529538 312382 529774
rect 312466 529538 312702 529774
rect 312146 529218 312382 529454
rect 312466 529218 312702 529454
rect 308426 489818 308662 490054
rect 308746 489818 308982 490054
rect 308426 489498 308662 489734
rect 308746 489498 308982 489734
rect 308426 453818 308662 454054
rect 308746 453818 308982 454054
rect 308426 453498 308662 453734
rect 308746 453498 308982 453734
rect 308426 417818 308662 418054
rect 308746 417818 308982 418054
rect 308426 417498 308662 417734
rect 308746 417498 308982 417734
rect 308426 381818 308662 382054
rect 308746 381818 308982 382054
rect 308426 381498 308662 381734
rect 308746 381498 308982 381734
rect 308426 345818 308662 346054
rect 308746 345818 308982 346054
rect 308426 345498 308662 345734
rect 308746 345498 308982 345734
rect 308426 309818 308662 310054
rect 308746 309818 308982 310054
rect 308426 309498 308662 309734
rect 308746 309498 308982 309734
rect 308426 273818 308662 274054
rect 308746 273818 308982 274054
rect 308426 273498 308662 273734
rect 308746 273498 308982 273734
rect 304706 234098 304942 234334
rect 305026 234098 305262 234334
rect 304706 233778 304942 234014
rect 305026 233778 305262 234014
rect 304706 198098 304942 198334
rect 305026 198098 305262 198334
rect 304706 197778 304942 198014
rect 305026 197778 305262 198014
rect 304706 162098 304942 162334
rect 305026 162098 305262 162334
rect 304706 161778 304942 162014
rect 305026 161778 305262 162014
rect 304706 126098 304942 126334
rect 305026 126098 305262 126334
rect 304706 125778 304942 126014
rect 305026 125778 305262 126014
rect 304706 90098 304942 90334
rect 305026 90098 305262 90334
rect 304706 89778 304942 90014
rect 305026 89778 305262 90014
rect 304706 54098 304942 54334
rect 305026 54098 305262 54334
rect 304706 53778 304942 54014
rect 305026 53778 305262 54014
rect 304706 18098 304942 18334
rect 305026 18098 305262 18334
rect 304706 17778 304942 18014
rect 305026 17778 305262 18014
rect 304706 -4422 304942 -4186
rect 305026 -4422 305262 -4186
rect 304706 -4742 304942 -4506
rect 305026 -4742 305262 -4506
rect 312146 493538 312382 493774
rect 312466 493538 312702 493774
rect 312146 493218 312382 493454
rect 312466 493218 312702 493454
rect 312146 457538 312382 457774
rect 312466 457538 312702 457774
rect 312146 457218 312382 457454
rect 312466 457218 312702 457454
rect 312146 421538 312382 421774
rect 312466 421538 312702 421774
rect 312146 421218 312382 421454
rect 312466 421218 312702 421454
rect 312146 385538 312382 385774
rect 312466 385538 312702 385774
rect 312146 385218 312382 385454
rect 312466 385218 312702 385454
rect 312146 349538 312382 349774
rect 312466 349538 312702 349774
rect 312146 349218 312382 349454
rect 312466 349218 312702 349454
rect 312146 313538 312382 313774
rect 312466 313538 312702 313774
rect 312146 313218 312382 313454
rect 312466 313218 312702 313454
rect 312146 277538 312382 277774
rect 312466 277538 312702 277774
rect 312146 277218 312382 277454
rect 312466 277218 312702 277454
rect 308426 237818 308662 238054
rect 308746 237818 308982 238054
rect 308426 237498 308662 237734
rect 308746 237498 308982 237734
rect 308426 201818 308662 202054
rect 308746 201818 308982 202054
rect 308426 201498 308662 201734
rect 308746 201498 308982 201734
rect 308426 165818 308662 166054
rect 308746 165818 308982 166054
rect 308426 165498 308662 165734
rect 308746 165498 308982 165734
rect 308426 129818 308662 130054
rect 308746 129818 308982 130054
rect 308426 129498 308662 129734
rect 308746 129498 308982 129734
rect 308426 93818 308662 94054
rect 308746 93818 308982 94054
rect 308426 93498 308662 93734
rect 308746 93498 308982 93734
rect 308426 57818 308662 58054
rect 308746 57818 308982 58054
rect 308426 57498 308662 57734
rect 308746 57498 308982 57734
rect 308426 21818 308662 22054
rect 308746 21818 308982 22054
rect 308426 21498 308662 21734
rect 308746 21498 308982 21734
rect 308426 -5382 308662 -5146
rect 308746 -5382 308982 -5146
rect 308426 -5702 308662 -5466
rect 308746 -5702 308982 -5466
rect 315866 569258 316102 569494
rect 316186 569258 316422 569494
rect 315866 568938 316102 569174
rect 316186 568938 316422 569174
rect 315866 533258 316102 533494
rect 316186 533258 316422 533494
rect 315866 532938 316102 533174
rect 316186 532938 316422 533174
rect 315866 497258 316102 497494
rect 316186 497258 316422 497494
rect 315866 496938 316102 497174
rect 316186 496938 316422 497174
rect 315866 461258 316102 461494
rect 316186 461258 316422 461494
rect 315866 460938 316102 461174
rect 316186 460938 316422 461174
rect 315866 425258 316102 425494
rect 316186 425258 316422 425494
rect 315866 424938 316102 425174
rect 316186 424938 316422 425174
rect 315866 389258 316102 389494
rect 316186 389258 316422 389494
rect 315866 388938 316102 389174
rect 316186 388938 316422 389174
rect 315866 353258 316102 353494
rect 316186 353258 316422 353494
rect 315866 352938 316102 353174
rect 316186 352938 316422 353174
rect 315866 317258 316102 317494
rect 316186 317258 316422 317494
rect 315866 316938 316102 317174
rect 316186 316938 316422 317174
rect 315866 281258 316102 281494
rect 316186 281258 316422 281494
rect 315866 280938 316102 281174
rect 316186 280938 316422 281174
rect 312146 241538 312382 241774
rect 312466 241538 312702 241774
rect 312146 241218 312382 241454
rect 312466 241218 312702 241454
rect 312146 205538 312382 205774
rect 312466 205538 312702 205774
rect 312146 205218 312382 205454
rect 312466 205218 312702 205454
rect 312146 169538 312382 169774
rect 312466 169538 312702 169774
rect 312146 169218 312382 169454
rect 312466 169218 312702 169454
rect 312146 133538 312382 133774
rect 312466 133538 312702 133774
rect 312146 133218 312382 133454
rect 312466 133218 312702 133454
rect 312146 97538 312382 97774
rect 312466 97538 312702 97774
rect 312146 97218 312382 97454
rect 312466 97218 312702 97454
rect 312146 61538 312382 61774
rect 312466 61538 312702 61774
rect 312146 61218 312382 61454
rect 312466 61218 312702 61454
rect 312146 25538 312382 25774
rect 312466 25538 312702 25774
rect 312146 25218 312382 25454
rect 312466 25218 312702 25454
rect 312146 -6342 312382 -6106
rect 312466 -6342 312702 -6106
rect 312146 -6662 312382 -6426
rect 312466 -6662 312702 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 315866 245258 316102 245494
rect 316186 245258 316422 245494
rect 315866 244938 316102 245174
rect 316186 244938 316422 245174
rect 315866 209258 316102 209494
rect 316186 209258 316422 209494
rect 315866 208938 316102 209174
rect 316186 208938 316422 209174
rect 315866 173258 316102 173494
rect 316186 173258 316422 173494
rect 315866 172938 316102 173174
rect 316186 172938 316422 173174
rect 315866 137258 316102 137494
rect 316186 137258 316422 137494
rect 315866 136938 316102 137174
rect 316186 136938 316422 137174
rect 315866 101258 316102 101494
rect 316186 101258 316422 101494
rect 315866 100938 316102 101174
rect 316186 100938 316422 101174
rect 315866 65258 316102 65494
rect 316186 65258 316422 65494
rect 315866 64938 316102 65174
rect 316186 64938 316422 65174
rect 315866 29258 316102 29494
rect 316186 29258 316422 29494
rect 315866 28938 316102 29174
rect 316186 28938 316422 29174
rect 315866 -7302 316102 -7066
rect 316186 -7302 316422 -7066
rect 315866 -7622 316102 -7386
rect 316186 -7622 316422 -7386
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 333266 706522 333502 706758
rect 333586 706522 333822 706758
rect 333266 706202 333502 706438
rect 333586 706202 333822 706438
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -2502 333502 -2266
rect 333586 -2502 333822 -2266
rect 333266 -2822 333502 -2586
rect 333586 -2822 333822 -2586
rect 336986 707482 337222 707718
rect 337306 707482 337542 707718
rect 336986 707162 337222 707398
rect 337306 707162 337542 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 336986 -3462 337222 -3226
rect 337306 -3462 337542 -3226
rect 336986 -3782 337222 -3546
rect 337306 -3782 337542 -3546
rect 340706 708442 340942 708678
rect 341026 708442 341262 708678
rect 340706 708122 340942 708358
rect 341026 708122 341262 708358
rect 340706 666098 340942 666334
rect 341026 666098 341262 666334
rect 340706 665778 340942 666014
rect 341026 665778 341262 666014
rect 340706 630098 340942 630334
rect 341026 630098 341262 630334
rect 340706 629778 340942 630014
rect 341026 629778 341262 630014
rect 340706 594098 340942 594334
rect 341026 594098 341262 594334
rect 340706 593778 340942 594014
rect 341026 593778 341262 594014
rect 340706 558098 340942 558334
rect 341026 558098 341262 558334
rect 340706 557778 340942 558014
rect 341026 557778 341262 558014
rect 340706 522098 340942 522334
rect 341026 522098 341262 522334
rect 340706 521778 340942 522014
rect 341026 521778 341262 522014
rect 340706 486098 340942 486334
rect 341026 486098 341262 486334
rect 340706 485778 340942 486014
rect 341026 485778 341262 486014
rect 340706 450098 340942 450334
rect 341026 450098 341262 450334
rect 340706 449778 340942 450014
rect 341026 449778 341262 450014
rect 340706 414098 340942 414334
rect 341026 414098 341262 414334
rect 340706 413778 340942 414014
rect 341026 413778 341262 414014
rect 340706 378098 340942 378334
rect 341026 378098 341262 378334
rect 340706 377778 340942 378014
rect 341026 377778 341262 378014
rect 340706 342098 340942 342334
rect 341026 342098 341262 342334
rect 340706 341778 340942 342014
rect 341026 341778 341262 342014
rect 340706 306098 340942 306334
rect 341026 306098 341262 306334
rect 340706 305778 340942 306014
rect 341026 305778 341262 306014
rect 340706 270098 340942 270334
rect 341026 270098 341262 270334
rect 340706 269778 340942 270014
rect 341026 269778 341262 270014
rect 340706 234098 340942 234334
rect 341026 234098 341262 234334
rect 340706 233778 340942 234014
rect 341026 233778 341262 234014
rect 340706 198098 340942 198334
rect 341026 198098 341262 198334
rect 340706 197778 340942 198014
rect 341026 197778 341262 198014
rect 340706 162098 340942 162334
rect 341026 162098 341262 162334
rect 340706 161778 340942 162014
rect 341026 161778 341262 162014
rect 340706 126098 340942 126334
rect 341026 126098 341262 126334
rect 340706 125778 340942 126014
rect 341026 125778 341262 126014
rect 340706 90098 340942 90334
rect 341026 90098 341262 90334
rect 340706 89778 340942 90014
rect 341026 89778 341262 90014
rect 340706 54098 340942 54334
rect 341026 54098 341262 54334
rect 340706 53778 340942 54014
rect 341026 53778 341262 54014
rect 340706 18098 340942 18334
rect 341026 18098 341262 18334
rect 340706 17778 340942 18014
rect 341026 17778 341262 18014
rect 340706 -4422 340942 -4186
rect 341026 -4422 341262 -4186
rect 340706 -4742 340942 -4506
rect 341026 -4742 341262 -4506
rect 344426 709402 344662 709638
rect 344746 709402 344982 709638
rect 344426 709082 344662 709318
rect 344746 709082 344982 709318
rect 344426 669818 344662 670054
rect 344746 669818 344982 670054
rect 344426 669498 344662 669734
rect 344746 669498 344982 669734
rect 344426 633818 344662 634054
rect 344746 633818 344982 634054
rect 344426 633498 344662 633734
rect 344746 633498 344982 633734
rect 344426 597818 344662 598054
rect 344746 597818 344982 598054
rect 344426 597498 344662 597734
rect 344746 597498 344982 597734
rect 344426 561818 344662 562054
rect 344746 561818 344982 562054
rect 344426 561498 344662 561734
rect 344746 561498 344982 561734
rect 344426 525818 344662 526054
rect 344746 525818 344982 526054
rect 344426 525498 344662 525734
rect 344746 525498 344982 525734
rect 344426 489818 344662 490054
rect 344746 489818 344982 490054
rect 344426 489498 344662 489734
rect 344746 489498 344982 489734
rect 344426 453818 344662 454054
rect 344746 453818 344982 454054
rect 344426 453498 344662 453734
rect 344746 453498 344982 453734
rect 344426 417818 344662 418054
rect 344746 417818 344982 418054
rect 344426 417498 344662 417734
rect 344746 417498 344982 417734
rect 344426 381818 344662 382054
rect 344746 381818 344982 382054
rect 344426 381498 344662 381734
rect 344746 381498 344982 381734
rect 344426 345818 344662 346054
rect 344746 345818 344982 346054
rect 344426 345498 344662 345734
rect 344746 345498 344982 345734
rect 344426 309818 344662 310054
rect 344746 309818 344982 310054
rect 344426 309498 344662 309734
rect 344746 309498 344982 309734
rect 344426 273818 344662 274054
rect 344746 273818 344982 274054
rect 344426 273498 344662 273734
rect 344746 273498 344982 273734
rect 348146 710362 348382 710598
rect 348466 710362 348702 710598
rect 348146 710042 348382 710278
rect 348466 710042 348702 710278
rect 348146 673538 348382 673774
rect 348466 673538 348702 673774
rect 348146 673218 348382 673454
rect 348466 673218 348702 673454
rect 348146 637538 348382 637774
rect 348466 637538 348702 637774
rect 348146 637218 348382 637454
rect 348466 637218 348702 637454
rect 348146 601538 348382 601774
rect 348466 601538 348702 601774
rect 348146 601218 348382 601454
rect 348466 601218 348702 601454
rect 348146 565538 348382 565774
rect 348466 565538 348702 565774
rect 348146 565218 348382 565454
rect 348466 565218 348702 565454
rect 348146 529538 348382 529774
rect 348466 529538 348702 529774
rect 348146 529218 348382 529454
rect 348466 529218 348702 529454
rect 348146 493538 348382 493774
rect 348466 493538 348702 493774
rect 348146 493218 348382 493454
rect 348466 493218 348702 493454
rect 348146 457538 348382 457774
rect 348466 457538 348702 457774
rect 348146 457218 348382 457454
rect 348466 457218 348702 457454
rect 348146 421538 348382 421774
rect 348466 421538 348702 421774
rect 348146 421218 348382 421454
rect 348466 421218 348702 421454
rect 348146 385538 348382 385774
rect 348466 385538 348702 385774
rect 348146 385218 348382 385454
rect 348466 385218 348702 385454
rect 348146 349538 348382 349774
rect 348466 349538 348702 349774
rect 348146 349218 348382 349454
rect 348466 349218 348702 349454
rect 348146 313538 348382 313774
rect 348466 313538 348702 313774
rect 348146 313218 348382 313454
rect 348466 313218 348702 313454
rect 348146 277538 348382 277774
rect 348466 277538 348702 277774
rect 348146 277218 348382 277454
rect 348466 277218 348702 277454
rect 344426 237818 344662 238054
rect 344746 237818 344982 238054
rect 344426 237498 344662 237734
rect 344746 237498 344982 237734
rect 344426 201818 344662 202054
rect 344746 201818 344982 202054
rect 344426 201498 344662 201734
rect 344746 201498 344982 201734
rect 344426 165818 344662 166054
rect 344746 165818 344982 166054
rect 344426 165498 344662 165734
rect 344746 165498 344982 165734
rect 348146 241538 348382 241774
rect 348466 241538 348702 241774
rect 348146 241218 348382 241454
rect 348466 241218 348702 241454
rect 348146 205538 348382 205774
rect 348466 205538 348702 205774
rect 348146 205218 348382 205454
rect 348466 205218 348702 205454
rect 348146 169538 348382 169774
rect 348466 169538 348702 169774
rect 348146 169218 348382 169454
rect 348466 169218 348702 169454
rect 344426 129818 344662 130054
rect 344746 129818 344982 130054
rect 344426 129498 344662 129734
rect 344746 129498 344982 129734
rect 344426 93818 344662 94054
rect 344746 93818 344982 94054
rect 344426 93498 344662 93734
rect 344746 93498 344982 93734
rect 344426 57818 344662 58054
rect 344746 57818 344982 58054
rect 344426 57498 344662 57734
rect 344746 57498 344982 57734
rect 344426 21818 344662 22054
rect 344746 21818 344982 22054
rect 344426 21498 344662 21734
rect 344746 21498 344982 21734
rect 344426 -5382 344662 -5146
rect 344746 -5382 344982 -5146
rect 344426 -5702 344662 -5466
rect 344746 -5702 344982 -5466
rect 348146 133538 348382 133774
rect 348466 133538 348702 133774
rect 348146 133218 348382 133454
rect 348466 133218 348702 133454
rect 348146 97538 348382 97774
rect 348466 97538 348702 97774
rect 348146 97218 348382 97454
rect 348466 97218 348702 97454
rect 348146 61538 348382 61774
rect 348466 61538 348702 61774
rect 348146 61218 348382 61454
rect 348466 61218 348702 61454
rect 348146 25538 348382 25774
rect 348466 25538 348702 25774
rect 348146 25218 348382 25454
rect 348466 25218 348702 25454
rect 348146 -6342 348382 -6106
rect 348466 -6342 348702 -6106
rect 348146 -6662 348382 -6426
rect 348466 -6662 348702 -6426
rect 351866 711322 352102 711558
rect 352186 711322 352422 711558
rect 351866 711002 352102 711238
rect 352186 711002 352422 711238
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 351866 677258 352102 677494
rect 352186 677258 352422 677494
rect 351866 676938 352102 677174
rect 352186 676938 352422 677174
rect 351866 641258 352102 641494
rect 352186 641258 352422 641494
rect 351866 640938 352102 641174
rect 352186 640938 352422 641174
rect 351866 605258 352102 605494
rect 352186 605258 352422 605494
rect 351866 604938 352102 605174
rect 352186 604938 352422 605174
rect 351866 569258 352102 569494
rect 352186 569258 352422 569494
rect 351866 568938 352102 569174
rect 352186 568938 352422 569174
rect 351866 533258 352102 533494
rect 352186 533258 352422 533494
rect 351866 532938 352102 533174
rect 352186 532938 352422 533174
rect 351866 497258 352102 497494
rect 352186 497258 352422 497494
rect 351866 496938 352102 497174
rect 352186 496938 352422 497174
rect 351866 461258 352102 461494
rect 352186 461258 352422 461494
rect 351866 460938 352102 461174
rect 352186 460938 352422 461174
rect 351866 425258 352102 425494
rect 352186 425258 352422 425494
rect 351866 424938 352102 425174
rect 352186 424938 352422 425174
rect 351866 389258 352102 389494
rect 352186 389258 352422 389494
rect 351866 388938 352102 389174
rect 352186 388938 352422 389174
rect 351866 353258 352102 353494
rect 352186 353258 352422 353494
rect 351866 352938 352102 353174
rect 352186 352938 352422 353174
rect 351866 317258 352102 317494
rect 352186 317258 352422 317494
rect 351866 316938 352102 317174
rect 352186 316938 352422 317174
rect 351866 281258 352102 281494
rect 352186 281258 352422 281494
rect 351866 280938 352102 281174
rect 352186 280938 352422 281174
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 351866 245258 352102 245494
rect 352186 245258 352422 245494
rect 351866 244938 352102 245174
rect 352186 244938 352422 245174
rect 351866 209258 352102 209494
rect 352186 209258 352422 209494
rect 351866 208938 352102 209174
rect 352186 208938 352422 209174
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 351866 173258 352102 173494
rect 352186 173258 352422 173494
rect 351866 172938 352102 173174
rect 352186 172938 352422 173174
rect 351866 137258 352102 137494
rect 352186 137258 352422 137494
rect 351866 136938 352102 137174
rect 352186 136938 352422 137174
rect 351866 101258 352102 101494
rect 352186 101258 352422 101494
rect 351866 100938 352102 101174
rect 352186 100938 352422 101174
rect 351866 65258 352102 65494
rect 352186 65258 352422 65494
rect 351866 64938 352102 65174
rect 352186 64938 352422 65174
rect 351866 29258 352102 29494
rect 352186 29258 352422 29494
rect 351866 28938 352102 29174
rect 352186 28938 352422 29174
rect 351866 -7302 352102 -7066
rect 352186 -7302 352422 -7066
rect 351866 -7622 352102 -7386
rect 352186 -7622 352422 -7386
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 369266 706522 369502 706758
rect 369586 706522 369822 706758
rect 369266 706202 369502 706438
rect 369586 706202 369822 706438
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -2502 369502 -2266
rect 369586 -2502 369822 -2266
rect 369266 -2822 369502 -2586
rect 369586 -2822 369822 -2586
rect 372986 707482 373222 707718
rect 373306 707482 373542 707718
rect 372986 707162 373222 707398
rect 373306 707162 373542 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 372986 -3462 373222 -3226
rect 373306 -3462 373542 -3226
rect 372986 -3782 373222 -3546
rect 373306 -3782 373542 -3546
rect 376706 708442 376942 708678
rect 377026 708442 377262 708678
rect 376706 708122 376942 708358
rect 377026 708122 377262 708358
rect 376706 666098 376942 666334
rect 377026 666098 377262 666334
rect 376706 665778 376942 666014
rect 377026 665778 377262 666014
rect 376706 630098 376942 630334
rect 377026 630098 377262 630334
rect 376706 629778 376942 630014
rect 377026 629778 377262 630014
rect 376706 594098 376942 594334
rect 377026 594098 377262 594334
rect 376706 593778 376942 594014
rect 377026 593778 377262 594014
rect 376706 558098 376942 558334
rect 377026 558098 377262 558334
rect 376706 557778 376942 558014
rect 377026 557778 377262 558014
rect 376706 522098 376942 522334
rect 377026 522098 377262 522334
rect 376706 521778 376942 522014
rect 377026 521778 377262 522014
rect 376706 486098 376942 486334
rect 377026 486098 377262 486334
rect 376706 485778 376942 486014
rect 377026 485778 377262 486014
rect 376706 450098 376942 450334
rect 377026 450098 377262 450334
rect 376706 449778 376942 450014
rect 377026 449778 377262 450014
rect 376706 414098 376942 414334
rect 377026 414098 377262 414334
rect 376706 413778 376942 414014
rect 377026 413778 377262 414014
rect 376706 378098 376942 378334
rect 377026 378098 377262 378334
rect 376706 377778 376942 378014
rect 377026 377778 377262 378014
rect 376706 342098 376942 342334
rect 377026 342098 377262 342334
rect 376706 341778 376942 342014
rect 377026 341778 377262 342014
rect 376706 306098 376942 306334
rect 377026 306098 377262 306334
rect 376706 305778 376942 306014
rect 377026 305778 377262 306014
rect 376706 270098 376942 270334
rect 377026 270098 377262 270334
rect 376706 269778 376942 270014
rect 377026 269778 377262 270014
rect 376706 234098 376942 234334
rect 377026 234098 377262 234334
rect 376706 233778 376942 234014
rect 377026 233778 377262 234014
rect 376706 198098 376942 198334
rect 377026 198098 377262 198334
rect 376706 197778 376942 198014
rect 377026 197778 377262 198014
rect 376706 162098 376942 162334
rect 377026 162098 377262 162334
rect 376706 161778 376942 162014
rect 377026 161778 377262 162014
rect 376706 126098 376942 126334
rect 377026 126098 377262 126334
rect 376706 125778 376942 126014
rect 377026 125778 377262 126014
rect 376706 90098 376942 90334
rect 377026 90098 377262 90334
rect 376706 89778 376942 90014
rect 377026 89778 377262 90014
rect 376706 54098 376942 54334
rect 377026 54098 377262 54334
rect 376706 53778 376942 54014
rect 377026 53778 377262 54014
rect 376706 18098 376942 18334
rect 377026 18098 377262 18334
rect 376706 17778 376942 18014
rect 377026 17778 377262 18014
rect 376706 -4422 376942 -4186
rect 377026 -4422 377262 -4186
rect 376706 -4742 376942 -4506
rect 377026 -4742 377262 -4506
rect 380426 709402 380662 709638
rect 380746 709402 380982 709638
rect 380426 709082 380662 709318
rect 380746 709082 380982 709318
rect 380426 669818 380662 670054
rect 380746 669818 380982 670054
rect 380426 669498 380662 669734
rect 380746 669498 380982 669734
rect 380426 633818 380662 634054
rect 380746 633818 380982 634054
rect 380426 633498 380662 633734
rect 380746 633498 380982 633734
rect 380426 597818 380662 598054
rect 380746 597818 380982 598054
rect 380426 597498 380662 597734
rect 380746 597498 380982 597734
rect 380426 561818 380662 562054
rect 380746 561818 380982 562054
rect 380426 561498 380662 561734
rect 380746 561498 380982 561734
rect 380426 525818 380662 526054
rect 380746 525818 380982 526054
rect 380426 525498 380662 525734
rect 380746 525498 380982 525734
rect 380426 489818 380662 490054
rect 380746 489818 380982 490054
rect 380426 489498 380662 489734
rect 380746 489498 380982 489734
rect 380426 453818 380662 454054
rect 380746 453818 380982 454054
rect 380426 453498 380662 453734
rect 380746 453498 380982 453734
rect 380426 417818 380662 418054
rect 380746 417818 380982 418054
rect 380426 417498 380662 417734
rect 380746 417498 380982 417734
rect 380426 381818 380662 382054
rect 380746 381818 380982 382054
rect 380426 381498 380662 381734
rect 380746 381498 380982 381734
rect 380426 345818 380662 346054
rect 380746 345818 380982 346054
rect 380426 345498 380662 345734
rect 380746 345498 380982 345734
rect 380426 309818 380662 310054
rect 380746 309818 380982 310054
rect 380426 309498 380662 309734
rect 380746 309498 380982 309734
rect 380426 273818 380662 274054
rect 380746 273818 380982 274054
rect 380426 273498 380662 273734
rect 380746 273498 380982 273734
rect 380426 237818 380662 238054
rect 380746 237818 380982 238054
rect 380426 237498 380662 237734
rect 380746 237498 380982 237734
rect 380426 201818 380662 202054
rect 380746 201818 380982 202054
rect 380426 201498 380662 201734
rect 380746 201498 380982 201734
rect 380426 165818 380662 166054
rect 380746 165818 380982 166054
rect 380426 165498 380662 165734
rect 380746 165498 380982 165734
rect 380426 129818 380662 130054
rect 380746 129818 380982 130054
rect 380426 129498 380662 129734
rect 380746 129498 380982 129734
rect 380426 93818 380662 94054
rect 380746 93818 380982 94054
rect 380426 93498 380662 93734
rect 380746 93498 380982 93734
rect 380426 57818 380662 58054
rect 380746 57818 380982 58054
rect 380426 57498 380662 57734
rect 380746 57498 380982 57734
rect 380426 21818 380662 22054
rect 380746 21818 380982 22054
rect 380426 21498 380662 21734
rect 380746 21498 380982 21734
rect 380426 -5382 380662 -5146
rect 380746 -5382 380982 -5146
rect 380426 -5702 380662 -5466
rect 380746 -5702 380982 -5466
rect 384146 710362 384382 710598
rect 384466 710362 384702 710598
rect 384146 710042 384382 710278
rect 384466 710042 384702 710278
rect 384146 673538 384382 673774
rect 384466 673538 384702 673774
rect 384146 673218 384382 673454
rect 384466 673218 384702 673454
rect 384146 637538 384382 637774
rect 384466 637538 384702 637774
rect 384146 637218 384382 637454
rect 384466 637218 384702 637454
rect 384146 601538 384382 601774
rect 384466 601538 384702 601774
rect 384146 601218 384382 601454
rect 384466 601218 384702 601454
rect 384146 565538 384382 565774
rect 384466 565538 384702 565774
rect 384146 565218 384382 565454
rect 384466 565218 384702 565454
rect 384146 529538 384382 529774
rect 384466 529538 384702 529774
rect 384146 529218 384382 529454
rect 384466 529218 384702 529454
rect 384146 493538 384382 493774
rect 384466 493538 384702 493774
rect 384146 493218 384382 493454
rect 384466 493218 384702 493454
rect 384146 457538 384382 457774
rect 384466 457538 384702 457774
rect 384146 457218 384382 457454
rect 384466 457218 384702 457454
rect 384146 421538 384382 421774
rect 384466 421538 384702 421774
rect 384146 421218 384382 421454
rect 384466 421218 384702 421454
rect 384146 385538 384382 385774
rect 384466 385538 384702 385774
rect 384146 385218 384382 385454
rect 384466 385218 384702 385454
rect 384146 349538 384382 349774
rect 384466 349538 384702 349774
rect 384146 349218 384382 349454
rect 384466 349218 384702 349454
rect 384146 313538 384382 313774
rect 384466 313538 384702 313774
rect 384146 313218 384382 313454
rect 384466 313218 384702 313454
rect 384146 277538 384382 277774
rect 384466 277538 384702 277774
rect 384146 277218 384382 277454
rect 384466 277218 384702 277454
rect 384146 241538 384382 241774
rect 384466 241538 384702 241774
rect 384146 241218 384382 241454
rect 384466 241218 384702 241454
rect 384146 205538 384382 205774
rect 384466 205538 384702 205774
rect 384146 205218 384382 205454
rect 384466 205218 384702 205454
rect 384146 169538 384382 169774
rect 384466 169538 384702 169774
rect 384146 169218 384382 169454
rect 384466 169218 384702 169454
rect 384146 133538 384382 133774
rect 384466 133538 384702 133774
rect 384146 133218 384382 133454
rect 384466 133218 384702 133454
rect 384146 97538 384382 97774
rect 384466 97538 384702 97774
rect 384146 97218 384382 97454
rect 384466 97218 384702 97454
rect 384146 61538 384382 61774
rect 384466 61538 384702 61774
rect 384146 61218 384382 61454
rect 384466 61218 384702 61454
rect 384146 25538 384382 25774
rect 384466 25538 384702 25774
rect 384146 25218 384382 25454
rect 384466 25218 384702 25454
rect 384146 -6342 384382 -6106
rect 384466 -6342 384702 -6106
rect 384146 -6662 384382 -6426
rect 384466 -6662 384702 -6426
rect 387866 711322 388102 711558
rect 388186 711322 388422 711558
rect 387866 711002 388102 711238
rect 388186 711002 388422 711238
rect 387866 677258 388102 677494
rect 388186 677258 388422 677494
rect 387866 676938 388102 677174
rect 388186 676938 388422 677174
rect 387866 641258 388102 641494
rect 388186 641258 388422 641494
rect 387866 640938 388102 641174
rect 388186 640938 388422 641174
rect 387866 605258 388102 605494
rect 388186 605258 388422 605494
rect 387866 604938 388102 605174
rect 388186 604938 388422 605174
rect 387866 569258 388102 569494
rect 388186 569258 388422 569494
rect 387866 568938 388102 569174
rect 388186 568938 388422 569174
rect 387866 533258 388102 533494
rect 388186 533258 388422 533494
rect 387866 532938 388102 533174
rect 388186 532938 388422 533174
rect 387866 497258 388102 497494
rect 388186 497258 388422 497494
rect 387866 496938 388102 497174
rect 388186 496938 388422 497174
rect 387866 461258 388102 461494
rect 388186 461258 388422 461494
rect 387866 460938 388102 461174
rect 388186 460938 388422 461174
rect 387866 425258 388102 425494
rect 388186 425258 388422 425494
rect 387866 424938 388102 425174
rect 388186 424938 388422 425174
rect 387866 389258 388102 389494
rect 388186 389258 388422 389494
rect 387866 388938 388102 389174
rect 388186 388938 388422 389174
rect 387866 353258 388102 353494
rect 388186 353258 388422 353494
rect 387866 352938 388102 353174
rect 388186 352938 388422 353174
rect 387866 317258 388102 317494
rect 388186 317258 388422 317494
rect 387866 316938 388102 317174
rect 388186 316938 388422 317174
rect 387866 281258 388102 281494
rect 388186 281258 388422 281494
rect 387866 280938 388102 281174
rect 388186 280938 388422 281174
rect 387866 245258 388102 245494
rect 388186 245258 388422 245494
rect 387866 244938 388102 245174
rect 388186 244938 388422 245174
rect 387866 209258 388102 209494
rect 388186 209258 388422 209494
rect 387866 208938 388102 209174
rect 388186 208938 388422 209174
rect 387866 173258 388102 173494
rect 388186 173258 388422 173494
rect 387866 172938 388102 173174
rect 388186 172938 388422 173174
rect 387866 137258 388102 137494
rect 388186 137258 388422 137494
rect 387866 136938 388102 137174
rect 388186 136938 388422 137174
rect 387866 101258 388102 101494
rect 388186 101258 388422 101494
rect 387866 100938 388102 101174
rect 388186 100938 388422 101174
rect 387866 65258 388102 65494
rect 388186 65258 388422 65494
rect 387866 64938 388102 65174
rect 388186 64938 388422 65174
rect 387866 29258 388102 29494
rect 388186 29258 388422 29494
rect 387866 28938 388102 29174
rect 388186 28938 388422 29174
rect 387866 -7302 388102 -7066
rect 388186 -7302 388422 -7066
rect 387866 -7622 388102 -7386
rect 388186 -7622 388422 -7386
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 405266 706522 405502 706758
rect 405586 706522 405822 706758
rect 405266 706202 405502 706438
rect 405586 706202 405822 706438
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -2502 405502 -2266
rect 405586 -2502 405822 -2266
rect 405266 -2822 405502 -2586
rect 405586 -2822 405822 -2586
rect 408986 707482 409222 707718
rect 409306 707482 409542 707718
rect 408986 707162 409222 707398
rect 409306 707162 409542 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 408986 -3462 409222 -3226
rect 409306 -3462 409542 -3226
rect 408986 -3782 409222 -3546
rect 409306 -3782 409542 -3546
rect 412706 708442 412942 708678
rect 413026 708442 413262 708678
rect 412706 708122 412942 708358
rect 413026 708122 413262 708358
rect 412706 666098 412942 666334
rect 413026 666098 413262 666334
rect 412706 665778 412942 666014
rect 413026 665778 413262 666014
rect 412706 630098 412942 630334
rect 413026 630098 413262 630334
rect 412706 629778 412942 630014
rect 413026 629778 413262 630014
rect 412706 594098 412942 594334
rect 413026 594098 413262 594334
rect 412706 593778 412942 594014
rect 413026 593778 413262 594014
rect 412706 558098 412942 558334
rect 413026 558098 413262 558334
rect 412706 557778 412942 558014
rect 413026 557778 413262 558014
rect 412706 522098 412942 522334
rect 413026 522098 413262 522334
rect 412706 521778 412942 522014
rect 413026 521778 413262 522014
rect 412706 486098 412942 486334
rect 413026 486098 413262 486334
rect 412706 485778 412942 486014
rect 413026 485778 413262 486014
rect 412706 450098 412942 450334
rect 413026 450098 413262 450334
rect 412706 449778 412942 450014
rect 413026 449778 413262 450014
rect 412706 414098 412942 414334
rect 413026 414098 413262 414334
rect 412706 413778 412942 414014
rect 413026 413778 413262 414014
rect 412706 378098 412942 378334
rect 413026 378098 413262 378334
rect 412706 377778 412942 378014
rect 413026 377778 413262 378014
rect 412706 342098 412942 342334
rect 413026 342098 413262 342334
rect 412706 341778 412942 342014
rect 413026 341778 413262 342014
rect 412706 306098 412942 306334
rect 413026 306098 413262 306334
rect 412706 305778 412942 306014
rect 413026 305778 413262 306014
rect 412706 270098 412942 270334
rect 413026 270098 413262 270334
rect 412706 269778 412942 270014
rect 413026 269778 413262 270014
rect 412706 234098 412942 234334
rect 413026 234098 413262 234334
rect 412706 233778 412942 234014
rect 413026 233778 413262 234014
rect 412706 198098 412942 198334
rect 413026 198098 413262 198334
rect 412706 197778 412942 198014
rect 413026 197778 413262 198014
rect 412706 162098 412942 162334
rect 413026 162098 413262 162334
rect 412706 161778 412942 162014
rect 413026 161778 413262 162014
rect 412706 126098 412942 126334
rect 413026 126098 413262 126334
rect 412706 125778 412942 126014
rect 413026 125778 413262 126014
rect 412706 90098 412942 90334
rect 413026 90098 413262 90334
rect 412706 89778 412942 90014
rect 413026 89778 413262 90014
rect 412706 54098 412942 54334
rect 413026 54098 413262 54334
rect 412706 53778 412942 54014
rect 413026 53778 413262 54014
rect 412706 18098 412942 18334
rect 413026 18098 413262 18334
rect 412706 17778 412942 18014
rect 413026 17778 413262 18014
rect 412706 -4422 412942 -4186
rect 413026 -4422 413262 -4186
rect 412706 -4742 412942 -4506
rect 413026 -4742 413262 -4506
rect 416426 709402 416662 709638
rect 416746 709402 416982 709638
rect 416426 709082 416662 709318
rect 416746 709082 416982 709318
rect 416426 669818 416662 670054
rect 416746 669818 416982 670054
rect 416426 669498 416662 669734
rect 416746 669498 416982 669734
rect 416426 633818 416662 634054
rect 416746 633818 416982 634054
rect 416426 633498 416662 633734
rect 416746 633498 416982 633734
rect 416426 597818 416662 598054
rect 416746 597818 416982 598054
rect 416426 597498 416662 597734
rect 416746 597498 416982 597734
rect 416426 561818 416662 562054
rect 416746 561818 416982 562054
rect 416426 561498 416662 561734
rect 416746 561498 416982 561734
rect 416426 525818 416662 526054
rect 416746 525818 416982 526054
rect 416426 525498 416662 525734
rect 416746 525498 416982 525734
rect 416426 489818 416662 490054
rect 416746 489818 416982 490054
rect 416426 489498 416662 489734
rect 416746 489498 416982 489734
rect 416426 453818 416662 454054
rect 416746 453818 416982 454054
rect 416426 453498 416662 453734
rect 416746 453498 416982 453734
rect 416426 417818 416662 418054
rect 416746 417818 416982 418054
rect 416426 417498 416662 417734
rect 416746 417498 416982 417734
rect 416426 381818 416662 382054
rect 416746 381818 416982 382054
rect 416426 381498 416662 381734
rect 416746 381498 416982 381734
rect 416426 345818 416662 346054
rect 416746 345818 416982 346054
rect 416426 345498 416662 345734
rect 416746 345498 416982 345734
rect 416426 309818 416662 310054
rect 416746 309818 416982 310054
rect 416426 309498 416662 309734
rect 416746 309498 416982 309734
rect 416426 273818 416662 274054
rect 416746 273818 416982 274054
rect 416426 273498 416662 273734
rect 416746 273498 416982 273734
rect 416426 237818 416662 238054
rect 416746 237818 416982 238054
rect 416426 237498 416662 237734
rect 416746 237498 416982 237734
rect 416426 201818 416662 202054
rect 416746 201818 416982 202054
rect 416426 201498 416662 201734
rect 416746 201498 416982 201734
rect 416426 165818 416662 166054
rect 416746 165818 416982 166054
rect 416426 165498 416662 165734
rect 416746 165498 416982 165734
rect 416426 129818 416662 130054
rect 416746 129818 416982 130054
rect 416426 129498 416662 129734
rect 416746 129498 416982 129734
rect 416426 93818 416662 94054
rect 416746 93818 416982 94054
rect 416426 93498 416662 93734
rect 416746 93498 416982 93734
rect 416426 57818 416662 58054
rect 416746 57818 416982 58054
rect 416426 57498 416662 57734
rect 416746 57498 416982 57734
rect 416426 21818 416662 22054
rect 416746 21818 416982 22054
rect 416426 21498 416662 21734
rect 416746 21498 416982 21734
rect 416426 -5382 416662 -5146
rect 416746 -5382 416982 -5146
rect 416426 -5702 416662 -5466
rect 416746 -5702 416982 -5466
rect 420146 710362 420382 710598
rect 420466 710362 420702 710598
rect 420146 710042 420382 710278
rect 420466 710042 420702 710278
rect 420146 673538 420382 673774
rect 420466 673538 420702 673774
rect 420146 673218 420382 673454
rect 420466 673218 420702 673454
rect 420146 637538 420382 637774
rect 420466 637538 420702 637774
rect 420146 637218 420382 637454
rect 420466 637218 420702 637454
rect 420146 601538 420382 601774
rect 420466 601538 420702 601774
rect 420146 601218 420382 601454
rect 420466 601218 420702 601454
rect 420146 565538 420382 565774
rect 420466 565538 420702 565774
rect 420146 565218 420382 565454
rect 420466 565218 420702 565454
rect 420146 529538 420382 529774
rect 420466 529538 420702 529774
rect 420146 529218 420382 529454
rect 420466 529218 420702 529454
rect 420146 493538 420382 493774
rect 420466 493538 420702 493774
rect 420146 493218 420382 493454
rect 420466 493218 420702 493454
rect 420146 457538 420382 457774
rect 420466 457538 420702 457774
rect 420146 457218 420382 457454
rect 420466 457218 420702 457454
rect 420146 421538 420382 421774
rect 420466 421538 420702 421774
rect 420146 421218 420382 421454
rect 420466 421218 420702 421454
rect 420146 385538 420382 385774
rect 420466 385538 420702 385774
rect 420146 385218 420382 385454
rect 420466 385218 420702 385454
rect 420146 349538 420382 349774
rect 420466 349538 420702 349774
rect 420146 349218 420382 349454
rect 420466 349218 420702 349454
rect 420146 313538 420382 313774
rect 420466 313538 420702 313774
rect 420146 313218 420382 313454
rect 420466 313218 420702 313454
rect 420146 277538 420382 277774
rect 420466 277538 420702 277774
rect 420146 277218 420382 277454
rect 420466 277218 420702 277454
rect 420146 241538 420382 241774
rect 420466 241538 420702 241774
rect 420146 241218 420382 241454
rect 420466 241218 420702 241454
rect 420146 205538 420382 205774
rect 420466 205538 420702 205774
rect 420146 205218 420382 205454
rect 420466 205218 420702 205454
rect 420146 169538 420382 169774
rect 420466 169538 420702 169774
rect 420146 169218 420382 169454
rect 420466 169218 420702 169454
rect 420146 133538 420382 133774
rect 420466 133538 420702 133774
rect 420146 133218 420382 133454
rect 420466 133218 420702 133454
rect 420146 97538 420382 97774
rect 420466 97538 420702 97774
rect 420146 97218 420382 97454
rect 420466 97218 420702 97454
rect 420146 61538 420382 61774
rect 420466 61538 420702 61774
rect 420146 61218 420382 61454
rect 420466 61218 420702 61454
rect 420146 25538 420382 25774
rect 420466 25538 420702 25774
rect 420146 25218 420382 25454
rect 420466 25218 420702 25454
rect 420146 -6342 420382 -6106
rect 420466 -6342 420702 -6106
rect 420146 -6662 420382 -6426
rect 420466 -6662 420702 -6426
rect 423866 711322 424102 711558
rect 424186 711322 424422 711558
rect 423866 711002 424102 711238
rect 424186 711002 424422 711238
rect 423866 677258 424102 677494
rect 424186 677258 424422 677494
rect 423866 676938 424102 677174
rect 424186 676938 424422 677174
rect 423866 641258 424102 641494
rect 424186 641258 424422 641494
rect 423866 640938 424102 641174
rect 424186 640938 424422 641174
rect 423866 605258 424102 605494
rect 424186 605258 424422 605494
rect 423866 604938 424102 605174
rect 424186 604938 424422 605174
rect 423866 569258 424102 569494
rect 424186 569258 424422 569494
rect 423866 568938 424102 569174
rect 424186 568938 424422 569174
rect 423866 533258 424102 533494
rect 424186 533258 424422 533494
rect 423866 532938 424102 533174
rect 424186 532938 424422 533174
rect 423866 497258 424102 497494
rect 424186 497258 424422 497494
rect 423866 496938 424102 497174
rect 424186 496938 424422 497174
rect 423866 461258 424102 461494
rect 424186 461258 424422 461494
rect 423866 460938 424102 461174
rect 424186 460938 424422 461174
rect 423866 425258 424102 425494
rect 424186 425258 424422 425494
rect 423866 424938 424102 425174
rect 424186 424938 424422 425174
rect 423866 389258 424102 389494
rect 424186 389258 424422 389494
rect 423866 388938 424102 389174
rect 424186 388938 424422 389174
rect 423866 353258 424102 353494
rect 424186 353258 424422 353494
rect 423866 352938 424102 353174
rect 424186 352938 424422 353174
rect 423866 317258 424102 317494
rect 424186 317258 424422 317494
rect 423866 316938 424102 317174
rect 424186 316938 424422 317174
rect 423866 281258 424102 281494
rect 424186 281258 424422 281494
rect 423866 280938 424102 281174
rect 424186 280938 424422 281174
rect 423866 245258 424102 245494
rect 424186 245258 424422 245494
rect 423866 244938 424102 245174
rect 424186 244938 424422 245174
rect 423866 209258 424102 209494
rect 424186 209258 424422 209494
rect 423866 208938 424102 209174
rect 424186 208938 424422 209174
rect 423866 173258 424102 173494
rect 424186 173258 424422 173494
rect 423866 172938 424102 173174
rect 424186 172938 424422 173174
rect 423866 137258 424102 137494
rect 424186 137258 424422 137494
rect 423866 136938 424102 137174
rect 424186 136938 424422 137174
rect 423866 101258 424102 101494
rect 424186 101258 424422 101494
rect 423866 100938 424102 101174
rect 424186 100938 424422 101174
rect 423866 65258 424102 65494
rect 424186 65258 424422 65494
rect 423866 64938 424102 65174
rect 424186 64938 424422 65174
rect 423866 29258 424102 29494
rect 424186 29258 424422 29494
rect 423866 28938 424102 29174
rect 424186 28938 424422 29174
rect 423866 -7302 424102 -7066
rect 424186 -7302 424422 -7066
rect 423866 -7622 424102 -7386
rect 424186 -7622 424422 -7386
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 441266 706522 441502 706758
rect 441586 706522 441822 706758
rect 441266 706202 441502 706438
rect 441586 706202 441822 706438
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -2502 441502 -2266
rect 441586 -2502 441822 -2266
rect 441266 -2822 441502 -2586
rect 441586 -2822 441822 -2586
rect 444986 707482 445222 707718
rect 445306 707482 445542 707718
rect 444986 707162 445222 707398
rect 445306 707162 445542 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 444986 -3462 445222 -3226
rect 445306 -3462 445542 -3226
rect 444986 -3782 445222 -3546
rect 445306 -3782 445542 -3546
rect 448706 708442 448942 708678
rect 449026 708442 449262 708678
rect 448706 708122 448942 708358
rect 449026 708122 449262 708358
rect 448706 666098 448942 666334
rect 449026 666098 449262 666334
rect 448706 665778 448942 666014
rect 449026 665778 449262 666014
rect 448706 630098 448942 630334
rect 449026 630098 449262 630334
rect 448706 629778 448942 630014
rect 449026 629778 449262 630014
rect 448706 594098 448942 594334
rect 449026 594098 449262 594334
rect 448706 593778 448942 594014
rect 449026 593778 449262 594014
rect 448706 558098 448942 558334
rect 449026 558098 449262 558334
rect 448706 557778 448942 558014
rect 449026 557778 449262 558014
rect 448706 522098 448942 522334
rect 449026 522098 449262 522334
rect 448706 521778 448942 522014
rect 449026 521778 449262 522014
rect 448706 486098 448942 486334
rect 449026 486098 449262 486334
rect 448706 485778 448942 486014
rect 449026 485778 449262 486014
rect 448706 450098 448942 450334
rect 449026 450098 449262 450334
rect 448706 449778 448942 450014
rect 449026 449778 449262 450014
rect 448706 414098 448942 414334
rect 449026 414098 449262 414334
rect 448706 413778 448942 414014
rect 449026 413778 449262 414014
rect 448706 378098 448942 378334
rect 449026 378098 449262 378334
rect 448706 377778 448942 378014
rect 449026 377778 449262 378014
rect 448706 342098 448942 342334
rect 449026 342098 449262 342334
rect 448706 341778 448942 342014
rect 449026 341778 449262 342014
rect 448706 306098 448942 306334
rect 449026 306098 449262 306334
rect 448706 305778 448942 306014
rect 449026 305778 449262 306014
rect 448706 270098 448942 270334
rect 449026 270098 449262 270334
rect 448706 269778 448942 270014
rect 449026 269778 449262 270014
rect 448706 234098 448942 234334
rect 449026 234098 449262 234334
rect 448706 233778 448942 234014
rect 449026 233778 449262 234014
rect 448706 198098 448942 198334
rect 449026 198098 449262 198334
rect 448706 197778 448942 198014
rect 449026 197778 449262 198014
rect 448706 162098 448942 162334
rect 449026 162098 449262 162334
rect 448706 161778 448942 162014
rect 449026 161778 449262 162014
rect 448706 126098 448942 126334
rect 449026 126098 449262 126334
rect 448706 125778 448942 126014
rect 449026 125778 449262 126014
rect 448706 90098 448942 90334
rect 449026 90098 449262 90334
rect 448706 89778 448942 90014
rect 449026 89778 449262 90014
rect 448706 54098 448942 54334
rect 449026 54098 449262 54334
rect 448706 53778 448942 54014
rect 449026 53778 449262 54014
rect 448706 18098 448942 18334
rect 449026 18098 449262 18334
rect 448706 17778 448942 18014
rect 449026 17778 449262 18014
rect 448706 -4422 448942 -4186
rect 449026 -4422 449262 -4186
rect 448706 -4742 448942 -4506
rect 449026 -4742 449262 -4506
rect 452426 709402 452662 709638
rect 452746 709402 452982 709638
rect 452426 709082 452662 709318
rect 452746 709082 452982 709318
rect 452426 669818 452662 670054
rect 452746 669818 452982 670054
rect 452426 669498 452662 669734
rect 452746 669498 452982 669734
rect 452426 633818 452662 634054
rect 452746 633818 452982 634054
rect 452426 633498 452662 633734
rect 452746 633498 452982 633734
rect 452426 597818 452662 598054
rect 452746 597818 452982 598054
rect 452426 597498 452662 597734
rect 452746 597498 452982 597734
rect 452426 561818 452662 562054
rect 452746 561818 452982 562054
rect 452426 561498 452662 561734
rect 452746 561498 452982 561734
rect 452426 525818 452662 526054
rect 452746 525818 452982 526054
rect 452426 525498 452662 525734
rect 452746 525498 452982 525734
rect 452426 489818 452662 490054
rect 452746 489818 452982 490054
rect 452426 489498 452662 489734
rect 452746 489498 452982 489734
rect 452426 453818 452662 454054
rect 452746 453818 452982 454054
rect 452426 453498 452662 453734
rect 452746 453498 452982 453734
rect 452426 417818 452662 418054
rect 452746 417818 452982 418054
rect 452426 417498 452662 417734
rect 452746 417498 452982 417734
rect 452426 381818 452662 382054
rect 452746 381818 452982 382054
rect 452426 381498 452662 381734
rect 452746 381498 452982 381734
rect 452426 345818 452662 346054
rect 452746 345818 452982 346054
rect 452426 345498 452662 345734
rect 452746 345498 452982 345734
rect 452426 309818 452662 310054
rect 452746 309818 452982 310054
rect 452426 309498 452662 309734
rect 452746 309498 452982 309734
rect 452426 273818 452662 274054
rect 452746 273818 452982 274054
rect 452426 273498 452662 273734
rect 452746 273498 452982 273734
rect 452426 237818 452662 238054
rect 452746 237818 452982 238054
rect 452426 237498 452662 237734
rect 452746 237498 452982 237734
rect 452426 201818 452662 202054
rect 452746 201818 452982 202054
rect 452426 201498 452662 201734
rect 452746 201498 452982 201734
rect 452426 165818 452662 166054
rect 452746 165818 452982 166054
rect 452426 165498 452662 165734
rect 452746 165498 452982 165734
rect 452426 129818 452662 130054
rect 452746 129818 452982 130054
rect 452426 129498 452662 129734
rect 452746 129498 452982 129734
rect 452426 93818 452662 94054
rect 452746 93818 452982 94054
rect 452426 93498 452662 93734
rect 452746 93498 452982 93734
rect 452426 57818 452662 58054
rect 452746 57818 452982 58054
rect 452426 57498 452662 57734
rect 452746 57498 452982 57734
rect 452426 21818 452662 22054
rect 452746 21818 452982 22054
rect 452426 21498 452662 21734
rect 452746 21498 452982 21734
rect 452426 -5382 452662 -5146
rect 452746 -5382 452982 -5146
rect 452426 -5702 452662 -5466
rect 452746 -5702 452982 -5466
rect 456146 710362 456382 710598
rect 456466 710362 456702 710598
rect 456146 710042 456382 710278
rect 456466 710042 456702 710278
rect 456146 673538 456382 673774
rect 456466 673538 456702 673774
rect 456146 673218 456382 673454
rect 456466 673218 456702 673454
rect 456146 637538 456382 637774
rect 456466 637538 456702 637774
rect 456146 637218 456382 637454
rect 456466 637218 456702 637454
rect 456146 601538 456382 601774
rect 456466 601538 456702 601774
rect 456146 601218 456382 601454
rect 456466 601218 456702 601454
rect 456146 565538 456382 565774
rect 456466 565538 456702 565774
rect 456146 565218 456382 565454
rect 456466 565218 456702 565454
rect 456146 529538 456382 529774
rect 456466 529538 456702 529774
rect 456146 529218 456382 529454
rect 456466 529218 456702 529454
rect 456146 493538 456382 493774
rect 456466 493538 456702 493774
rect 456146 493218 456382 493454
rect 456466 493218 456702 493454
rect 456146 457538 456382 457774
rect 456466 457538 456702 457774
rect 456146 457218 456382 457454
rect 456466 457218 456702 457454
rect 456146 421538 456382 421774
rect 456466 421538 456702 421774
rect 456146 421218 456382 421454
rect 456466 421218 456702 421454
rect 456146 385538 456382 385774
rect 456466 385538 456702 385774
rect 456146 385218 456382 385454
rect 456466 385218 456702 385454
rect 456146 349538 456382 349774
rect 456466 349538 456702 349774
rect 456146 349218 456382 349454
rect 456466 349218 456702 349454
rect 456146 313538 456382 313774
rect 456466 313538 456702 313774
rect 456146 313218 456382 313454
rect 456466 313218 456702 313454
rect 456146 277538 456382 277774
rect 456466 277538 456702 277774
rect 456146 277218 456382 277454
rect 456466 277218 456702 277454
rect 456146 241538 456382 241774
rect 456466 241538 456702 241774
rect 456146 241218 456382 241454
rect 456466 241218 456702 241454
rect 459866 711322 460102 711558
rect 460186 711322 460422 711558
rect 459866 711002 460102 711238
rect 460186 711002 460422 711238
rect 459866 677258 460102 677494
rect 460186 677258 460422 677494
rect 459866 676938 460102 677174
rect 460186 676938 460422 677174
rect 459866 641258 460102 641494
rect 460186 641258 460422 641494
rect 459866 640938 460102 641174
rect 460186 640938 460422 641174
rect 459866 605258 460102 605494
rect 460186 605258 460422 605494
rect 459866 604938 460102 605174
rect 460186 604938 460422 605174
rect 459866 569258 460102 569494
rect 460186 569258 460422 569494
rect 459866 568938 460102 569174
rect 460186 568938 460422 569174
rect 459866 533258 460102 533494
rect 460186 533258 460422 533494
rect 459866 532938 460102 533174
rect 460186 532938 460422 533174
rect 459866 497258 460102 497494
rect 460186 497258 460422 497494
rect 459866 496938 460102 497174
rect 460186 496938 460422 497174
rect 459866 461258 460102 461494
rect 460186 461258 460422 461494
rect 459866 460938 460102 461174
rect 460186 460938 460422 461174
rect 459866 425258 460102 425494
rect 460186 425258 460422 425494
rect 459866 424938 460102 425174
rect 460186 424938 460422 425174
rect 459866 389258 460102 389494
rect 460186 389258 460422 389494
rect 459866 388938 460102 389174
rect 460186 388938 460422 389174
rect 459866 353258 460102 353494
rect 460186 353258 460422 353494
rect 459866 352938 460102 353174
rect 460186 352938 460422 353174
rect 459866 317258 460102 317494
rect 460186 317258 460422 317494
rect 459866 316938 460102 317174
rect 460186 316938 460422 317174
rect 459866 281258 460102 281494
rect 460186 281258 460422 281494
rect 459866 280938 460102 281174
rect 460186 280938 460422 281174
rect 459866 245258 460102 245494
rect 460186 245258 460422 245494
rect 459866 244938 460102 245174
rect 460186 244938 460422 245174
rect 456146 205538 456382 205774
rect 456466 205538 456702 205774
rect 456146 205218 456382 205454
rect 456466 205218 456702 205454
rect 456146 169538 456382 169774
rect 456466 169538 456702 169774
rect 456146 169218 456382 169454
rect 456466 169218 456702 169454
rect 456146 133538 456382 133774
rect 456466 133538 456702 133774
rect 456146 133218 456382 133454
rect 456466 133218 456702 133454
rect 456146 97538 456382 97774
rect 456466 97538 456702 97774
rect 456146 97218 456382 97454
rect 456466 97218 456702 97454
rect 456146 61538 456382 61774
rect 456466 61538 456702 61774
rect 456146 61218 456382 61454
rect 456466 61218 456702 61454
rect 456146 25538 456382 25774
rect 456466 25538 456702 25774
rect 456146 25218 456382 25454
rect 456466 25218 456702 25454
rect 459866 209258 460102 209494
rect 460186 209258 460422 209494
rect 459866 208938 460102 209174
rect 460186 208938 460422 209174
rect 459866 173258 460102 173494
rect 460186 173258 460422 173494
rect 459866 172938 460102 173174
rect 460186 172938 460422 173174
rect 459866 137258 460102 137494
rect 460186 137258 460422 137494
rect 459866 136938 460102 137174
rect 460186 136938 460422 137174
rect 459866 101258 460102 101494
rect 460186 101258 460422 101494
rect 459866 100938 460102 101174
rect 460186 100938 460422 101174
rect 459866 65258 460102 65494
rect 460186 65258 460422 65494
rect 459866 64938 460102 65174
rect 460186 64938 460422 65174
rect 459866 29258 460102 29494
rect 460186 29258 460422 29494
rect 459866 28938 460102 29174
rect 460186 28938 460422 29174
rect 456146 -6342 456382 -6106
rect 456466 -6342 456702 -6106
rect 456146 -6662 456382 -6426
rect 456466 -6662 456702 -6426
rect 459866 -7302 460102 -7066
rect 460186 -7302 460422 -7066
rect 459866 -7622 460102 -7386
rect 460186 -7622 460422 -7386
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 477266 706522 477502 706758
rect 477586 706522 477822 706758
rect 477266 706202 477502 706438
rect 477586 706202 477822 706438
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -2502 477502 -2266
rect 477586 -2502 477822 -2266
rect 477266 -2822 477502 -2586
rect 477586 -2822 477822 -2586
rect 480986 707482 481222 707718
rect 481306 707482 481542 707718
rect 480986 707162 481222 707398
rect 481306 707162 481542 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 480986 -3462 481222 -3226
rect 481306 -3462 481542 -3226
rect 480986 -3782 481222 -3546
rect 481306 -3782 481542 -3546
rect 484706 708442 484942 708678
rect 485026 708442 485262 708678
rect 484706 708122 484942 708358
rect 485026 708122 485262 708358
rect 484706 666098 484942 666334
rect 485026 666098 485262 666334
rect 484706 665778 484942 666014
rect 485026 665778 485262 666014
rect 484706 630098 484942 630334
rect 485026 630098 485262 630334
rect 484706 629778 484942 630014
rect 485026 629778 485262 630014
rect 484706 594098 484942 594334
rect 485026 594098 485262 594334
rect 484706 593778 484942 594014
rect 485026 593778 485262 594014
rect 484706 558098 484942 558334
rect 485026 558098 485262 558334
rect 484706 557778 484942 558014
rect 485026 557778 485262 558014
rect 484706 522098 484942 522334
rect 485026 522098 485262 522334
rect 484706 521778 484942 522014
rect 485026 521778 485262 522014
rect 484706 486098 484942 486334
rect 485026 486098 485262 486334
rect 484706 485778 484942 486014
rect 485026 485778 485262 486014
rect 484706 450098 484942 450334
rect 485026 450098 485262 450334
rect 484706 449778 484942 450014
rect 485026 449778 485262 450014
rect 484706 414098 484942 414334
rect 485026 414098 485262 414334
rect 484706 413778 484942 414014
rect 485026 413778 485262 414014
rect 484706 378098 484942 378334
rect 485026 378098 485262 378334
rect 484706 377778 484942 378014
rect 485026 377778 485262 378014
rect 484706 342098 484942 342334
rect 485026 342098 485262 342334
rect 484706 341778 484942 342014
rect 485026 341778 485262 342014
rect 484706 306098 484942 306334
rect 485026 306098 485262 306334
rect 484706 305778 484942 306014
rect 485026 305778 485262 306014
rect 484706 270098 484942 270334
rect 485026 270098 485262 270334
rect 484706 269778 484942 270014
rect 485026 269778 485262 270014
rect 484706 234098 484942 234334
rect 485026 234098 485262 234334
rect 484706 233778 484942 234014
rect 485026 233778 485262 234014
rect 484706 198098 484942 198334
rect 485026 198098 485262 198334
rect 484706 197778 484942 198014
rect 485026 197778 485262 198014
rect 484706 162098 484942 162334
rect 485026 162098 485262 162334
rect 484706 161778 484942 162014
rect 485026 161778 485262 162014
rect 484706 126098 484942 126334
rect 485026 126098 485262 126334
rect 484706 125778 484942 126014
rect 485026 125778 485262 126014
rect 484706 90098 484942 90334
rect 485026 90098 485262 90334
rect 484706 89778 484942 90014
rect 485026 89778 485262 90014
rect 484706 54098 484942 54334
rect 485026 54098 485262 54334
rect 484706 53778 484942 54014
rect 485026 53778 485262 54014
rect 484706 18098 484942 18334
rect 485026 18098 485262 18334
rect 484706 17778 484942 18014
rect 485026 17778 485262 18014
rect 484706 -4422 484942 -4186
rect 485026 -4422 485262 -4186
rect 484706 -4742 484942 -4506
rect 485026 -4742 485262 -4506
rect 488426 709402 488662 709638
rect 488746 709402 488982 709638
rect 488426 709082 488662 709318
rect 488746 709082 488982 709318
rect 488426 669818 488662 670054
rect 488746 669818 488982 670054
rect 488426 669498 488662 669734
rect 488746 669498 488982 669734
rect 488426 633818 488662 634054
rect 488746 633818 488982 634054
rect 488426 633498 488662 633734
rect 488746 633498 488982 633734
rect 488426 597818 488662 598054
rect 488746 597818 488982 598054
rect 488426 597498 488662 597734
rect 488746 597498 488982 597734
rect 488426 561818 488662 562054
rect 488746 561818 488982 562054
rect 488426 561498 488662 561734
rect 488746 561498 488982 561734
rect 488426 525818 488662 526054
rect 488746 525818 488982 526054
rect 488426 525498 488662 525734
rect 488746 525498 488982 525734
rect 488426 489818 488662 490054
rect 488746 489818 488982 490054
rect 488426 489498 488662 489734
rect 488746 489498 488982 489734
rect 488426 453818 488662 454054
rect 488746 453818 488982 454054
rect 488426 453498 488662 453734
rect 488746 453498 488982 453734
rect 488426 417818 488662 418054
rect 488746 417818 488982 418054
rect 488426 417498 488662 417734
rect 488746 417498 488982 417734
rect 488426 381818 488662 382054
rect 488746 381818 488982 382054
rect 488426 381498 488662 381734
rect 488746 381498 488982 381734
rect 488426 345818 488662 346054
rect 488746 345818 488982 346054
rect 488426 345498 488662 345734
rect 488746 345498 488982 345734
rect 488426 309818 488662 310054
rect 488746 309818 488982 310054
rect 488426 309498 488662 309734
rect 488746 309498 488982 309734
rect 488426 273818 488662 274054
rect 488746 273818 488982 274054
rect 488426 273498 488662 273734
rect 488746 273498 488982 273734
rect 488426 237818 488662 238054
rect 488746 237818 488982 238054
rect 488426 237498 488662 237734
rect 488746 237498 488982 237734
rect 488426 201818 488662 202054
rect 488746 201818 488982 202054
rect 488426 201498 488662 201734
rect 488746 201498 488982 201734
rect 488426 165818 488662 166054
rect 488746 165818 488982 166054
rect 488426 165498 488662 165734
rect 488746 165498 488982 165734
rect 488426 129818 488662 130054
rect 488746 129818 488982 130054
rect 488426 129498 488662 129734
rect 488746 129498 488982 129734
rect 488426 93818 488662 94054
rect 488746 93818 488982 94054
rect 488426 93498 488662 93734
rect 488746 93498 488982 93734
rect 488426 57818 488662 58054
rect 488746 57818 488982 58054
rect 488426 57498 488662 57734
rect 488746 57498 488982 57734
rect 488426 21818 488662 22054
rect 488746 21818 488982 22054
rect 488426 21498 488662 21734
rect 488746 21498 488982 21734
rect 488426 -5382 488662 -5146
rect 488746 -5382 488982 -5146
rect 488426 -5702 488662 -5466
rect 488746 -5702 488982 -5466
rect 492146 710362 492382 710598
rect 492466 710362 492702 710598
rect 492146 710042 492382 710278
rect 492466 710042 492702 710278
rect 492146 673538 492382 673774
rect 492466 673538 492702 673774
rect 492146 673218 492382 673454
rect 492466 673218 492702 673454
rect 495866 711322 496102 711558
rect 496186 711322 496422 711558
rect 495866 711002 496102 711238
rect 496186 711002 496422 711238
rect 495866 677258 496102 677494
rect 496186 677258 496422 677494
rect 495866 676938 496102 677174
rect 496186 676938 496422 677174
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 513266 706522 513502 706758
rect 513586 706522 513822 706758
rect 513266 706202 513502 706438
rect 513586 706202 513822 706438
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 516986 707482 517222 707718
rect 517306 707482 517542 707718
rect 516986 707162 517222 707398
rect 517306 707162 517542 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 520706 708442 520942 708678
rect 521026 708442 521262 708678
rect 520706 708122 520942 708358
rect 521026 708122 521262 708358
rect 520706 666098 520942 666334
rect 521026 666098 521262 666334
rect 520706 665778 520942 666014
rect 521026 665778 521262 666014
rect 524426 709402 524662 709638
rect 524746 709402 524982 709638
rect 524426 709082 524662 709318
rect 524746 709082 524982 709318
rect 524426 669818 524662 670054
rect 524746 669818 524982 670054
rect 524426 669498 524662 669734
rect 524746 669498 524982 669734
rect 528146 710362 528382 710598
rect 528466 710362 528702 710598
rect 528146 710042 528382 710278
rect 528466 710042 528702 710278
rect 528146 673538 528382 673774
rect 528466 673538 528702 673774
rect 528146 673218 528382 673454
rect 528466 673218 528702 673454
rect 531866 711322 532102 711558
rect 532186 711322 532422 711558
rect 531866 711002 532102 711238
rect 532186 711002 532422 711238
rect 531866 677258 532102 677494
rect 532186 677258 532422 677494
rect 531866 676938 532102 677174
rect 532186 676938 532422 677174
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 494250 651218 494486 651454
rect 494250 650898 494486 651134
rect 524970 651218 525206 651454
rect 524970 650898 525206 651134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 492146 637538 492382 637774
rect 492466 637538 492702 637774
rect 492146 637218 492382 637454
rect 492466 637218 492702 637454
rect 509610 618938 509846 619174
rect 509610 618618 509846 618854
rect 494250 615218 494486 615454
rect 494250 614898 494486 615134
rect 524970 615218 525206 615454
rect 524970 614898 525206 615134
rect 492146 601538 492382 601774
rect 492466 601538 492702 601774
rect 492146 601218 492382 601454
rect 492466 601218 492702 601454
rect 492146 565538 492382 565774
rect 492466 565538 492702 565774
rect 492146 565218 492382 565454
rect 492466 565218 492702 565454
rect 492146 529538 492382 529774
rect 492466 529538 492702 529774
rect 492146 529218 492382 529454
rect 492466 529218 492702 529454
rect 492146 493538 492382 493774
rect 492466 493538 492702 493774
rect 492146 493218 492382 493454
rect 492466 493218 492702 493454
rect 492146 457538 492382 457774
rect 492466 457538 492702 457774
rect 492146 457218 492382 457454
rect 492466 457218 492702 457454
rect 492146 421538 492382 421774
rect 492466 421538 492702 421774
rect 492146 421218 492382 421454
rect 492466 421218 492702 421454
rect 492146 385538 492382 385774
rect 492466 385538 492702 385774
rect 492146 385218 492382 385454
rect 492466 385218 492702 385454
rect 492146 349538 492382 349774
rect 492466 349538 492702 349774
rect 492146 349218 492382 349454
rect 492466 349218 492702 349454
rect 492146 313538 492382 313774
rect 492466 313538 492702 313774
rect 492146 313218 492382 313454
rect 492466 313218 492702 313454
rect 492146 277538 492382 277774
rect 492466 277538 492702 277774
rect 492146 277218 492382 277454
rect 492466 277218 492702 277454
rect 492146 241538 492382 241774
rect 492466 241538 492702 241774
rect 492146 241218 492382 241454
rect 492466 241218 492702 241454
rect 492146 205538 492382 205774
rect 492466 205538 492702 205774
rect 492146 205218 492382 205454
rect 492466 205218 492702 205454
rect 492146 169538 492382 169774
rect 492466 169538 492702 169774
rect 492146 169218 492382 169454
rect 492466 169218 492702 169454
rect 492146 133538 492382 133774
rect 492466 133538 492702 133774
rect 492146 133218 492382 133454
rect 492466 133218 492702 133454
rect 492146 97538 492382 97774
rect 492466 97538 492702 97774
rect 492146 97218 492382 97454
rect 492466 97218 492702 97454
rect 492146 61538 492382 61774
rect 492466 61538 492702 61774
rect 492146 61218 492382 61454
rect 492466 61218 492702 61454
rect 492146 25538 492382 25774
rect 492466 25538 492702 25774
rect 492146 25218 492382 25454
rect 492466 25218 492702 25454
rect 492146 -6342 492382 -6106
rect 492466 -6342 492702 -6106
rect 492146 -6662 492382 -6426
rect 492466 -6662 492702 -6426
rect 495866 569258 496102 569494
rect 496186 569258 496422 569494
rect 495866 568938 496102 569174
rect 496186 568938 496422 569174
rect 495866 533258 496102 533494
rect 496186 533258 496422 533494
rect 495866 532938 496102 533174
rect 496186 532938 496422 533174
rect 495866 497258 496102 497494
rect 496186 497258 496422 497494
rect 495866 496938 496102 497174
rect 496186 496938 496422 497174
rect 495866 461258 496102 461494
rect 496186 461258 496422 461494
rect 495866 460938 496102 461174
rect 496186 460938 496422 461174
rect 495866 425258 496102 425494
rect 496186 425258 496422 425494
rect 495866 424938 496102 425174
rect 496186 424938 496422 425174
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 495866 389258 496102 389494
rect 496186 389258 496422 389494
rect 495866 388938 496102 389174
rect 496186 388938 496422 389174
rect 495866 353258 496102 353494
rect 496186 353258 496422 353494
rect 495866 352938 496102 353174
rect 496186 352938 496422 353174
rect 495866 317258 496102 317494
rect 496186 317258 496422 317494
rect 495866 316938 496102 317174
rect 496186 316938 496422 317174
rect 495866 281258 496102 281494
rect 496186 281258 496422 281494
rect 495866 280938 496102 281174
rect 496186 280938 496422 281174
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 495866 245258 496102 245494
rect 496186 245258 496422 245494
rect 495866 244938 496102 245174
rect 496186 244938 496422 245174
rect 495866 209258 496102 209494
rect 496186 209258 496422 209494
rect 495866 208938 496102 209174
rect 496186 208938 496422 209174
rect 495866 173258 496102 173494
rect 496186 173258 496422 173494
rect 495866 172938 496102 173174
rect 496186 172938 496422 173174
rect 495866 137258 496102 137494
rect 496186 137258 496422 137494
rect 495866 136938 496102 137174
rect 496186 136938 496422 137174
rect 495866 101258 496102 101494
rect 496186 101258 496422 101494
rect 495866 100938 496102 101174
rect 496186 100938 496422 101174
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 495866 65258 496102 65494
rect 496186 65258 496422 65494
rect 495866 64938 496102 65174
rect 496186 64938 496422 65174
rect 495866 29258 496102 29494
rect 496186 29258 496422 29494
rect 495866 28938 496102 29174
rect 496186 28938 496422 29174
rect 495866 -7302 496102 -7066
rect 496186 -7302 496422 -7066
rect 495866 -7622 496102 -7386
rect 496186 -7622 496422 -7386
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -2502 513502 -2266
rect 513586 -2502 513822 -2266
rect 513266 -2822 513502 -2586
rect 513586 -2822 513822 -2586
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 516986 -3462 517222 -3226
rect 517306 -3462 517542 -3226
rect 516986 -3782 517222 -3546
rect 517306 -3782 517542 -3546
rect 520706 594098 520942 594334
rect 521026 594098 521262 594334
rect 520706 593778 520942 594014
rect 521026 593778 521262 594014
rect 520706 558098 520942 558334
rect 521026 558098 521262 558334
rect 520706 557778 520942 558014
rect 521026 557778 521262 558014
rect 520706 522098 520942 522334
rect 521026 522098 521262 522334
rect 520706 521778 520942 522014
rect 521026 521778 521262 522014
rect 520706 486098 520942 486334
rect 521026 486098 521262 486334
rect 520706 485778 520942 486014
rect 521026 485778 521262 486014
rect 520706 450098 520942 450334
rect 521026 450098 521262 450334
rect 520706 449778 520942 450014
rect 521026 449778 521262 450014
rect 520706 414098 520942 414334
rect 521026 414098 521262 414334
rect 520706 413778 520942 414014
rect 521026 413778 521262 414014
rect 520706 378098 520942 378334
rect 521026 378098 521262 378334
rect 520706 377778 520942 378014
rect 521026 377778 521262 378014
rect 520706 342098 520942 342334
rect 521026 342098 521262 342334
rect 520706 341778 520942 342014
rect 521026 341778 521262 342014
rect 520706 306098 520942 306334
rect 521026 306098 521262 306334
rect 520706 305778 520942 306014
rect 521026 305778 521262 306014
rect 520706 270098 520942 270334
rect 521026 270098 521262 270334
rect 520706 269778 520942 270014
rect 521026 269778 521262 270014
rect 520706 234098 520942 234334
rect 521026 234098 521262 234334
rect 520706 233778 520942 234014
rect 521026 233778 521262 234014
rect 520706 198098 520942 198334
rect 521026 198098 521262 198334
rect 520706 197778 520942 198014
rect 521026 197778 521262 198014
rect 520706 162098 520942 162334
rect 521026 162098 521262 162334
rect 520706 161778 520942 162014
rect 521026 161778 521262 162014
rect 520706 126098 520942 126334
rect 521026 126098 521262 126334
rect 520706 125778 520942 126014
rect 521026 125778 521262 126014
rect 520706 90098 520942 90334
rect 521026 90098 521262 90334
rect 520706 89778 520942 90014
rect 521026 89778 521262 90014
rect 520706 54098 520942 54334
rect 521026 54098 521262 54334
rect 520706 53778 520942 54014
rect 521026 53778 521262 54014
rect 520706 18098 520942 18334
rect 521026 18098 521262 18334
rect 520706 17778 520942 18014
rect 521026 17778 521262 18014
rect 520706 -4422 520942 -4186
rect 521026 -4422 521262 -4186
rect 520706 -4742 520942 -4506
rect 521026 -4742 521262 -4506
rect 524426 597818 524662 598054
rect 524746 597818 524982 598054
rect 524426 597498 524662 597734
rect 524746 597498 524982 597734
rect 524426 561818 524662 562054
rect 524746 561818 524982 562054
rect 524426 561498 524662 561734
rect 524746 561498 524982 561734
rect 524426 525818 524662 526054
rect 524746 525818 524982 526054
rect 524426 525498 524662 525734
rect 524746 525498 524982 525734
rect 524426 489818 524662 490054
rect 524746 489818 524982 490054
rect 524426 489498 524662 489734
rect 524746 489498 524982 489734
rect 524426 453818 524662 454054
rect 524746 453818 524982 454054
rect 524426 453498 524662 453734
rect 524746 453498 524982 453734
rect 524426 417818 524662 418054
rect 524746 417818 524982 418054
rect 524426 417498 524662 417734
rect 524746 417498 524982 417734
rect 524426 381818 524662 382054
rect 524746 381818 524982 382054
rect 524426 381498 524662 381734
rect 524746 381498 524982 381734
rect 524426 345818 524662 346054
rect 524746 345818 524982 346054
rect 524426 345498 524662 345734
rect 524746 345498 524982 345734
rect 524426 309818 524662 310054
rect 524746 309818 524982 310054
rect 524426 309498 524662 309734
rect 524746 309498 524982 309734
rect 524426 273818 524662 274054
rect 524746 273818 524982 274054
rect 524426 273498 524662 273734
rect 524746 273498 524982 273734
rect 524426 237818 524662 238054
rect 524746 237818 524982 238054
rect 524426 237498 524662 237734
rect 524746 237498 524982 237734
rect 524426 201818 524662 202054
rect 524746 201818 524982 202054
rect 524426 201498 524662 201734
rect 524746 201498 524982 201734
rect 524426 165818 524662 166054
rect 524746 165818 524982 166054
rect 524426 165498 524662 165734
rect 524746 165498 524982 165734
rect 524426 129818 524662 130054
rect 524746 129818 524982 130054
rect 524426 129498 524662 129734
rect 524746 129498 524982 129734
rect 524426 93818 524662 94054
rect 524746 93818 524982 94054
rect 524426 93498 524662 93734
rect 524746 93498 524982 93734
rect 524426 57818 524662 58054
rect 524746 57818 524982 58054
rect 524426 57498 524662 57734
rect 524746 57498 524982 57734
rect 524426 21818 524662 22054
rect 524746 21818 524982 22054
rect 524426 21498 524662 21734
rect 524746 21498 524982 21734
rect 524426 -5382 524662 -5146
rect 524746 -5382 524982 -5146
rect 524426 -5702 524662 -5466
rect 524746 -5702 524982 -5466
rect 528146 565538 528382 565774
rect 528466 565538 528702 565774
rect 528146 565218 528382 565454
rect 528466 565218 528702 565454
rect 528146 529538 528382 529774
rect 528466 529538 528702 529774
rect 528146 529218 528382 529454
rect 528466 529218 528702 529454
rect 528146 493538 528382 493774
rect 528466 493538 528702 493774
rect 528146 493218 528382 493454
rect 528466 493218 528702 493454
rect 528146 457538 528382 457774
rect 528466 457538 528702 457774
rect 528146 457218 528382 457454
rect 528466 457218 528702 457454
rect 528146 421538 528382 421774
rect 528466 421538 528702 421774
rect 528146 421218 528382 421454
rect 528466 421218 528702 421454
rect 528146 385538 528382 385774
rect 528466 385538 528702 385774
rect 528146 385218 528382 385454
rect 528466 385218 528702 385454
rect 528146 349538 528382 349774
rect 528466 349538 528702 349774
rect 528146 349218 528382 349454
rect 528466 349218 528702 349454
rect 528146 313538 528382 313774
rect 528466 313538 528702 313774
rect 528146 313218 528382 313454
rect 528466 313218 528702 313454
rect 528146 277538 528382 277774
rect 528466 277538 528702 277774
rect 528146 277218 528382 277454
rect 528466 277218 528702 277454
rect 528146 241538 528382 241774
rect 528466 241538 528702 241774
rect 528146 241218 528382 241454
rect 528466 241218 528702 241454
rect 528146 205538 528382 205774
rect 528466 205538 528702 205774
rect 528146 205218 528382 205454
rect 528466 205218 528702 205454
rect 528146 169538 528382 169774
rect 528466 169538 528702 169774
rect 528146 169218 528382 169454
rect 528466 169218 528702 169454
rect 528146 133538 528382 133774
rect 528466 133538 528702 133774
rect 528146 133218 528382 133454
rect 528466 133218 528702 133454
rect 528146 97538 528382 97774
rect 528466 97538 528702 97774
rect 528146 97218 528382 97454
rect 528466 97218 528702 97454
rect 528146 61538 528382 61774
rect 528466 61538 528702 61774
rect 528146 61218 528382 61454
rect 528466 61218 528702 61454
rect 528146 25538 528382 25774
rect 528466 25538 528702 25774
rect 528146 25218 528382 25454
rect 528466 25218 528702 25454
rect 528146 -6342 528382 -6106
rect 528466 -6342 528702 -6106
rect 528146 -6662 528382 -6426
rect 528466 -6662 528702 -6426
rect 531866 569258 532102 569494
rect 532186 569258 532422 569494
rect 531866 568938 532102 569174
rect 532186 568938 532422 569174
rect 531866 533258 532102 533494
rect 532186 533258 532422 533494
rect 531866 532938 532102 533174
rect 532186 532938 532422 533174
rect 531866 497258 532102 497494
rect 532186 497258 532422 497494
rect 531866 496938 532102 497174
rect 532186 496938 532422 497174
rect 531866 461258 532102 461494
rect 532186 461258 532422 461494
rect 531866 460938 532102 461174
rect 532186 460938 532422 461174
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 531866 425258 532102 425494
rect 532186 425258 532422 425494
rect 531866 424938 532102 425174
rect 532186 424938 532422 425174
rect 531866 389258 532102 389494
rect 532186 389258 532422 389494
rect 531866 388938 532102 389174
rect 532186 388938 532422 389174
rect 531866 353258 532102 353494
rect 532186 353258 532422 353494
rect 531866 352938 532102 353174
rect 532186 352938 532422 353174
rect 531866 317258 532102 317494
rect 532186 317258 532422 317494
rect 531866 316938 532102 317174
rect 532186 316938 532422 317174
rect 531866 281258 532102 281494
rect 532186 281258 532422 281494
rect 531866 280938 532102 281174
rect 532186 280938 532422 281174
rect 531866 245258 532102 245494
rect 532186 245258 532422 245494
rect 531866 244938 532102 245174
rect 532186 244938 532422 245174
rect 531866 209258 532102 209494
rect 532186 209258 532422 209494
rect 531866 208938 532102 209174
rect 532186 208938 532422 209174
rect 531866 173258 532102 173494
rect 532186 173258 532422 173494
rect 531866 172938 532102 173174
rect 532186 172938 532422 173174
rect 531866 137258 532102 137494
rect 532186 137258 532422 137494
rect 531866 136938 532102 137174
rect 532186 136938 532422 137174
rect 531866 101258 532102 101494
rect 532186 101258 532422 101494
rect 531866 100938 532102 101174
rect 532186 100938 532422 101174
rect 531866 65258 532102 65494
rect 532186 65258 532422 65494
rect 531866 64938 532102 65174
rect 532186 64938 532422 65174
rect 531866 29258 532102 29494
rect 532186 29258 532422 29494
rect 531866 28938 532102 29174
rect 532186 28938 532422 29174
rect 531866 -7302 532102 -7066
rect 532186 -7302 532422 -7066
rect 531866 -7622 532102 -7386
rect 532186 -7622 532422 -7386
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 549266 706522 549502 706758
rect 549586 706522 549822 706758
rect 549266 706202 549502 706438
rect 549586 706202 549822 706438
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -2502 549502 -2266
rect 549586 -2502 549822 -2266
rect 549266 -2822 549502 -2586
rect 549586 -2822 549822 -2586
rect 552986 707482 553222 707718
rect 553306 707482 553542 707718
rect 552986 707162 553222 707398
rect 553306 707162 553542 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 552986 -3462 553222 -3226
rect 553306 -3462 553542 -3226
rect 552986 -3782 553222 -3546
rect 553306 -3782 553542 -3546
rect 556706 708442 556942 708678
rect 557026 708442 557262 708678
rect 556706 708122 556942 708358
rect 557026 708122 557262 708358
rect 556706 666098 556942 666334
rect 557026 666098 557262 666334
rect 556706 665778 556942 666014
rect 557026 665778 557262 666014
rect 556706 630098 556942 630334
rect 557026 630098 557262 630334
rect 556706 629778 556942 630014
rect 557026 629778 557262 630014
rect 556706 594098 556942 594334
rect 557026 594098 557262 594334
rect 556706 593778 556942 594014
rect 557026 593778 557262 594014
rect 556706 558098 556942 558334
rect 557026 558098 557262 558334
rect 556706 557778 556942 558014
rect 557026 557778 557262 558014
rect 556706 522098 556942 522334
rect 557026 522098 557262 522334
rect 556706 521778 556942 522014
rect 557026 521778 557262 522014
rect 556706 486098 556942 486334
rect 557026 486098 557262 486334
rect 556706 485778 556942 486014
rect 557026 485778 557262 486014
rect 556706 450098 556942 450334
rect 557026 450098 557262 450334
rect 556706 449778 556942 450014
rect 557026 449778 557262 450014
rect 556706 414098 556942 414334
rect 557026 414098 557262 414334
rect 556706 413778 556942 414014
rect 557026 413778 557262 414014
rect 556706 378098 556942 378334
rect 557026 378098 557262 378334
rect 556706 377778 556942 378014
rect 557026 377778 557262 378014
rect 556706 342098 556942 342334
rect 557026 342098 557262 342334
rect 556706 341778 556942 342014
rect 557026 341778 557262 342014
rect 556706 306098 556942 306334
rect 557026 306098 557262 306334
rect 556706 305778 556942 306014
rect 557026 305778 557262 306014
rect 556706 270098 556942 270334
rect 557026 270098 557262 270334
rect 556706 269778 556942 270014
rect 557026 269778 557262 270014
rect 560426 709402 560662 709638
rect 560746 709402 560982 709638
rect 560426 709082 560662 709318
rect 560746 709082 560982 709318
rect 560426 669818 560662 670054
rect 560746 669818 560982 670054
rect 560426 669498 560662 669734
rect 560746 669498 560982 669734
rect 560426 633818 560662 634054
rect 560746 633818 560982 634054
rect 560426 633498 560662 633734
rect 560746 633498 560982 633734
rect 560426 597818 560662 598054
rect 560746 597818 560982 598054
rect 560426 597498 560662 597734
rect 560746 597498 560982 597734
rect 560426 561818 560662 562054
rect 560746 561818 560982 562054
rect 560426 561498 560662 561734
rect 560746 561498 560982 561734
rect 560426 525818 560662 526054
rect 560746 525818 560982 526054
rect 560426 525498 560662 525734
rect 560746 525498 560982 525734
rect 560426 489818 560662 490054
rect 560746 489818 560982 490054
rect 560426 489498 560662 489734
rect 560746 489498 560982 489734
rect 560426 453818 560662 454054
rect 560746 453818 560982 454054
rect 560426 453498 560662 453734
rect 560746 453498 560982 453734
rect 560426 417818 560662 418054
rect 560746 417818 560982 418054
rect 560426 417498 560662 417734
rect 560746 417498 560982 417734
rect 560426 381818 560662 382054
rect 560746 381818 560982 382054
rect 560426 381498 560662 381734
rect 560746 381498 560982 381734
rect 560426 345818 560662 346054
rect 560746 345818 560982 346054
rect 560426 345498 560662 345734
rect 560746 345498 560982 345734
rect 560426 309818 560662 310054
rect 560746 309818 560982 310054
rect 560426 309498 560662 309734
rect 560746 309498 560982 309734
rect 560426 273818 560662 274054
rect 560746 273818 560982 274054
rect 560426 273498 560662 273734
rect 560746 273498 560982 273734
rect 556706 234098 556942 234334
rect 557026 234098 557262 234334
rect 556706 233778 556942 234014
rect 557026 233778 557262 234014
rect 556706 198098 556942 198334
rect 557026 198098 557262 198334
rect 556706 197778 556942 198014
rect 557026 197778 557262 198014
rect 556706 162098 556942 162334
rect 557026 162098 557262 162334
rect 556706 161778 556942 162014
rect 557026 161778 557262 162014
rect 556706 126098 556942 126334
rect 557026 126098 557262 126334
rect 556706 125778 556942 126014
rect 557026 125778 557262 126014
rect 556706 90098 556942 90334
rect 557026 90098 557262 90334
rect 556706 89778 556942 90014
rect 557026 89778 557262 90014
rect 560426 237818 560662 238054
rect 560746 237818 560982 238054
rect 560426 237498 560662 237734
rect 560746 237498 560982 237734
rect 560426 201818 560662 202054
rect 560746 201818 560982 202054
rect 560426 201498 560662 201734
rect 560746 201498 560982 201734
rect 560426 165818 560662 166054
rect 560746 165818 560982 166054
rect 560426 165498 560662 165734
rect 560746 165498 560982 165734
rect 560426 129818 560662 130054
rect 560746 129818 560982 130054
rect 560426 129498 560662 129734
rect 560746 129498 560982 129734
rect 560426 93818 560662 94054
rect 560746 93818 560982 94054
rect 560426 93498 560662 93734
rect 560746 93498 560982 93734
rect 556706 54098 556942 54334
rect 557026 54098 557262 54334
rect 556706 53778 556942 54014
rect 557026 53778 557262 54014
rect 556706 18098 556942 18334
rect 557026 18098 557262 18334
rect 556706 17778 556942 18014
rect 557026 17778 557262 18014
rect 556706 -4422 556942 -4186
rect 557026 -4422 557262 -4186
rect 556706 -4742 556942 -4506
rect 557026 -4742 557262 -4506
rect 560426 57818 560662 58054
rect 560746 57818 560982 58054
rect 560426 57498 560662 57734
rect 560746 57498 560982 57734
rect 560426 21818 560662 22054
rect 560746 21818 560982 22054
rect 560426 21498 560662 21734
rect 560746 21498 560982 21734
rect 560426 -5382 560662 -5146
rect 560746 -5382 560982 -5146
rect 560426 -5702 560662 -5466
rect 560746 -5702 560982 -5466
rect 564146 710362 564382 710598
rect 564466 710362 564702 710598
rect 564146 710042 564382 710278
rect 564466 710042 564702 710278
rect 564146 673538 564382 673774
rect 564466 673538 564702 673774
rect 564146 673218 564382 673454
rect 564466 673218 564702 673454
rect 564146 637538 564382 637774
rect 564466 637538 564702 637774
rect 564146 637218 564382 637454
rect 564466 637218 564702 637454
rect 564146 601538 564382 601774
rect 564466 601538 564702 601774
rect 564146 601218 564382 601454
rect 564466 601218 564702 601454
rect 564146 565538 564382 565774
rect 564466 565538 564702 565774
rect 564146 565218 564382 565454
rect 564466 565218 564702 565454
rect 564146 529538 564382 529774
rect 564466 529538 564702 529774
rect 564146 529218 564382 529454
rect 564466 529218 564702 529454
rect 564146 493538 564382 493774
rect 564466 493538 564702 493774
rect 564146 493218 564382 493454
rect 564466 493218 564702 493454
rect 564146 457538 564382 457774
rect 564466 457538 564702 457774
rect 564146 457218 564382 457454
rect 564466 457218 564702 457454
rect 564146 421538 564382 421774
rect 564466 421538 564702 421774
rect 564146 421218 564382 421454
rect 564466 421218 564702 421454
rect 564146 385538 564382 385774
rect 564466 385538 564702 385774
rect 564146 385218 564382 385454
rect 564466 385218 564702 385454
rect 564146 349538 564382 349774
rect 564466 349538 564702 349774
rect 564146 349218 564382 349454
rect 564466 349218 564702 349454
rect 564146 313538 564382 313774
rect 564466 313538 564702 313774
rect 564146 313218 564382 313454
rect 564466 313218 564702 313454
rect 564146 277538 564382 277774
rect 564466 277538 564702 277774
rect 564146 277218 564382 277454
rect 564466 277218 564702 277454
rect 564146 241538 564382 241774
rect 564466 241538 564702 241774
rect 564146 241218 564382 241454
rect 564466 241218 564702 241454
rect 564146 205538 564382 205774
rect 564466 205538 564702 205774
rect 564146 205218 564382 205454
rect 564466 205218 564702 205454
rect 564146 169538 564382 169774
rect 564466 169538 564702 169774
rect 564146 169218 564382 169454
rect 564466 169218 564702 169454
rect 564146 133538 564382 133774
rect 564466 133538 564702 133774
rect 564146 133218 564382 133454
rect 564466 133218 564702 133454
rect 564146 97538 564382 97774
rect 564466 97538 564702 97774
rect 564146 97218 564382 97454
rect 564466 97218 564702 97454
rect 564146 61538 564382 61774
rect 564466 61538 564702 61774
rect 564146 61218 564382 61454
rect 564466 61218 564702 61454
rect 564146 25538 564382 25774
rect 564466 25538 564702 25774
rect 564146 25218 564382 25454
rect 564466 25218 564702 25454
rect 564146 -6342 564382 -6106
rect 564466 -6342 564702 -6106
rect 564146 -6662 564382 -6426
rect 564466 -6662 564702 -6426
rect 567866 711322 568102 711558
rect 568186 711322 568422 711558
rect 567866 711002 568102 711238
rect 568186 711002 568422 711238
rect 567866 677258 568102 677494
rect 568186 677258 568422 677494
rect 567866 676938 568102 677174
rect 568186 676938 568422 677174
rect 567866 641258 568102 641494
rect 568186 641258 568422 641494
rect 567866 640938 568102 641174
rect 568186 640938 568422 641174
rect 567866 605258 568102 605494
rect 568186 605258 568422 605494
rect 567866 604938 568102 605174
rect 568186 604938 568422 605174
rect 567866 569258 568102 569494
rect 568186 569258 568422 569494
rect 567866 568938 568102 569174
rect 568186 568938 568422 569174
rect 567866 533258 568102 533494
rect 568186 533258 568422 533494
rect 567866 532938 568102 533174
rect 568186 532938 568422 533174
rect 567866 497258 568102 497494
rect 568186 497258 568422 497494
rect 567866 496938 568102 497174
rect 568186 496938 568422 497174
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 567866 461258 568102 461494
rect 568186 461258 568422 461494
rect 567866 460938 568102 461174
rect 568186 460938 568422 461174
rect 567866 425258 568102 425494
rect 568186 425258 568422 425494
rect 567866 424938 568102 425174
rect 568186 424938 568422 425174
rect 567866 389258 568102 389494
rect 568186 389258 568422 389494
rect 567866 388938 568102 389174
rect 568186 388938 568422 389174
rect 567866 353258 568102 353494
rect 568186 353258 568422 353494
rect 567866 352938 568102 353174
rect 568186 352938 568422 353174
rect 567866 317258 568102 317494
rect 568186 317258 568422 317494
rect 567866 316938 568102 317174
rect 568186 316938 568422 317174
rect 567866 281258 568102 281494
rect 568186 281258 568422 281494
rect 567866 280938 568102 281174
rect 568186 280938 568422 281174
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 567866 245258 568102 245494
rect 568186 245258 568422 245494
rect 567866 244938 568102 245174
rect 568186 244938 568422 245174
rect 567866 209258 568102 209494
rect 568186 209258 568422 209494
rect 567866 208938 568102 209174
rect 568186 208938 568422 209174
rect 567866 173258 568102 173494
rect 568186 173258 568422 173494
rect 567866 172938 568102 173174
rect 568186 172938 568422 173174
rect 567866 137258 568102 137494
rect 568186 137258 568422 137494
rect 567866 136938 568102 137174
rect 568186 136938 568422 137174
rect 567866 101258 568102 101494
rect 568186 101258 568422 101494
rect 567866 100938 568102 101174
rect 568186 100938 568422 101174
rect 567866 65258 568102 65494
rect 568186 65258 568422 65494
rect 567866 64938 568102 65174
rect 568186 64938 568422 65174
rect 567866 29258 568102 29494
rect 568186 29258 568422 29494
rect 567866 28938 568102 29174
rect 568186 28938 568422 29174
rect 567866 -7302 568102 -7066
rect 568186 -7302 568422 -7066
rect 567866 -7622 568102 -7386
rect 568186 -7622 568422 -7386
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 694658 587498 694894
rect 587582 694658 587818 694894
rect 587262 694338 587498 694574
rect 587582 694338 587818 694574
rect 587262 658658 587498 658894
rect 587582 658658 587818 658894
rect 587262 658338 587498 658574
rect 587582 658338 587818 658574
rect 587262 622658 587498 622894
rect 587582 622658 587818 622894
rect 587262 622338 587498 622574
rect 587582 622338 587818 622574
rect 587262 586658 587498 586894
rect 587582 586658 587818 586894
rect 587262 586338 587498 586574
rect 587582 586338 587818 586574
rect 587262 550658 587498 550894
rect 587582 550658 587818 550894
rect 587262 550338 587498 550574
rect 587582 550338 587818 550574
rect 587262 514658 587498 514894
rect 587582 514658 587818 514894
rect 587262 514338 587498 514574
rect 587582 514338 587818 514574
rect 587262 478658 587498 478894
rect 587582 478658 587818 478894
rect 587262 478338 587498 478574
rect 587582 478338 587818 478574
rect 587262 442658 587498 442894
rect 587582 442658 587818 442894
rect 587262 442338 587498 442574
rect 587582 442338 587818 442574
rect 587262 406658 587498 406894
rect 587582 406658 587818 406894
rect 587262 406338 587498 406574
rect 587582 406338 587818 406574
rect 587262 370658 587498 370894
rect 587582 370658 587818 370894
rect 587262 370338 587498 370574
rect 587582 370338 587818 370574
rect 587262 334658 587498 334894
rect 587582 334658 587818 334894
rect 587262 334338 587498 334574
rect 587582 334338 587818 334574
rect 587262 298658 587498 298894
rect 587582 298658 587818 298894
rect 587262 298338 587498 298574
rect 587582 298338 587818 298574
rect 587262 262658 587498 262894
rect 587582 262658 587818 262894
rect 587262 262338 587498 262574
rect 587582 262338 587818 262574
rect 587262 226658 587498 226894
rect 587582 226658 587818 226894
rect 587262 226338 587498 226574
rect 587582 226338 587818 226574
rect 587262 190658 587498 190894
rect 587582 190658 587818 190894
rect 587262 190338 587498 190574
rect 587582 190338 587818 190574
rect 587262 154658 587498 154894
rect 587582 154658 587818 154894
rect 587262 154338 587498 154574
rect 587582 154338 587818 154574
rect 587262 118658 587498 118894
rect 587582 118658 587818 118894
rect 587262 118338 587498 118574
rect 587582 118338 587818 118574
rect 587262 82658 587498 82894
rect 587582 82658 587818 82894
rect 587262 82338 587498 82574
rect 587582 82338 587818 82574
rect 587262 46658 587498 46894
rect 587582 46658 587818 46894
rect 587262 46338 587498 46574
rect 587582 46338 587818 46574
rect 587262 10658 587498 10894
rect 587582 10658 587818 10894
rect 587262 10338 587498 10574
rect 587582 10338 587818 10574
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 698378 588458 698614
rect 588542 698378 588778 698614
rect 588222 698058 588458 698294
rect 588542 698058 588778 698294
rect 588222 662378 588458 662614
rect 588542 662378 588778 662614
rect 588222 662058 588458 662294
rect 588542 662058 588778 662294
rect 588222 626378 588458 626614
rect 588542 626378 588778 626614
rect 588222 626058 588458 626294
rect 588542 626058 588778 626294
rect 588222 590378 588458 590614
rect 588542 590378 588778 590614
rect 588222 590058 588458 590294
rect 588542 590058 588778 590294
rect 588222 554378 588458 554614
rect 588542 554378 588778 554614
rect 588222 554058 588458 554294
rect 588542 554058 588778 554294
rect 588222 518378 588458 518614
rect 588542 518378 588778 518614
rect 588222 518058 588458 518294
rect 588542 518058 588778 518294
rect 588222 482378 588458 482614
rect 588542 482378 588778 482614
rect 588222 482058 588458 482294
rect 588542 482058 588778 482294
rect 588222 446378 588458 446614
rect 588542 446378 588778 446614
rect 588222 446058 588458 446294
rect 588542 446058 588778 446294
rect 588222 410378 588458 410614
rect 588542 410378 588778 410614
rect 588222 410058 588458 410294
rect 588542 410058 588778 410294
rect 588222 374378 588458 374614
rect 588542 374378 588778 374614
rect 588222 374058 588458 374294
rect 588542 374058 588778 374294
rect 588222 338378 588458 338614
rect 588542 338378 588778 338614
rect 588222 338058 588458 338294
rect 588542 338058 588778 338294
rect 588222 302378 588458 302614
rect 588542 302378 588778 302614
rect 588222 302058 588458 302294
rect 588542 302058 588778 302294
rect 588222 266378 588458 266614
rect 588542 266378 588778 266614
rect 588222 266058 588458 266294
rect 588542 266058 588778 266294
rect 588222 230378 588458 230614
rect 588542 230378 588778 230614
rect 588222 230058 588458 230294
rect 588542 230058 588778 230294
rect 588222 194378 588458 194614
rect 588542 194378 588778 194614
rect 588222 194058 588458 194294
rect 588542 194058 588778 194294
rect 588222 158378 588458 158614
rect 588542 158378 588778 158614
rect 588222 158058 588458 158294
rect 588542 158058 588778 158294
rect 588222 122378 588458 122614
rect 588542 122378 588778 122614
rect 588222 122058 588458 122294
rect 588542 122058 588778 122294
rect 588222 86378 588458 86614
rect 588542 86378 588778 86614
rect 588222 86058 588458 86294
rect 588542 86058 588778 86294
rect 588222 50378 588458 50614
rect 588542 50378 588778 50614
rect 588222 50058 588458 50294
rect 588542 50058 588778 50294
rect 588222 14378 588458 14614
rect 588542 14378 588778 14614
rect 588222 14058 588458 14294
rect 588542 14058 588778 14294
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 666098 589418 666334
rect 589502 666098 589738 666334
rect 589182 665778 589418 666014
rect 589502 665778 589738 666014
rect 589182 630098 589418 630334
rect 589502 630098 589738 630334
rect 589182 629778 589418 630014
rect 589502 629778 589738 630014
rect 589182 594098 589418 594334
rect 589502 594098 589738 594334
rect 589182 593778 589418 594014
rect 589502 593778 589738 594014
rect 589182 558098 589418 558334
rect 589502 558098 589738 558334
rect 589182 557778 589418 558014
rect 589502 557778 589738 558014
rect 589182 522098 589418 522334
rect 589502 522098 589738 522334
rect 589182 521778 589418 522014
rect 589502 521778 589738 522014
rect 589182 486098 589418 486334
rect 589502 486098 589738 486334
rect 589182 485778 589418 486014
rect 589502 485778 589738 486014
rect 589182 450098 589418 450334
rect 589502 450098 589738 450334
rect 589182 449778 589418 450014
rect 589502 449778 589738 450014
rect 589182 414098 589418 414334
rect 589502 414098 589738 414334
rect 589182 413778 589418 414014
rect 589502 413778 589738 414014
rect 589182 378098 589418 378334
rect 589502 378098 589738 378334
rect 589182 377778 589418 378014
rect 589502 377778 589738 378014
rect 589182 342098 589418 342334
rect 589502 342098 589738 342334
rect 589182 341778 589418 342014
rect 589502 341778 589738 342014
rect 589182 306098 589418 306334
rect 589502 306098 589738 306334
rect 589182 305778 589418 306014
rect 589502 305778 589738 306014
rect 589182 270098 589418 270334
rect 589502 270098 589738 270334
rect 589182 269778 589418 270014
rect 589502 269778 589738 270014
rect 589182 234098 589418 234334
rect 589502 234098 589738 234334
rect 589182 233778 589418 234014
rect 589502 233778 589738 234014
rect 589182 198098 589418 198334
rect 589502 198098 589738 198334
rect 589182 197778 589418 198014
rect 589502 197778 589738 198014
rect 589182 162098 589418 162334
rect 589502 162098 589738 162334
rect 589182 161778 589418 162014
rect 589502 161778 589738 162014
rect 589182 126098 589418 126334
rect 589502 126098 589738 126334
rect 589182 125778 589418 126014
rect 589502 125778 589738 126014
rect 589182 90098 589418 90334
rect 589502 90098 589738 90334
rect 589182 89778 589418 90014
rect 589502 89778 589738 90014
rect 589182 54098 589418 54334
rect 589502 54098 589738 54334
rect 589182 53778 589418 54014
rect 589502 53778 589738 54014
rect 589182 18098 589418 18334
rect 589502 18098 589738 18334
rect 589182 17778 589418 18014
rect 589502 17778 589738 18014
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 669818 590378 670054
rect 590462 669818 590698 670054
rect 590142 669498 590378 669734
rect 590462 669498 590698 669734
rect 590142 633818 590378 634054
rect 590462 633818 590698 634054
rect 590142 633498 590378 633734
rect 590462 633498 590698 633734
rect 590142 597818 590378 598054
rect 590462 597818 590698 598054
rect 590142 597498 590378 597734
rect 590462 597498 590698 597734
rect 590142 561818 590378 562054
rect 590462 561818 590698 562054
rect 590142 561498 590378 561734
rect 590462 561498 590698 561734
rect 590142 525818 590378 526054
rect 590462 525818 590698 526054
rect 590142 525498 590378 525734
rect 590462 525498 590698 525734
rect 590142 489818 590378 490054
rect 590462 489818 590698 490054
rect 590142 489498 590378 489734
rect 590462 489498 590698 489734
rect 590142 453818 590378 454054
rect 590462 453818 590698 454054
rect 590142 453498 590378 453734
rect 590462 453498 590698 453734
rect 590142 417818 590378 418054
rect 590462 417818 590698 418054
rect 590142 417498 590378 417734
rect 590462 417498 590698 417734
rect 590142 381818 590378 382054
rect 590462 381818 590698 382054
rect 590142 381498 590378 381734
rect 590462 381498 590698 381734
rect 590142 345818 590378 346054
rect 590462 345818 590698 346054
rect 590142 345498 590378 345734
rect 590462 345498 590698 345734
rect 590142 309818 590378 310054
rect 590462 309818 590698 310054
rect 590142 309498 590378 309734
rect 590462 309498 590698 309734
rect 590142 273818 590378 274054
rect 590462 273818 590698 274054
rect 590142 273498 590378 273734
rect 590462 273498 590698 273734
rect 590142 237818 590378 238054
rect 590462 237818 590698 238054
rect 590142 237498 590378 237734
rect 590462 237498 590698 237734
rect 590142 201818 590378 202054
rect 590462 201818 590698 202054
rect 590142 201498 590378 201734
rect 590462 201498 590698 201734
rect 590142 165818 590378 166054
rect 590462 165818 590698 166054
rect 590142 165498 590378 165734
rect 590462 165498 590698 165734
rect 590142 129818 590378 130054
rect 590462 129818 590698 130054
rect 590142 129498 590378 129734
rect 590462 129498 590698 129734
rect 590142 93818 590378 94054
rect 590462 93818 590698 94054
rect 590142 93498 590378 93734
rect 590462 93498 590698 93734
rect 590142 57818 590378 58054
rect 590462 57818 590698 58054
rect 590142 57498 590378 57734
rect 590462 57498 590698 57734
rect 590142 21818 590378 22054
rect 590462 21818 590698 22054
rect 590142 21498 590378 21734
rect 590462 21498 590698 21734
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673538 591338 673774
rect 591422 673538 591658 673774
rect 591102 673218 591338 673454
rect 591422 673218 591658 673454
rect 591102 637538 591338 637774
rect 591422 637538 591658 637774
rect 591102 637218 591338 637454
rect 591422 637218 591658 637454
rect 591102 601538 591338 601774
rect 591422 601538 591658 601774
rect 591102 601218 591338 601454
rect 591422 601218 591658 601454
rect 591102 565538 591338 565774
rect 591422 565538 591658 565774
rect 591102 565218 591338 565454
rect 591422 565218 591658 565454
rect 591102 529538 591338 529774
rect 591422 529538 591658 529774
rect 591102 529218 591338 529454
rect 591422 529218 591658 529454
rect 591102 493538 591338 493774
rect 591422 493538 591658 493774
rect 591102 493218 591338 493454
rect 591422 493218 591658 493454
rect 591102 457538 591338 457774
rect 591422 457538 591658 457774
rect 591102 457218 591338 457454
rect 591422 457218 591658 457454
rect 591102 421538 591338 421774
rect 591422 421538 591658 421774
rect 591102 421218 591338 421454
rect 591422 421218 591658 421454
rect 591102 385538 591338 385774
rect 591422 385538 591658 385774
rect 591102 385218 591338 385454
rect 591422 385218 591658 385454
rect 591102 349538 591338 349774
rect 591422 349538 591658 349774
rect 591102 349218 591338 349454
rect 591422 349218 591658 349454
rect 591102 313538 591338 313774
rect 591422 313538 591658 313774
rect 591102 313218 591338 313454
rect 591422 313218 591658 313454
rect 591102 277538 591338 277774
rect 591422 277538 591658 277774
rect 591102 277218 591338 277454
rect 591422 277218 591658 277454
rect 591102 241538 591338 241774
rect 591422 241538 591658 241774
rect 591102 241218 591338 241454
rect 591422 241218 591658 241454
rect 591102 205538 591338 205774
rect 591422 205538 591658 205774
rect 591102 205218 591338 205454
rect 591422 205218 591658 205454
rect 591102 169538 591338 169774
rect 591422 169538 591658 169774
rect 591102 169218 591338 169454
rect 591422 169218 591658 169454
rect 591102 133538 591338 133774
rect 591422 133538 591658 133774
rect 591102 133218 591338 133454
rect 591422 133218 591658 133454
rect 591102 97538 591338 97774
rect 591422 97538 591658 97774
rect 591102 97218 591338 97454
rect 591422 97218 591658 97454
rect 591102 61538 591338 61774
rect 591422 61538 591658 61774
rect 591102 61218 591338 61454
rect 591422 61218 591658 61454
rect 591102 25538 591338 25774
rect 591422 25538 591658 25774
rect 591102 25218 591338 25454
rect 591422 25218 591658 25454
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 677258 592298 677494
rect 592382 677258 592618 677494
rect 592062 676938 592298 677174
rect 592382 676938 592618 677174
rect 592062 641258 592298 641494
rect 592382 641258 592618 641494
rect 592062 640938 592298 641174
rect 592382 640938 592618 641174
rect 592062 605258 592298 605494
rect 592382 605258 592618 605494
rect 592062 604938 592298 605174
rect 592382 604938 592618 605174
rect 592062 569258 592298 569494
rect 592382 569258 592618 569494
rect 592062 568938 592298 569174
rect 592382 568938 592618 569174
rect 592062 533258 592298 533494
rect 592382 533258 592618 533494
rect 592062 532938 592298 533174
rect 592382 532938 592618 533174
rect 592062 497258 592298 497494
rect 592382 497258 592618 497494
rect 592062 496938 592298 497174
rect 592382 496938 592618 497174
rect 592062 461258 592298 461494
rect 592382 461258 592618 461494
rect 592062 460938 592298 461174
rect 592382 460938 592618 461174
rect 592062 425258 592298 425494
rect 592382 425258 592618 425494
rect 592062 424938 592298 425174
rect 592382 424938 592618 425174
rect 592062 389258 592298 389494
rect 592382 389258 592618 389494
rect 592062 388938 592298 389174
rect 592382 388938 592618 389174
rect 592062 353258 592298 353494
rect 592382 353258 592618 353494
rect 592062 352938 592298 353174
rect 592382 352938 592618 353174
rect 592062 317258 592298 317494
rect 592382 317258 592618 317494
rect 592062 316938 592298 317174
rect 592382 316938 592618 317174
rect 592062 281258 592298 281494
rect 592382 281258 592618 281494
rect 592062 280938 592298 281174
rect 592382 280938 592618 281174
rect 592062 245258 592298 245494
rect 592382 245258 592618 245494
rect 592062 244938 592298 245174
rect 592382 244938 592618 245174
rect 592062 209258 592298 209494
rect 592382 209258 592618 209494
rect 592062 208938 592298 209174
rect 592382 208938 592618 209174
rect 592062 173258 592298 173494
rect 592382 173258 592618 173494
rect 592062 172938 592298 173174
rect 592382 172938 592618 173174
rect 592062 137258 592298 137494
rect 592382 137258 592618 137494
rect 592062 136938 592298 137174
rect 592382 136938 592618 137174
rect 592062 101258 592298 101494
rect 592382 101258 592618 101494
rect 592062 100938 592298 101174
rect 592382 100938 592618 101174
rect 592062 65258 592298 65494
rect 592382 65258 592618 65494
rect 592062 64938 592298 65174
rect 592382 64938 592618 65174
rect 592062 29258 592298 29494
rect 592382 29258 592618 29494
rect 592062 28938 592298 29174
rect 592382 28938 592618 29174
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 315866 711558
rect 316102 711322 316186 711558
rect 316422 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 315866 711238
rect 316102 711002 316186 711238
rect 316422 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 60146 710598
rect 60382 710362 60466 710598
rect 60702 710362 96146 710598
rect 96382 710362 96466 710598
rect 96702 710362 132146 710598
rect 132382 710362 132466 710598
rect 132702 710362 168146 710598
rect 168382 710362 168466 710598
rect 168702 710362 204146 710598
rect 204382 710362 204466 710598
rect 204702 710362 240146 710598
rect 240382 710362 240466 710598
rect 240702 710362 276146 710598
rect 276382 710362 276466 710598
rect 276702 710362 312146 710598
rect 312382 710362 312466 710598
rect 312702 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 60146 710278
rect 60382 710042 60466 710278
rect 60702 710042 96146 710278
rect 96382 710042 96466 710278
rect 96702 710042 132146 710278
rect 132382 710042 132466 710278
rect 132702 710042 168146 710278
rect 168382 710042 168466 710278
rect 168702 710042 204146 710278
rect 204382 710042 204466 710278
rect 204702 710042 240146 710278
rect 240382 710042 240466 710278
rect 240702 710042 276146 710278
rect 276382 710042 276466 710278
rect 276702 710042 312146 710278
rect 312382 710042 312466 710278
rect 312702 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 56426 709638
rect 56662 709402 56746 709638
rect 56982 709402 92426 709638
rect 92662 709402 92746 709638
rect 92982 709402 128426 709638
rect 128662 709402 128746 709638
rect 128982 709402 164426 709638
rect 164662 709402 164746 709638
rect 164982 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 236426 709638
rect 236662 709402 236746 709638
rect 236982 709402 272426 709638
rect 272662 709402 272746 709638
rect 272982 709402 308426 709638
rect 308662 709402 308746 709638
rect 308982 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 56426 709318
rect 56662 709082 56746 709318
rect 56982 709082 92426 709318
rect 92662 709082 92746 709318
rect 92982 709082 128426 709318
rect 128662 709082 128746 709318
rect 128982 709082 164426 709318
rect 164662 709082 164746 709318
rect 164982 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 236426 709318
rect 236662 709082 236746 709318
rect 236982 709082 272426 709318
rect 272662 709082 272746 709318
rect 272982 709082 308426 709318
rect 308662 709082 308746 709318
rect 308982 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 52706 708678
rect 52942 708442 53026 708678
rect 53262 708442 88706 708678
rect 88942 708442 89026 708678
rect 89262 708442 124706 708678
rect 124942 708442 125026 708678
rect 125262 708442 160706 708678
rect 160942 708442 161026 708678
rect 161262 708442 196706 708678
rect 196942 708442 197026 708678
rect 197262 708442 232706 708678
rect 232942 708442 233026 708678
rect 233262 708442 268706 708678
rect 268942 708442 269026 708678
rect 269262 708442 304706 708678
rect 304942 708442 305026 708678
rect 305262 708442 340706 708678
rect 340942 708442 341026 708678
rect 341262 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 484706 708678
rect 484942 708442 485026 708678
rect 485262 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 52706 708358
rect 52942 708122 53026 708358
rect 53262 708122 88706 708358
rect 88942 708122 89026 708358
rect 89262 708122 124706 708358
rect 124942 708122 125026 708358
rect 125262 708122 160706 708358
rect 160942 708122 161026 708358
rect 161262 708122 196706 708358
rect 196942 708122 197026 708358
rect 197262 708122 232706 708358
rect 232942 708122 233026 708358
rect 233262 708122 268706 708358
rect 268942 708122 269026 708358
rect 269262 708122 304706 708358
rect 304942 708122 305026 708358
rect 305262 708122 340706 708358
rect 340942 708122 341026 708358
rect 341262 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 484706 708358
rect 484942 708122 485026 708358
rect 485262 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 592650 698294
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 592650 694894
rect -8726 694574 592650 694658
rect -8726 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 592650 694574
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 592650 691174
rect -8726 690854 592650 690938
rect -8726 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 592650 690854
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 315866 677494
rect 316102 677258 316186 677494
rect 316422 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect -8726 677174 592650 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 315866 677174
rect 316102 676938 316186 677174
rect 316422 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 24146 673774
rect 24382 673538 24466 673774
rect 24702 673538 60146 673774
rect 60382 673538 60466 673774
rect 60702 673538 96146 673774
rect 96382 673538 96466 673774
rect 96702 673538 132146 673774
rect 132382 673538 132466 673774
rect 132702 673538 168146 673774
rect 168382 673538 168466 673774
rect 168702 673538 204146 673774
rect 204382 673538 204466 673774
rect 204702 673538 240146 673774
rect 240382 673538 240466 673774
rect 240702 673538 276146 673774
rect 276382 673538 276466 673774
rect 276702 673538 312146 673774
rect 312382 673538 312466 673774
rect 312702 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 592650 673774
rect -8726 673454 592650 673538
rect -8726 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 24146 673454
rect 24382 673218 24466 673454
rect 24702 673218 60146 673454
rect 60382 673218 60466 673454
rect 60702 673218 96146 673454
rect 96382 673218 96466 673454
rect 96702 673218 132146 673454
rect 132382 673218 132466 673454
rect 132702 673218 168146 673454
rect 168382 673218 168466 673454
rect 168702 673218 204146 673454
rect 204382 673218 204466 673454
rect 204702 673218 240146 673454
rect 240382 673218 240466 673454
rect 240702 673218 276146 673454
rect 276382 673218 276466 673454
rect 276702 673218 312146 673454
rect 312382 673218 312466 673454
rect 312702 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 592650 673454
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 56426 670054
rect 56662 669818 56746 670054
rect 56982 669818 92426 670054
rect 92662 669818 92746 670054
rect 92982 669818 128426 670054
rect 128662 669818 128746 670054
rect 128982 669818 164426 670054
rect 164662 669818 164746 670054
rect 164982 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 236426 670054
rect 236662 669818 236746 670054
rect 236982 669818 272426 670054
rect 272662 669818 272746 670054
rect 272982 669818 308426 670054
rect 308662 669818 308746 670054
rect 308982 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 592650 670054
rect -8726 669734 592650 669818
rect -8726 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 56426 669734
rect 56662 669498 56746 669734
rect 56982 669498 92426 669734
rect 92662 669498 92746 669734
rect 92982 669498 128426 669734
rect 128662 669498 128746 669734
rect 128982 669498 164426 669734
rect 164662 669498 164746 669734
rect 164982 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 236426 669734
rect 236662 669498 236746 669734
rect 236982 669498 272426 669734
rect 272662 669498 272746 669734
rect 272982 669498 308426 669734
rect 308662 669498 308746 669734
rect 308982 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 592650 669734
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 52706 666334
rect 52942 666098 53026 666334
rect 53262 666098 88706 666334
rect 88942 666098 89026 666334
rect 89262 666098 124706 666334
rect 124942 666098 125026 666334
rect 125262 666098 160706 666334
rect 160942 666098 161026 666334
rect 161262 666098 196706 666334
rect 196942 666098 197026 666334
rect 197262 666098 232706 666334
rect 232942 666098 233026 666334
rect 233262 666098 268706 666334
rect 268942 666098 269026 666334
rect 269262 666098 304706 666334
rect 304942 666098 305026 666334
rect 305262 666098 340706 666334
rect 340942 666098 341026 666334
rect 341262 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 484706 666334
rect 484942 666098 485026 666334
rect 485262 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 592650 666334
rect -8726 666014 592650 666098
rect -8726 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 52706 666014
rect 52942 665778 53026 666014
rect 53262 665778 88706 666014
rect 88942 665778 89026 666014
rect 89262 665778 124706 666014
rect 124942 665778 125026 666014
rect 125262 665778 160706 666014
rect 160942 665778 161026 666014
rect 161262 665778 196706 666014
rect 196942 665778 197026 666014
rect 197262 665778 232706 666014
rect 232942 665778 233026 666014
rect 233262 665778 268706 666014
rect 268942 665778 269026 666014
rect 269262 665778 304706 666014
rect 304942 665778 305026 666014
rect 305262 665778 340706 666014
rect 340942 665778 341026 666014
rect 341262 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 484706 666014
rect 484942 665778 485026 666014
rect 485262 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 592650 666014
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 592650 662294
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 592650 658894
rect -8726 658574 592650 658658
rect -8726 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 592650 658574
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 592650 655174
rect -8726 654854 592650 654938
rect -8726 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 592650 654854
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 494250 651454
rect 494486 651218 524970 651454
rect 525206 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 494250 651134
rect 494486 650898 524970 651134
rect 525206 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 63866 641494
rect 64102 641258 64186 641494
rect 64422 641258 99866 641494
rect 100102 641258 100186 641494
rect 100422 641258 135866 641494
rect 136102 641258 136186 641494
rect 136422 641258 171866 641494
rect 172102 641258 172186 641494
rect 172422 641258 207866 641494
rect 208102 641258 208186 641494
rect 208422 641258 243866 641494
rect 244102 641258 244186 641494
rect 244422 641258 279866 641494
rect 280102 641258 280186 641494
rect 280422 641258 315866 641494
rect 316102 641258 316186 641494
rect 316422 641258 351866 641494
rect 352102 641258 352186 641494
rect 352422 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 459866 641494
rect 460102 641258 460186 641494
rect 460422 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect -8726 641174 592650 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 63866 641174
rect 64102 640938 64186 641174
rect 64422 640938 99866 641174
rect 100102 640938 100186 641174
rect 100422 640938 135866 641174
rect 136102 640938 136186 641174
rect 136422 640938 171866 641174
rect 172102 640938 172186 641174
rect 172422 640938 207866 641174
rect 208102 640938 208186 641174
rect 208422 640938 243866 641174
rect 244102 640938 244186 641174
rect 244422 640938 279866 641174
rect 280102 640938 280186 641174
rect 280422 640938 315866 641174
rect 316102 640938 316186 641174
rect 316422 640938 351866 641174
rect 352102 640938 352186 641174
rect 352422 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 459866 641174
rect 460102 640938 460186 641174
rect 460422 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 24146 637774
rect 24382 637538 24466 637774
rect 24702 637538 60146 637774
rect 60382 637538 60466 637774
rect 60702 637538 96146 637774
rect 96382 637538 96466 637774
rect 96702 637538 132146 637774
rect 132382 637538 132466 637774
rect 132702 637538 168146 637774
rect 168382 637538 168466 637774
rect 168702 637538 204146 637774
rect 204382 637538 204466 637774
rect 204702 637538 240146 637774
rect 240382 637538 240466 637774
rect 240702 637538 276146 637774
rect 276382 637538 276466 637774
rect 276702 637538 312146 637774
rect 312382 637538 312466 637774
rect 312702 637538 348146 637774
rect 348382 637538 348466 637774
rect 348702 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 492146 637774
rect 492382 637538 492466 637774
rect 492702 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 592650 637774
rect -8726 637454 592650 637538
rect -8726 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 24146 637454
rect 24382 637218 24466 637454
rect 24702 637218 60146 637454
rect 60382 637218 60466 637454
rect 60702 637218 96146 637454
rect 96382 637218 96466 637454
rect 96702 637218 132146 637454
rect 132382 637218 132466 637454
rect 132702 637218 168146 637454
rect 168382 637218 168466 637454
rect 168702 637218 204146 637454
rect 204382 637218 204466 637454
rect 204702 637218 240146 637454
rect 240382 637218 240466 637454
rect 240702 637218 276146 637454
rect 276382 637218 276466 637454
rect 276702 637218 312146 637454
rect 312382 637218 312466 637454
rect 312702 637218 348146 637454
rect 348382 637218 348466 637454
rect 348702 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 492146 637454
rect 492382 637218 492466 637454
rect 492702 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 592650 637454
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 56426 634054
rect 56662 633818 56746 634054
rect 56982 633818 92426 634054
rect 92662 633818 92746 634054
rect 92982 633818 128426 634054
rect 128662 633818 128746 634054
rect 128982 633818 164426 634054
rect 164662 633818 164746 634054
rect 164982 633818 200426 634054
rect 200662 633818 200746 634054
rect 200982 633818 236426 634054
rect 236662 633818 236746 634054
rect 236982 633818 272426 634054
rect 272662 633818 272746 634054
rect 272982 633818 308426 634054
rect 308662 633818 308746 634054
rect 308982 633818 344426 634054
rect 344662 633818 344746 634054
rect 344982 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 488426 634054
rect 488662 633818 488746 634054
rect 488982 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 592650 634054
rect -8726 633734 592650 633818
rect -8726 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 56426 633734
rect 56662 633498 56746 633734
rect 56982 633498 92426 633734
rect 92662 633498 92746 633734
rect 92982 633498 128426 633734
rect 128662 633498 128746 633734
rect 128982 633498 164426 633734
rect 164662 633498 164746 633734
rect 164982 633498 200426 633734
rect 200662 633498 200746 633734
rect 200982 633498 236426 633734
rect 236662 633498 236746 633734
rect 236982 633498 272426 633734
rect 272662 633498 272746 633734
rect 272982 633498 308426 633734
rect 308662 633498 308746 633734
rect 308982 633498 344426 633734
rect 344662 633498 344746 633734
rect 344982 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 488426 633734
rect 488662 633498 488746 633734
rect 488982 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 592650 633734
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 52706 630334
rect 52942 630098 53026 630334
rect 53262 630098 88706 630334
rect 88942 630098 89026 630334
rect 89262 630098 124706 630334
rect 124942 630098 125026 630334
rect 125262 630098 160706 630334
rect 160942 630098 161026 630334
rect 161262 630098 196706 630334
rect 196942 630098 197026 630334
rect 197262 630098 232706 630334
rect 232942 630098 233026 630334
rect 233262 630098 268706 630334
rect 268942 630098 269026 630334
rect 269262 630098 304706 630334
rect 304942 630098 305026 630334
rect 305262 630098 340706 630334
rect 340942 630098 341026 630334
rect 341262 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 484706 630334
rect 484942 630098 485026 630334
rect 485262 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 592650 630334
rect -8726 630014 592650 630098
rect -8726 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 52706 630014
rect 52942 629778 53026 630014
rect 53262 629778 88706 630014
rect 88942 629778 89026 630014
rect 89262 629778 124706 630014
rect 124942 629778 125026 630014
rect 125262 629778 160706 630014
rect 160942 629778 161026 630014
rect 161262 629778 196706 630014
rect 196942 629778 197026 630014
rect 197262 629778 232706 630014
rect 232942 629778 233026 630014
rect 233262 629778 268706 630014
rect 268942 629778 269026 630014
rect 269262 629778 304706 630014
rect 304942 629778 305026 630014
rect 305262 629778 340706 630014
rect 340942 629778 341026 630014
rect 341262 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 484706 630014
rect 484942 629778 485026 630014
rect 485262 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 592650 630014
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 592650 626294
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 592650 622894
rect -8726 622574 592650 622658
rect -8726 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 592650 622574
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 89610 619174
rect 89846 618938 120330 619174
rect 120566 618938 151050 619174
rect 151286 618938 181770 619174
rect 182006 618938 212490 619174
rect 212726 618938 243210 619174
rect 243446 618938 273930 619174
rect 274166 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509610 619174
rect 509846 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 592650 619174
rect -8726 618854 592650 618938
rect -8726 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 89610 618854
rect 89846 618618 120330 618854
rect 120566 618618 151050 618854
rect 151286 618618 181770 618854
rect 182006 618618 212490 618854
rect 212726 618618 243210 618854
rect 243446 618618 273930 618854
rect 274166 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509610 618854
rect 509846 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 592650 618854
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 74250 615454
rect 74486 615218 104970 615454
rect 105206 615218 135690 615454
rect 135926 615218 166410 615454
rect 166646 615218 197130 615454
rect 197366 615218 227850 615454
rect 228086 615218 258570 615454
rect 258806 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 494250 615454
rect 494486 615218 524970 615454
rect 525206 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 74250 615134
rect 74486 614898 104970 615134
rect 105206 614898 135690 615134
rect 135926 614898 166410 615134
rect 166646 614898 197130 615134
rect 197366 614898 227850 615134
rect 228086 614898 258570 615134
rect 258806 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 494250 615134
rect 494486 614898 524970 615134
rect 525206 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 63866 605494
rect 64102 605258 64186 605494
rect 64422 605258 315866 605494
rect 316102 605258 316186 605494
rect 316422 605258 351866 605494
rect 352102 605258 352186 605494
rect 352422 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 459866 605494
rect 460102 605258 460186 605494
rect 460422 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect -8726 605174 592650 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 63866 605174
rect 64102 604938 64186 605174
rect 64422 604938 315866 605174
rect 316102 604938 316186 605174
rect 316422 604938 351866 605174
rect 352102 604938 352186 605174
rect 352422 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 459866 605174
rect 460102 604938 460186 605174
rect 460422 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 24146 601774
rect 24382 601538 24466 601774
rect 24702 601538 60146 601774
rect 60382 601538 60466 601774
rect 60702 601538 312146 601774
rect 312382 601538 312466 601774
rect 312702 601538 348146 601774
rect 348382 601538 348466 601774
rect 348702 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 492146 601774
rect 492382 601538 492466 601774
rect 492702 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 592650 601774
rect -8726 601454 592650 601538
rect -8726 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 24146 601454
rect 24382 601218 24466 601454
rect 24702 601218 60146 601454
rect 60382 601218 60466 601454
rect 60702 601218 312146 601454
rect 312382 601218 312466 601454
rect 312702 601218 348146 601454
rect 348382 601218 348466 601454
rect 348702 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 492146 601454
rect 492382 601218 492466 601454
rect 492702 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 592650 601454
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 56426 598054
rect 56662 597818 56746 598054
rect 56982 597818 308426 598054
rect 308662 597818 308746 598054
rect 308982 597818 344426 598054
rect 344662 597818 344746 598054
rect 344982 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 592650 598054
rect -8726 597734 592650 597818
rect -8726 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 56426 597734
rect 56662 597498 56746 597734
rect 56982 597498 308426 597734
rect 308662 597498 308746 597734
rect 308982 597498 344426 597734
rect 344662 597498 344746 597734
rect 344982 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 592650 597734
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 52706 594334
rect 52942 594098 53026 594334
rect 53262 594098 304706 594334
rect 304942 594098 305026 594334
rect 305262 594098 340706 594334
rect 340942 594098 341026 594334
rect 341262 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 592650 594334
rect -8726 594014 592650 594098
rect -8726 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 52706 594014
rect 52942 593778 53026 594014
rect 53262 593778 304706 594014
rect 304942 593778 305026 594014
rect 305262 593778 340706 594014
rect 340942 593778 341026 594014
rect 341262 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 592650 594014
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 592650 590294
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 592650 586894
rect -8726 586574 592650 586658
rect -8726 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 592650 586574
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 89610 583174
rect 89846 582938 120330 583174
rect 120566 582938 151050 583174
rect 151286 582938 181770 583174
rect 182006 582938 212490 583174
rect 212726 582938 243210 583174
rect 243446 582938 273930 583174
rect 274166 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 592650 583174
rect -8726 582854 592650 582938
rect -8726 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 89610 582854
rect 89846 582618 120330 582854
rect 120566 582618 151050 582854
rect 151286 582618 181770 582854
rect 182006 582618 212490 582854
rect 212726 582618 243210 582854
rect 243446 582618 273930 582854
rect 274166 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 592650 582854
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 74250 579454
rect 74486 579218 104970 579454
rect 105206 579218 135690 579454
rect 135926 579218 166410 579454
rect 166646 579218 197130 579454
rect 197366 579218 227850 579454
rect 228086 579218 258570 579454
rect 258806 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 74250 579134
rect 74486 578898 104970 579134
rect 105206 578898 135690 579134
rect 135926 578898 166410 579134
rect 166646 578898 197130 579134
rect 197366 578898 227850 579134
rect 228086 578898 258570 579134
rect 258806 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 63866 569494
rect 64102 569258 64186 569494
rect 64422 569258 315866 569494
rect 316102 569258 316186 569494
rect 316422 569258 351866 569494
rect 352102 569258 352186 569494
rect 352422 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect -8726 569174 592650 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 63866 569174
rect 64102 568938 64186 569174
rect 64422 568938 315866 569174
rect 316102 568938 316186 569174
rect 316422 568938 351866 569174
rect 352102 568938 352186 569174
rect 352422 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 24146 565774
rect 24382 565538 24466 565774
rect 24702 565538 60146 565774
rect 60382 565538 60466 565774
rect 60702 565538 312146 565774
rect 312382 565538 312466 565774
rect 312702 565538 348146 565774
rect 348382 565538 348466 565774
rect 348702 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 592650 565774
rect -8726 565454 592650 565538
rect -8726 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 24146 565454
rect 24382 565218 24466 565454
rect 24702 565218 60146 565454
rect 60382 565218 60466 565454
rect 60702 565218 312146 565454
rect 312382 565218 312466 565454
rect 312702 565218 348146 565454
rect 348382 565218 348466 565454
rect 348702 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 592650 565454
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 56426 562054
rect 56662 561818 56746 562054
rect 56982 561818 308426 562054
rect 308662 561818 308746 562054
rect 308982 561818 344426 562054
rect 344662 561818 344746 562054
rect 344982 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 592650 562054
rect -8726 561734 592650 561818
rect -8726 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 56426 561734
rect 56662 561498 56746 561734
rect 56982 561498 308426 561734
rect 308662 561498 308746 561734
rect 308982 561498 344426 561734
rect 344662 561498 344746 561734
rect 344982 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 592650 561734
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 52706 558334
rect 52942 558098 53026 558334
rect 53262 558098 304706 558334
rect 304942 558098 305026 558334
rect 305262 558098 340706 558334
rect 340942 558098 341026 558334
rect 341262 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 592650 558334
rect -8726 558014 592650 558098
rect -8726 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 52706 558014
rect 52942 557778 53026 558014
rect 53262 557778 304706 558014
rect 304942 557778 305026 558014
rect 305262 557778 340706 558014
rect 340942 557778 341026 558014
rect 341262 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 592650 558014
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 592650 554294
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 592650 550894
rect -8726 550574 592650 550658
rect -8726 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 592650 550574
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 89610 547174
rect 89846 546938 120330 547174
rect 120566 546938 151050 547174
rect 151286 546938 181770 547174
rect 182006 546938 212490 547174
rect 212726 546938 243210 547174
rect 243446 546938 273930 547174
rect 274166 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 592650 547174
rect -8726 546854 592650 546938
rect -8726 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 89610 546854
rect 89846 546618 120330 546854
rect 120566 546618 151050 546854
rect 151286 546618 181770 546854
rect 182006 546618 212490 546854
rect 212726 546618 243210 546854
rect 243446 546618 273930 546854
rect 274166 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 592650 546854
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 74250 543454
rect 74486 543218 104970 543454
rect 105206 543218 135690 543454
rect 135926 543218 166410 543454
rect 166646 543218 197130 543454
rect 197366 543218 227850 543454
rect 228086 543218 258570 543454
rect 258806 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 74250 543134
rect 74486 542898 104970 543134
rect 105206 542898 135690 543134
rect 135926 542898 166410 543134
rect 166646 542898 197130 543134
rect 197366 542898 227850 543134
rect 228086 542898 258570 543134
rect 258806 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 63866 533494
rect 64102 533258 64186 533494
rect 64422 533258 315866 533494
rect 316102 533258 316186 533494
rect 316422 533258 351866 533494
rect 352102 533258 352186 533494
rect 352422 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect -8726 533174 592650 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 63866 533174
rect 64102 532938 64186 533174
rect 64422 532938 315866 533174
rect 316102 532938 316186 533174
rect 316422 532938 351866 533174
rect 352102 532938 352186 533174
rect 352422 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 24146 529774
rect 24382 529538 24466 529774
rect 24702 529538 60146 529774
rect 60382 529538 60466 529774
rect 60702 529538 312146 529774
rect 312382 529538 312466 529774
rect 312702 529538 348146 529774
rect 348382 529538 348466 529774
rect 348702 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 592650 529774
rect -8726 529454 592650 529538
rect -8726 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 24146 529454
rect 24382 529218 24466 529454
rect 24702 529218 60146 529454
rect 60382 529218 60466 529454
rect 60702 529218 312146 529454
rect 312382 529218 312466 529454
rect 312702 529218 348146 529454
rect 348382 529218 348466 529454
rect 348702 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 592650 529454
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 56426 526054
rect 56662 525818 56746 526054
rect 56982 525818 308426 526054
rect 308662 525818 308746 526054
rect 308982 525818 344426 526054
rect 344662 525818 344746 526054
rect 344982 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 592650 526054
rect -8726 525734 592650 525818
rect -8726 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 56426 525734
rect 56662 525498 56746 525734
rect 56982 525498 308426 525734
rect 308662 525498 308746 525734
rect 308982 525498 344426 525734
rect 344662 525498 344746 525734
rect 344982 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 592650 525734
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 52706 522334
rect 52942 522098 53026 522334
rect 53262 522098 304706 522334
rect 304942 522098 305026 522334
rect 305262 522098 340706 522334
rect 340942 522098 341026 522334
rect 341262 522098 376706 522334
rect 376942 522098 377026 522334
rect 377262 522098 412706 522334
rect 412942 522098 413026 522334
rect 413262 522098 448706 522334
rect 448942 522098 449026 522334
rect 449262 522098 484706 522334
rect 484942 522098 485026 522334
rect 485262 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 592650 522334
rect -8726 522014 592650 522098
rect -8726 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 52706 522014
rect 52942 521778 53026 522014
rect 53262 521778 304706 522014
rect 304942 521778 305026 522014
rect 305262 521778 340706 522014
rect 340942 521778 341026 522014
rect 341262 521778 376706 522014
rect 376942 521778 377026 522014
rect 377262 521778 412706 522014
rect 412942 521778 413026 522014
rect 413262 521778 448706 522014
rect 448942 521778 449026 522014
rect 449262 521778 484706 522014
rect 484942 521778 485026 522014
rect 485262 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 592650 522014
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 592650 518294
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 592650 514894
rect -8726 514574 592650 514658
rect -8726 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 592650 514574
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 89610 511174
rect 89846 510938 120330 511174
rect 120566 510938 151050 511174
rect 151286 510938 181770 511174
rect 182006 510938 212490 511174
rect 212726 510938 243210 511174
rect 243446 510938 273930 511174
rect 274166 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 592650 511174
rect -8726 510854 592650 510938
rect -8726 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 89610 510854
rect 89846 510618 120330 510854
rect 120566 510618 151050 510854
rect 151286 510618 181770 510854
rect 182006 510618 212490 510854
rect 212726 510618 243210 510854
rect 243446 510618 273930 510854
rect 274166 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 592650 510854
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 74250 507454
rect 74486 507218 104970 507454
rect 105206 507218 135690 507454
rect 135926 507218 166410 507454
rect 166646 507218 197130 507454
rect 197366 507218 227850 507454
rect 228086 507218 258570 507454
rect 258806 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 74250 507134
rect 74486 506898 104970 507134
rect 105206 506898 135690 507134
rect 135926 506898 166410 507134
rect 166646 506898 197130 507134
rect 197366 506898 227850 507134
rect 228086 506898 258570 507134
rect 258806 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 63866 497494
rect 64102 497258 64186 497494
rect 64422 497258 315866 497494
rect 316102 497258 316186 497494
rect 316422 497258 351866 497494
rect 352102 497258 352186 497494
rect 352422 497258 387866 497494
rect 388102 497258 388186 497494
rect 388422 497258 423866 497494
rect 424102 497258 424186 497494
rect 424422 497258 459866 497494
rect 460102 497258 460186 497494
rect 460422 497258 495866 497494
rect 496102 497258 496186 497494
rect 496422 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect -8726 497174 592650 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 63866 497174
rect 64102 496938 64186 497174
rect 64422 496938 315866 497174
rect 316102 496938 316186 497174
rect 316422 496938 351866 497174
rect 352102 496938 352186 497174
rect 352422 496938 387866 497174
rect 388102 496938 388186 497174
rect 388422 496938 423866 497174
rect 424102 496938 424186 497174
rect 424422 496938 459866 497174
rect 460102 496938 460186 497174
rect 460422 496938 495866 497174
rect 496102 496938 496186 497174
rect 496422 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 24146 493774
rect 24382 493538 24466 493774
rect 24702 493538 60146 493774
rect 60382 493538 60466 493774
rect 60702 493538 312146 493774
rect 312382 493538 312466 493774
rect 312702 493538 348146 493774
rect 348382 493538 348466 493774
rect 348702 493538 384146 493774
rect 384382 493538 384466 493774
rect 384702 493538 420146 493774
rect 420382 493538 420466 493774
rect 420702 493538 456146 493774
rect 456382 493538 456466 493774
rect 456702 493538 492146 493774
rect 492382 493538 492466 493774
rect 492702 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 592650 493774
rect -8726 493454 592650 493538
rect -8726 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 24146 493454
rect 24382 493218 24466 493454
rect 24702 493218 60146 493454
rect 60382 493218 60466 493454
rect 60702 493218 312146 493454
rect 312382 493218 312466 493454
rect 312702 493218 348146 493454
rect 348382 493218 348466 493454
rect 348702 493218 384146 493454
rect 384382 493218 384466 493454
rect 384702 493218 420146 493454
rect 420382 493218 420466 493454
rect 420702 493218 456146 493454
rect 456382 493218 456466 493454
rect 456702 493218 492146 493454
rect 492382 493218 492466 493454
rect 492702 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 592650 493454
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 56426 490054
rect 56662 489818 56746 490054
rect 56982 489818 308426 490054
rect 308662 489818 308746 490054
rect 308982 489818 344426 490054
rect 344662 489818 344746 490054
rect 344982 489818 380426 490054
rect 380662 489818 380746 490054
rect 380982 489818 416426 490054
rect 416662 489818 416746 490054
rect 416982 489818 452426 490054
rect 452662 489818 452746 490054
rect 452982 489818 488426 490054
rect 488662 489818 488746 490054
rect 488982 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 592650 490054
rect -8726 489734 592650 489818
rect -8726 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 56426 489734
rect 56662 489498 56746 489734
rect 56982 489498 308426 489734
rect 308662 489498 308746 489734
rect 308982 489498 344426 489734
rect 344662 489498 344746 489734
rect 344982 489498 380426 489734
rect 380662 489498 380746 489734
rect 380982 489498 416426 489734
rect 416662 489498 416746 489734
rect 416982 489498 452426 489734
rect 452662 489498 452746 489734
rect 452982 489498 488426 489734
rect 488662 489498 488746 489734
rect 488982 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 592650 489734
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 52706 486334
rect 52942 486098 53026 486334
rect 53262 486098 304706 486334
rect 304942 486098 305026 486334
rect 305262 486098 340706 486334
rect 340942 486098 341026 486334
rect 341262 486098 376706 486334
rect 376942 486098 377026 486334
rect 377262 486098 412706 486334
rect 412942 486098 413026 486334
rect 413262 486098 448706 486334
rect 448942 486098 449026 486334
rect 449262 486098 484706 486334
rect 484942 486098 485026 486334
rect 485262 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 592650 486334
rect -8726 486014 592650 486098
rect -8726 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 52706 486014
rect 52942 485778 53026 486014
rect 53262 485778 304706 486014
rect 304942 485778 305026 486014
rect 305262 485778 340706 486014
rect 340942 485778 341026 486014
rect 341262 485778 376706 486014
rect 376942 485778 377026 486014
rect 377262 485778 412706 486014
rect 412942 485778 413026 486014
rect 413262 485778 448706 486014
rect 448942 485778 449026 486014
rect 449262 485778 484706 486014
rect 484942 485778 485026 486014
rect 485262 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 592650 486014
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 592650 482294
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 592650 478894
rect -8726 478574 592650 478658
rect -8726 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 592650 478574
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 592650 475174
rect -8726 474854 592650 474938
rect -8726 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 592650 474854
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 63866 461494
rect 64102 461258 64186 461494
rect 64422 461258 99866 461494
rect 100102 461258 100186 461494
rect 100422 461258 135866 461494
rect 136102 461258 136186 461494
rect 136422 461258 171866 461494
rect 172102 461258 172186 461494
rect 172422 461258 207866 461494
rect 208102 461258 208186 461494
rect 208422 461258 279866 461494
rect 280102 461258 280186 461494
rect 280422 461258 315866 461494
rect 316102 461258 316186 461494
rect 316422 461258 351866 461494
rect 352102 461258 352186 461494
rect 352422 461258 387866 461494
rect 388102 461258 388186 461494
rect 388422 461258 423866 461494
rect 424102 461258 424186 461494
rect 424422 461258 459866 461494
rect 460102 461258 460186 461494
rect 460422 461258 495866 461494
rect 496102 461258 496186 461494
rect 496422 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect -8726 461174 592650 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 63866 461174
rect 64102 460938 64186 461174
rect 64422 460938 99866 461174
rect 100102 460938 100186 461174
rect 100422 460938 135866 461174
rect 136102 460938 136186 461174
rect 136422 460938 171866 461174
rect 172102 460938 172186 461174
rect 172422 460938 207866 461174
rect 208102 460938 208186 461174
rect 208422 460938 279866 461174
rect 280102 460938 280186 461174
rect 280422 460938 315866 461174
rect 316102 460938 316186 461174
rect 316422 460938 351866 461174
rect 352102 460938 352186 461174
rect 352422 460938 387866 461174
rect 388102 460938 388186 461174
rect 388422 460938 423866 461174
rect 424102 460938 424186 461174
rect 424422 460938 459866 461174
rect 460102 460938 460186 461174
rect 460422 460938 495866 461174
rect 496102 460938 496186 461174
rect 496422 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 24146 457774
rect 24382 457538 24466 457774
rect 24702 457538 60146 457774
rect 60382 457538 60466 457774
rect 60702 457538 96146 457774
rect 96382 457538 96466 457774
rect 96702 457538 132146 457774
rect 132382 457538 132466 457774
rect 132702 457538 168146 457774
rect 168382 457538 168466 457774
rect 168702 457538 204146 457774
rect 204382 457538 204466 457774
rect 204702 457538 240146 457774
rect 240382 457538 240466 457774
rect 240702 457538 276146 457774
rect 276382 457538 276466 457774
rect 276702 457538 312146 457774
rect 312382 457538 312466 457774
rect 312702 457538 348146 457774
rect 348382 457538 348466 457774
rect 348702 457538 384146 457774
rect 384382 457538 384466 457774
rect 384702 457538 420146 457774
rect 420382 457538 420466 457774
rect 420702 457538 456146 457774
rect 456382 457538 456466 457774
rect 456702 457538 492146 457774
rect 492382 457538 492466 457774
rect 492702 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 592650 457774
rect -8726 457454 592650 457538
rect -8726 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 24146 457454
rect 24382 457218 24466 457454
rect 24702 457218 60146 457454
rect 60382 457218 60466 457454
rect 60702 457218 96146 457454
rect 96382 457218 96466 457454
rect 96702 457218 132146 457454
rect 132382 457218 132466 457454
rect 132702 457218 168146 457454
rect 168382 457218 168466 457454
rect 168702 457218 204146 457454
rect 204382 457218 204466 457454
rect 204702 457218 240146 457454
rect 240382 457218 240466 457454
rect 240702 457218 276146 457454
rect 276382 457218 276466 457454
rect 276702 457218 312146 457454
rect 312382 457218 312466 457454
rect 312702 457218 348146 457454
rect 348382 457218 348466 457454
rect 348702 457218 384146 457454
rect 384382 457218 384466 457454
rect 384702 457218 420146 457454
rect 420382 457218 420466 457454
rect 420702 457218 456146 457454
rect 456382 457218 456466 457454
rect 456702 457218 492146 457454
rect 492382 457218 492466 457454
rect 492702 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 592650 457454
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 56426 454054
rect 56662 453818 56746 454054
rect 56982 453818 92426 454054
rect 92662 453818 92746 454054
rect 92982 453818 128426 454054
rect 128662 453818 128746 454054
rect 128982 453818 164426 454054
rect 164662 453818 164746 454054
rect 164982 453818 200426 454054
rect 200662 453818 200746 454054
rect 200982 453818 236426 454054
rect 236662 453818 236746 454054
rect 236982 453818 272426 454054
rect 272662 453818 272746 454054
rect 272982 453818 308426 454054
rect 308662 453818 308746 454054
rect 308982 453818 344426 454054
rect 344662 453818 344746 454054
rect 344982 453818 380426 454054
rect 380662 453818 380746 454054
rect 380982 453818 416426 454054
rect 416662 453818 416746 454054
rect 416982 453818 452426 454054
rect 452662 453818 452746 454054
rect 452982 453818 488426 454054
rect 488662 453818 488746 454054
rect 488982 453818 524426 454054
rect 524662 453818 524746 454054
rect 524982 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 592650 454054
rect -8726 453734 592650 453818
rect -8726 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 56426 453734
rect 56662 453498 56746 453734
rect 56982 453498 92426 453734
rect 92662 453498 92746 453734
rect 92982 453498 128426 453734
rect 128662 453498 128746 453734
rect 128982 453498 164426 453734
rect 164662 453498 164746 453734
rect 164982 453498 200426 453734
rect 200662 453498 200746 453734
rect 200982 453498 236426 453734
rect 236662 453498 236746 453734
rect 236982 453498 272426 453734
rect 272662 453498 272746 453734
rect 272982 453498 308426 453734
rect 308662 453498 308746 453734
rect 308982 453498 344426 453734
rect 344662 453498 344746 453734
rect 344982 453498 380426 453734
rect 380662 453498 380746 453734
rect 380982 453498 416426 453734
rect 416662 453498 416746 453734
rect 416982 453498 452426 453734
rect 452662 453498 452746 453734
rect 452982 453498 488426 453734
rect 488662 453498 488746 453734
rect 488982 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 592650 453734
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 52706 450334
rect 52942 450098 53026 450334
rect 53262 450098 88706 450334
rect 88942 450098 89026 450334
rect 89262 450098 124706 450334
rect 124942 450098 125026 450334
rect 125262 450098 160706 450334
rect 160942 450098 161026 450334
rect 161262 450098 196706 450334
rect 196942 450098 197026 450334
rect 197262 450098 232706 450334
rect 232942 450098 233026 450334
rect 233262 450098 268706 450334
rect 268942 450098 269026 450334
rect 269262 450098 304706 450334
rect 304942 450098 305026 450334
rect 305262 450098 340706 450334
rect 340942 450098 341026 450334
rect 341262 450098 376706 450334
rect 376942 450098 377026 450334
rect 377262 450098 412706 450334
rect 412942 450098 413026 450334
rect 413262 450098 448706 450334
rect 448942 450098 449026 450334
rect 449262 450098 484706 450334
rect 484942 450098 485026 450334
rect 485262 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 592650 450334
rect -8726 450014 592650 450098
rect -8726 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 52706 450014
rect 52942 449778 53026 450014
rect 53262 449778 88706 450014
rect 88942 449778 89026 450014
rect 89262 449778 124706 450014
rect 124942 449778 125026 450014
rect 125262 449778 160706 450014
rect 160942 449778 161026 450014
rect 161262 449778 196706 450014
rect 196942 449778 197026 450014
rect 197262 449778 232706 450014
rect 232942 449778 233026 450014
rect 233262 449778 268706 450014
rect 268942 449778 269026 450014
rect 269262 449778 304706 450014
rect 304942 449778 305026 450014
rect 305262 449778 340706 450014
rect 340942 449778 341026 450014
rect 341262 449778 376706 450014
rect 376942 449778 377026 450014
rect 377262 449778 412706 450014
rect 412942 449778 413026 450014
rect 413262 449778 448706 450014
rect 448942 449778 449026 450014
rect 449262 449778 484706 450014
rect 484942 449778 485026 450014
rect 485262 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 592650 450014
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 592650 446294
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 592650 442894
rect -8726 442574 592650 442658
rect -8726 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 592650 442574
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 592650 439174
rect -8726 438854 592650 438938
rect -8726 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 592650 438854
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 244250 435454
rect 244486 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 274970 435454
rect 275206 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 244250 435134
rect 244486 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 274970 435134
rect 275206 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 63866 425494
rect 64102 425258 64186 425494
rect 64422 425258 99866 425494
rect 100102 425258 100186 425494
rect 100422 425258 135866 425494
rect 136102 425258 136186 425494
rect 136422 425258 171866 425494
rect 172102 425258 172186 425494
rect 172422 425258 207866 425494
rect 208102 425258 208186 425494
rect 208422 425258 279866 425494
rect 280102 425258 280186 425494
rect 280422 425258 315866 425494
rect 316102 425258 316186 425494
rect 316422 425258 351866 425494
rect 352102 425258 352186 425494
rect 352422 425258 387866 425494
rect 388102 425258 388186 425494
rect 388422 425258 423866 425494
rect 424102 425258 424186 425494
rect 424422 425258 459866 425494
rect 460102 425258 460186 425494
rect 460422 425258 495866 425494
rect 496102 425258 496186 425494
rect 496422 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect -8726 425174 592650 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 63866 425174
rect 64102 424938 64186 425174
rect 64422 424938 99866 425174
rect 100102 424938 100186 425174
rect 100422 424938 135866 425174
rect 136102 424938 136186 425174
rect 136422 424938 171866 425174
rect 172102 424938 172186 425174
rect 172422 424938 207866 425174
rect 208102 424938 208186 425174
rect 208422 424938 279866 425174
rect 280102 424938 280186 425174
rect 280422 424938 315866 425174
rect 316102 424938 316186 425174
rect 316422 424938 351866 425174
rect 352102 424938 352186 425174
rect 352422 424938 387866 425174
rect 388102 424938 388186 425174
rect 388422 424938 423866 425174
rect 424102 424938 424186 425174
rect 424422 424938 459866 425174
rect 460102 424938 460186 425174
rect 460422 424938 495866 425174
rect 496102 424938 496186 425174
rect 496422 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 24146 421774
rect 24382 421538 24466 421774
rect 24702 421538 60146 421774
rect 60382 421538 60466 421774
rect 60702 421538 96146 421774
rect 96382 421538 96466 421774
rect 96702 421538 132146 421774
rect 132382 421538 132466 421774
rect 132702 421538 168146 421774
rect 168382 421538 168466 421774
rect 168702 421538 204146 421774
rect 204382 421538 204466 421774
rect 204702 421538 240146 421774
rect 240382 421538 240466 421774
rect 240702 421538 276146 421774
rect 276382 421538 276466 421774
rect 276702 421538 312146 421774
rect 312382 421538 312466 421774
rect 312702 421538 348146 421774
rect 348382 421538 348466 421774
rect 348702 421538 384146 421774
rect 384382 421538 384466 421774
rect 384702 421538 420146 421774
rect 420382 421538 420466 421774
rect 420702 421538 456146 421774
rect 456382 421538 456466 421774
rect 456702 421538 492146 421774
rect 492382 421538 492466 421774
rect 492702 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 592650 421774
rect -8726 421454 592650 421538
rect -8726 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 24146 421454
rect 24382 421218 24466 421454
rect 24702 421218 60146 421454
rect 60382 421218 60466 421454
rect 60702 421218 96146 421454
rect 96382 421218 96466 421454
rect 96702 421218 132146 421454
rect 132382 421218 132466 421454
rect 132702 421218 168146 421454
rect 168382 421218 168466 421454
rect 168702 421218 204146 421454
rect 204382 421218 204466 421454
rect 204702 421218 240146 421454
rect 240382 421218 240466 421454
rect 240702 421218 276146 421454
rect 276382 421218 276466 421454
rect 276702 421218 312146 421454
rect 312382 421218 312466 421454
rect 312702 421218 348146 421454
rect 348382 421218 348466 421454
rect 348702 421218 384146 421454
rect 384382 421218 384466 421454
rect 384702 421218 420146 421454
rect 420382 421218 420466 421454
rect 420702 421218 456146 421454
rect 456382 421218 456466 421454
rect 456702 421218 492146 421454
rect 492382 421218 492466 421454
rect 492702 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 592650 421454
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 56426 418054
rect 56662 417818 56746 418054
rect 56982 417818 92426 418054
rect 92662 417818 92746 418054
rect 92982 417818 128426 418054
rect 128662 417818 128746 418054
rect 128982 417818 164426 418054
rect 164662 417818 164746 418054
rect 164982 417818 200426 418054
rect 200662 417818 200746 418054
rect 200982 417818 236426 418054
rect 236662 417818 236746 418054
rect 236982 417818 272426 418054
rect 272662 417818 272746 418054
rect 272982 417818 308426 418054
rect 308662 417818 308746 418054
rect 308982 417818 344426 418054
rect 344662 417818 344746 418054
rect 344982 417818 380426 418054
rect 380662 417818 380746 418054
rect 380982 417818 416426 418054
rect 416662 417818 416746 418054
rect 416982 417818 452426 418054
rect 452662 417818 452746 418054
rect 452982 417818 488426 418054
rect 488662 417818 488746 418054
rect 488982 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 592650 418054
rect -8726 417734 592650 417818
rect -8726 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 56426 417734
rect 56662 417498 56746 417734
rect 56982 417498 92426 417734
rect 92662 417498 92746 417734
rect 92982 417498 128426 417734
rect 128662 417498 128746 417734
rect 128982 417498 164426 417734
rect 164662 417498 164746 417734
rect 164982 417498 200426 417734
rect 200662 417498 200746 417734
rect 200982 417498 236426 417734
rect 236662 417498 236746 417734
rect 236982 417498 272426 417734
rect 272662 417498 272746 417734
rect 272982 417498 308426 417734
rect 308662 417498 308746 417734
rect 308982 417498 344426 417734
rect 344662 417498 344746 417734
rect 344982 417498 380426 417734
rect 380662 417498 380746 417734
rect 380982 417498 416426 417734
rect 416662 417498 416746 417734
rect 416982 417498 452426 417734
rect 452662 417498 452746 417734
rect 452982 417498 488426 417734
rect 488662 417498 488746 417734
rect 488982 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 592650 417734
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 52706 414334
rect 52942 414098 53026 414334
rect 53262 414098 88706 414334
rect 88942 414098 89026 414334
rect 89262 414098 124706 414334
rect 124942 414098 125026 414334
rect 125262 414098 160706 414334
rect 160942 414098 161026 414334
rect 161262 414098 196706 414334
rect 196942 414098 197026 414334
rect 197262 414098 232706 414334
rect 232942 414098 233026 414334
rect 233262 414098 268706 414334
rect 268942 414098 269026 414334
rect 269262 414098 304706 414334
rect 304942 414098 305026 414334
rect 305262 414098 340706 414334
rect 340942 414098 341026 414334
rect 341262 414098 376706 414334
rect 376942 414098 377026 414334
rect 377262 414098 412706 414334
rect 412942 414098 413026 414334
rect 413262 414098 448706 414334
rect 448942 414098 449026 414334
rect 449262 414098 484706 414334
rect 484942 414098 485026 414334
rect 485262 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 592650 414334
rect -8726 414014 592650 414098
rect -8726 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 52706 414014
rect 52942 413778 53026 414014
rect 53262 413778 88706 414014
rect 88942 413778 89026 414014
rect 89262 413778 124706 414014
rect 124942 413778 125026 414014
rect 125262 413778 160706 414014
rect 160942 413778 161026 414014
rect 161262 413778 196706 414014
rect 196942 413778 197026 414014
rect 197262 413778 232706 414014
rect 232942 413778 233026 414014
rect 233262 413778 268706 414014
rect 268942 413778 269026 414014
rect 269262 413778 304706 414014
rect 304942 413778 305026 414014
rect 305262 413778 340706 414014
rect 340942 413778 341026 414014
rect 341262 413778 376706 414014
rect 376942 413778 377026 414014
rect 377262 413778 412706 414014
rect 412942 413778 413026 414014
rect 413262 413778 448706 414014
rect 448942 413778 449026 414014
rect 449262 413778 484706 414014
rect 484942 413778 485026 414014
rect 485262 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 592650 414014
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 592650 410294
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 592650 406894
rect -8726 406574 592650 406658
rect -8726 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 592650 406574
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 259610 403174
rect 259846 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 592650 403174
rect -8726 402854 592650 402938
rect -8726 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 259610 402854
rect 259846 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 592650 402854
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 109826 399454
rect 110062 399218 110146 399454
rect 110382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 244250 399454
rect 244486 399218 274970 399454
rect 275206 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 109826 399134
rect 110062 398898 110146 399134
rect 110382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 244250 399134
rect 244486 398898 274970 399134
rect 275206 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 63866 389494
rect 64102 389258 64186 389494
rect 64422 389258 99866 389494
rect 100102 389258 100186 389494
rect 100422 389258 135866 389494
rect 136102 389258 136186 389494
rect 136422 389258 171866 389494
rect 172102 389258 172186 389494
rect 172422 389258 207866 389494
rect 208102 389258 208186 389494
rect 208422 389258 279866 389494
rect 280102 389258 280186 389494
rect 280422 389258 315866 389494
rect 316102 389258 316186 389494
rect 316422 389258 351866 389494
rect 352102 389258 352186 389494
rect 352422 389258 387866 389494
rect 388102 389258 388186 389494
rect 388422 389258 423866 389494
rect 424102 389258 424186 389494
rect 424422 389258 459866 389494
rect 460102 389258 460186 389494
rect 460422 389258 495866 389494
rect 496102 389258 496186 389494
rect 496422 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect -8726 389174 592650 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 63866 389174
rect 64102 388938 64186 389174
rect 64422 388938 99866 389174
rect 100102 388938 100186 389174
rect 100422 388938 135866 389174
rect 136102 388938 136186 389174
rect 136422 388938 171866 389174
rect 172102 388938 172186 389174
rect 172422 388938 207866 389174
rect 208102 388938 208186 389174
rect 208422 388938 279866 389174
rect 280102 388938 280186 389174
rect 280422 388938 315866 389174
rect 316102 388938 316186 389174
rect 316422 388938 351866 389174
rect 352102 388938 352186 389174
rect 352422 388938 387866 389174
rect 388102 388938 388186 389174
rect 388422 388938 423866 389174
rect 424102 388938 424186 389174
rect 424422 388938 459866 389174
rect 460102 388938 460186 389174
rect 460422 388938 495866 389174
rect 496102 388938 496186 389174
rect 496422 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 24146 385774
rect 24382 385538 24466 385774
rect 24702 385538 60146 385774
rect 60382 385538 60466 385774
rect 60702 385538 96146 385774
rect 96382 385538 96466 385774
rect 96702 385538 132146 385774
rect 132382 385538 132466 385774
rect 132702 385538 168146 385774
rect 168382 385538 168466 385774
rect 168702 385538 204146 385774
rect 204382 385538 204466 385774
rect 204702 385538 312146 385774
rect 312382 385538 312466 385774
rect 312702 385538 348146 385774
rect 348382 385538 348466 385774
rect 348702 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 492146 385774
rect 492382 385538 492466 385774
rect 492702 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 592650 385774
rect -8726 385454 592650 385538
rect -8726 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 24146 385454
rect 24382 385218 24466 385454
rect 24702 385218 60146 385454
rect 60382 385218 60466 385454
rect 60702 385218 96146 385454
rect 96382 385218 96466 385454
rect 96702 385218 132146 385454
rect 132382 385218 132466 385454
rect 132702 385218 168146 385454
rect 168382 385218 168466 385454
rect 168702 385218 204146 385454
rect 204382 385218 204466 385454
rect 204702 385218 312146 385454
rect 312382 385218 312466 385454
rect 312702 385218 348146 385454
rect 348382 385218 348466 385454
rect 348702 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 492146 385454
rect 492382 385218 492466 385454
rect 492702 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 592650 385454
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 56426 382054
rect 56662 381818 56746 382054
rect 56982 381818 92426 382054
rect 92662 381818 92746 382054
rect 92982 381818 128426 382054
rect 128662 381818 128746 382054
rect 128982 381818 164426 382054
rect 164662 381818 164746 382054
rect 164982 381818 200426 382054
rect 200662 381818 200746 382054
rect 200982 381818 236426 382054
rect 236662 381818 236746 382054
rect 236982 381818 308426 382054
rect 308662 381818 308746 382054
rect 308982 381818 344426 382054
rect 344662 381818 344746 382054
rect 344982 381818 380426 382054
rect 380662 381818 380746 382054
rect 380982 381818 416426 382054
rect 416662 381818 416746 382054
rect 416982 381818 452426 382054
rect 452662 381818 452746 382054
rect 452982 381818 488426 382054
rect 488662 381818 488746 382054
rect 488982 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 592650 382054
rect -8726 381734 592650 381818
rect -8726 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 56426 381734
rect 56662 381498 56746 381734
rect 56982 381498 92426 381734
rect 92662 381498 92746 381734
rect 92982 381498 128426 381734
rect 128662 381498 128746 381734
rect 128982 381498 164426 381734
rect 164662 381498 164746 381734
rect 164982 381498 200426 381734
rect 200662 381498 200746 381734
rect 200982 381498 236426 381734
rect 236662 381498 236746 381734
rect 236982 381498 308426 381734
rect 308662 381498 308746 381734
rect 308982 381498 344426 381734
rect 344662 381498 344746 381734
rect 344982 381498 380426 381734
rect 380662 381498 380746 381734
rect 380982 381498 416426 381734
rect 416662 381498 416746 381734
rect 416982 381498 452426 381734
rect 452662 381498 452746 381734
rect 452982 381498 488426 381734
rect 488662 381498 488746 381734
rect 488982 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 592650 381734
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 52706 378334
rect 52942 378098 53026 378334
rect 53262 378098 88706 378334
rect 88942 378098 89026 378334
rect 89262 378098 124706 378334
rect 124942 378098 125026 378334
rect 125262 378098 160706 378334
rect 160942 378098 161026 378334
rect 161262 378098 196706 378334
rect 196942 378098 197026 378334
rect 197262 378098 232706 378334
rect 232942 378098 233026 378334
rect 233262 378098 304706 378334
rect 304942 378098 305026 378334
rect 305262 378098 340706 378334
rect 340942 378098 341026 378334
rect 341262 378098 376706 378334
rect 376942 378098 377026 378334
rect 377262 378098 412706 378334
rect 412942 378098 413026 378334
rect 413262 378098 448706 378334
rect 448942 378098 449026 378334
rect 449262 378098 484706 378334
rect 484942 378098 485026 378334
rect 485262 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 556706 378334
rect 556942 378098 557026 378334
rect 557262 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 592650 378334
rect -8726 378014 592650 378098
rect -8726 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 52706 378014
rect 52942 377778 53026 378014
rect 53262 377778 88706 378014
rect 88942 377778 89026 378014
rect 89262 377778 124706 378014
rect 124942 377778 125026 378014
rect 125262 377778 160706 378014
rect 160942 377778 161026 378014
rect 161262 377778 196706 378014
rect 196942 377778 197026 378014
rect 197262 377778 232706 378014
rect 232942 377778 233026 378014
rect 233262 377778 304706 378014
rect 304942 377778 305026 378014
rect 305262 377778 340706 378014
rect 340942 377778 341026 378014
rect 341262 377778 376706 378014
rect 376942 377778 377026 378014
rect 377262 377778 412706 378014
rect 412942 377778 413026 378014
rect 413262 377778 448706 378014
rect 448942 377778 449026 378014
rect 449262 377778 484706 378014
rect 484942 377778 485026 378014
rect 485262 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 556706 378014
rect 556942 377778 557026 378014
rect 557262 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 592650 378014
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 592650 374294
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 592650 370894
rect -8726 370574 592650 370658
rect -8726 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 592650 370574
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 259610 367174
rect 259846 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 592650 367174
rect -8726 366854 592650 366938
rect -8726 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 259610 366854
rect 259846 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 592650 366854
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 244250 363454
rect 244486 363218 274970 363454
rect 275206 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 244250 363134
rect 244486 362898 274970 363134
rect 275206 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 63866 353494
rect 64102 353258 64186 353494
rect 64422 353258 99866 353494
rect 100102 353258 100186 353494
rect 100422 353258 135866 353494
rect 136102 353258 136186 353494
rect 136422 353258 171866 353494
rect 172102 353258 172186 353494
rect 172422 353258 207866 353494
rect 208102 353258 208186 353494
rect 208422 353258 279866 353494
rect 280102 353258 280186 353494
rect 280422 353258 315866 353494
rect 316102 353258 316186 353494
rect 316422 353258 351866 353494
rect 352102 353258 352186 353494
rect 352422 353258 387866 353494
rect 388102 353258 388186 353494
rect 388422 353258 423866 353494
rect 424102 353258 424186 353494
rect 424422 353258 459866 353494
rect 460102 353258 460186 353494
rect 460422 353258 495866 353494
rect 496102 353258 496186 353494
rect 496422 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect -8726 353174 592650 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 63866 353174
rect 64102 352938 64186 353174
rect 64422 352938 99866 353174
rect 100102 352938 100186 353174
rect 100422 352938 135866 353174
rect 136102 352938 136186 353174
rect 136422 352938 171866 353174
rect 172102 352938 172186 353174
rect 172422 352938 207866 353174
rect 208102 352938 208186 353174
rect 208422 352938 279866 353174
rect 280102 352938 280186 353174
rect 280422 352938 315866 353174
rect 316102 352938 316186 353174
rect 316422 352938 351866 353174
rect 352102 352938 352186 353174
rect 352422 352938 387866 353174
rect 388102 352938 388186 353174
rect 388422 352938 423866 353174
rect 424102 352938 424186 353174
rect 424422 352938 459866 353174
rect 460102 352938 460186 353174
rect 460422 352938 495866 353174
rect 496102 352938 496186 353174
rect 496422 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 24146 349774
rect 24382 349538 24466 349774
rect 24702 349538 60146 349774
rect 60382 349538 60466 349774
rect 60702 349538 96146 349774
rect 96382 349538 96466 349774
rect 96702 349538 132146 349774
rect 132382 349538 132466 349774
rect 132702 349538 168146 349774
rect 168382 349538 168466 349774
rect 168702 349538 204146 349774
rect 204382 349538 204466 349774
rect 204702 349538 312146 349774
rect 312382 349538 312466 349774
rect 312702 349538 348146 349774
rect 348382 349538 348466 349774
rect 348702 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 456146 349774
rect 456382 349538 456466 349774
rect 456702 349538 492146 349774
rect 492382 349538 492466 349774
rect 492702 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 592650 349774
rect -8726 349454 592650 349538
rect -8726 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 24146 349454
rect 24382 349218 24466 349454
rect 24702 349218 60146 349454
rect 60382 349218 60466 349454
rect 60702 349218 96146 349454
rect 96382 349218 96466 349454
rect 96702 349218 132146 349454
rect 132382 349218 132466 349454
rect 132702 349218 168146 349454
rect 168382 349218 168466 349454
rect 168702 349218 204146 349454
rect 204382 349218 204466 349454
rect 204702 349218 312146 349454
rect 312382 349218 312466 349454
rect 312702 349218 348146 349454
rect 348382 349218 348466 349454
rect 348702 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 456146 349454
rect 456382 349218 456466 349454
rect 456702 349218 492146 349454
rect 492382 349218 492466 349454
rect 492702 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 592650 349454
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 56426 346054
rect 56662 345818 56746 346054
rect 56982 345818 92426 346054
rect 92662 345818 92746 346054
rect 92982 345818 128426 346054
rect 128662 345818 128746 346054
rect 128982 345818 164426 346054
rect 164662 345818 164746 346054
rect 164982 345818 200426 346054
rect 200662 345818 200746 346054
rect 200982 345818 236426 346054
rect 236662 345818 236746 346054
rect 236982 345818 308426 346054
rect 308662 345818 308746 346054
rect 308982 345818 344426 346054
rect 344662 345818 344746 346054
rect 344982 345818 380426 346054
rect 380662 345818 380746 346054
rect 380982 345818 416426 346054
rect 416662 345818 416746 346054
rect 416982 345818 452426 346054
rect 452662 345818 452746 346054
rect 452982 345818 488426 346054
rect 488662 345818 488746 346054
rect 488982 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 592650 346054
rect -8726 345734 592650 345818
rect -8726 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 56426 345734
rect 56662 345498 56746 345734
rect 56982 345498 92426 345734
rect 92662 345498 92746 345734
rect 92982 345498 128426 345734
rect 128662 345498 128746 345734
rect 128982 345498 164426 345734
rect 164662 345498 164746 345734
rect 164982 345498 200426 345734
rect 200662 345498 200746 345734
rect 200982 345498 236426 345734
rect 236662 345498 236746 345734
rect 236982 345498 308426 345734
rect 308662 345498 308746 345734
rect 308982 345498 344426 345734
rect 344662 345498 344746 345734
rect 344982 345498 380426 345734
rect 380662 345498 380746 345734
rect 380982 345498 416426 345734
rect 416662 345498 416746 345734
rect 416982 345498 452426 345734
rect 452662 345498 452746 345734
rect 452982 345498 488426 345734
rect 488662 345498 488746 345734
rect 488982 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 592650 345734
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 52706 342334
rect 52942 342098 53026 342334
rect 53262 342098 88706 342334
rect 88942 342098 89026 342334
rect 89262 342098 124706 342334
rect 124942 342098 125026 342334
rect 125262 342098 160706 342334
rect 160942 342098 161026 342334
rect 161262 342098 196706 342334
rect 196942 342098 197026 342334
rect 197262 342098 232706 342334
rect 232942 342098 233026 342334
rect 233262 342098 304706 342334
rect 304942 342098 305026 342334
rect 305262 342098 340706 342334
rect 340942 342098 341026 342334
rect 341262 342098 376706 342334
rect 376942 342098 377026 342334
rect 377262 342098 412706 342334
rect 412942 342098 413026 342334
rect 413262 342098 448706 342334
rect 448942 342098 449026 342334
rect 449262 342098 484706 342334
rect 484942 342098 485026 342334
rect 485262 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 592650 342334
rect -8726 342014 592650 342098
rect -8726 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 52706 342014
rect 52942 341778 53026 342014
rect 53262 341778 88706 342014
rect 88942 341778 89026 342014
rect 89262 341778 124706 342014
rect 124942 341778 125026 342014
rect 125262 341778 160706 342014
rect 160942 341778 161026 342014
rect 161262 341778 196706 342014
rect 196942 341778 197026 342014
rect 197262 341778 232706 342014
rect 232942 341778 233026 342014
rect 233262 341778 304706 342014
rect 304942 341778 305026 342014
rect 305262 341778 340706 342014
rect 340942 341778 341026 342014
rect 341262 341778 376706 342014
rect 376942 341778 377026 342014
rect 377262 341778 412706 342014
rect 412942 341778 413026 342014
rect 413262 341778 448706 342014
rect 448942 341778 449026 342014
rect 449262 341778 484706 342014
rect 484942 341778 485026 342014
rect 485262 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 592650 342014
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 592650 338294
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 592650 334894
rect -8726 334574 592650 334658
rect -8726 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 592650 334574
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 69610 331174
rect 69846 330938 100330 331174
rect 100566 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 259610 331174
rect 259846 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 592650 331174
rect -8726 330854 592650 330938
rect -8726 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 69610 330854
rect 69846 330618 100330 330854
rect 100566 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 259610 330854
rect 259846 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 592650 330854
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 54250 327454
rect 54486 327218 84970 327454
rect 85206 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 244250 327454
rect 244486 327218 274970 327454
rect 275206 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 54250 327134
rect 54486 326898 84970 327134
rect 85206 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 244250 327134
rect 244486 326898 274970 327134
rect 275206 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 135866 317494
rect 136102 317258 136186 317494
rect 136422 317258 171866 317494
rect 172102 317258 172186 317494
rect 172422 317258 207866 317494
rect 208102 317258 208186 317494
rect 208422 317258 279866 317494
rect 280102 317258 280186 317494
rect 280422 317258 315866 317494
rect 316102 317258 316186 317494
rect 316422 317258 351866 317494
rect 352102 317258 352186 317494
rect 352422 317258 387866 317494
rect 388102 317258 388186 317494
rect 388422 317258 423866 317494
rect 424102 317258 424186 317494
rect 424422 317258 459866 317494
rect 460102 317258 460186 317494
rect 460422 317258 495866 317494
rect 496102 317258 496186 317494
rect 496422 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect -8726 317174 592650 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 135866 317174
rect 136102 316938 136186 317174
rect 136422 316938 171866 317174
rect 172102 316938 172186 317174
rect 172422 316938 207866 317174
rect 208102 316938 208186 317174
rect 208422 316938 279866 317174
rect 280102 316938 280186 317174
rect 280422 316938 315866 317174
rect 316102 316938 316186 317174
rect 316422 316938 351866 317174
rect 352102 316938 352186 317174
rect 352422 316938 387866 317174
rect 388102 316938 388186 317174
rect 388422 316938 423866 317174
rect 424102 316938 424186 317174
rect 424422 316938 459866 317174
rect 460102 316938 460186 317174
rect 460422 316938 495866 317174
rect 496102 316938 496186 317174
rect 496422 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 24146 313774
rect 24382 313538 24466 313774
rect 24702 313538 132146 313774
rect 132382 313538 132466 313774
rect 132702 313538 168146 313774
rect 168382 313538 168466 313774
rect 168702 313538 204146 313774
rect 204382 313538 204466 313774
rect 204702 313538 312146 313774
rect 312382 313538 312466 313774
rect 312702 313538 348146 313774
rect 348382 313538 348466 313774
rect 348702 313538 384146 313774
rect 384382 313538 384466 313774
rect 384702 313538 420146 313774
rect 420382 313538 420466 313774
rect 420702 313538 456146 313774
rect 456382 313538 456466 313774
rect 456702 313538 492146 313774
rect 492382 313538 492466 313774
rect 492702 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 592650 313774
rect -8726 313454 592650 313538
rect -8726 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 24146 313454
rect 24382 313218 24466 313454
rect 24702 313218 132146 313454
rect 132382 313218 132466 313454
rect 132702 313218 168146 313454
rect 168382 313218 168466 313454
rect 168702 313218 204146 313454
rect 204382 313218 204466 313454
rect 204702 313218 312146 313454
rect 312382 313218 312466 313454
rect 312702 313218 348146 313454
rect 348382 313218 348466 313454
rect 348702 313218 384146 313454
rect 384382 313218 384466 313454
rect 384702 313218 420146 313454
rect 420382 313218 420466 313454
rect 420702 313218 456146 313454
rect 456382 313218 456466 313454
rect 456702 313218 492146 313454
rect 492382 313218 492466 313454
rect 492702 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 592650 313454
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 56426 310054
rect 56662 309818 56746 310054
rect 56982 309818 128426 310054
rect 128662 309818 128746 310054
rect 128982 309818 164426 310054
rect 164662 309818 164746 310054
rect 164982 309818 200426 310054
rect 200662 309818 200746 310054
rect 200982 309818 236426 310054
rect 236662 309818 236746 310054
rect 236982 309818 308426 310054
rect 308662 309818 308746 310054
rect 308982 309818 344426 310054
rect 344662 309818 344746 310054
rect 344982 309818 380426 310054
rect 380662 309818 380746 310054
rect 380982 309818 416426 310054
rect 416662 309818 416746 310054
rect 416982 309818 452426 310054
rect 452662 309818 452746 310054
rect 452982 309818 488426 310054
rect 488662 309818 488746 310054
rect 488982 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 592650 310054
rect -8726 309734 592650 309818
rect -8726 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 56426 309734
rect 56662 309498 56746 309734
rect 56982 309498 128426 309734
rect 128662 309498 128746 309734
rect 128982 309498 164426 309734
rect 164662 309498 164746 309734
rect 164982 309498 200426 309734
rect 200662 309498 200746 309734
rect 200982 309498 236426 309734
rect 236662 309498 236746 309734
rect 236982 309498 308426 309734
rect 308662 309498 308746 309734
rect 308982 309498 344426 309734
rect 344662 309498 344746 309734
rect 344982 309498 380426 309734
rect 380662 309498 380746 309734
rect 380982 309498 416426 309734
rect 416662 309498 416746 309734
rect 416982 309498 452426 309734
rect 452662 309498 452746 309734
rect 452982 309498 488426 309734
rect 488662 309498 488746 309734
rect 488982 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 592650 309734
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 52706 306334
rect 52942 306098 53026 306334
rect 53262 306098 124706 306334
rect 124942 306098 125026 306334
rect 125262 306098 160706 306334
rect 160942 306098 161026 306334
rect 161262 306098 196706 306334
rect 196942 306098 197026 306334
rect 197262 306098 232706 306334
rect 232942 306098 233026 306334
rect 233262 306098 304706 306334
rect 304942 306098 305026 306334
rect 305262 306098 340706 306334
rect 340942 306098 341026 306334
rect 341262 306098 376706 306334
rect 376942 306098 377026 306334
rect 377262 306098 412706 306334
rect 412942 306098 413026 306334
rect 413262 306098 448706 306334
rect 448942 306098 449026 306334
rect 449262 306098 484706 306334
rect 484942 306098 485026 306334
rect 485262 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 592650 306334
rect -8726 306014 592650 306098
rect -8726 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 52706 306014
rect 52942 305778 53026 306014
rect 53262 305778 124706 306014
rect 124942 305778 125026 306014
rect 125262 305778 160706 306014
rect 160942 305778 161026 306014
rect 161262 305778 196706 306014
rect 196942 305778 197026 306014
rect 197262 305778 232706 306014
rect 232942 305778 233026 306014
rect 233262 305778 304706 306014
rect 304942 305778 305026 306014
rect 305262 305778 340706 306014
rect 340942 305778 341026 306014
rect 341262 305778 376706 306014
rect 376942 305778 377026 306014
rect 377262 305778 412706 306014
rect 412942 305778 413026 306014
rect 413262 305778 448706 306014
rect 448942 305778 449026 306014
rect 449262 305778 484706 306014
rect 484942 305778 485026 306014
rect 485262 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 592650 306014
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 592650 302294
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 592650 298894
rect -8726 298574 592650 298658
rect -8726 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 592650 298574
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 69610 295174
rect 69846 294938 100330 295174
rect 100566 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 259610 295174
rect 259846 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 592650 295174
rect -8726 294854 592650 294938
rect -8726 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 69610 294854
rect 69846 294618 100330 294854
rect 100566 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 259610 294854
rect 259846 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 592650 294854
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 54250 291454
rect 54486 291218 84970 291454
rect 85206 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 244250 291454
rect 244486 291218 274970 291454
rect 275206 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 54250 291134
rect 54486 290898 84970 291134
rect 85206 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 244250 291134
rect 244486 290898 274970 291134
rect 275206 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 135866 281494
rect 136102 281258 136186 281494
rect 136422 281258 171866 281494
rect 172102 281258 172186 281494
rect 172422 281258 207866 281494
rect 208102 281258 208186 281494
rect 208422 281258 279866 281494
rect 280102 281258 280186 281494
rect 280422 281258 315866 281494
rect 316102 281258 316186 281494
rect 316422 281258 351866 281494
rect 352102 281258 352186 281494
rect 352422 281258 387866 281494
rect 388102 281258 388186 281494
rect 388422 281258 423866 281494
rect 424102 281258 424186 281494
rect 424422 281258 459866 281494
rect 460102 281258 460186 281494
rect 460422 281258 495866 281494
rect 496102 281258 496186 281494
rect 496422 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect -8726 281174 592650 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 135866 281174
rect 136102 280938 136186 281174
rect 136422 280938 171866 281174
rect 172102 280938 172186 281174
rect 172422 280938 207866 281174
rect 208102 280938 208186 281174
rect 208422 280938 279866 281174
rect 280102 280938 280186 281174
rect 280422 280938 315866 281174
rect 316102 280938 316186 281174
rect 316422 280938 351866 281174
rect 352102 280938 352186 281174
rect 352422 280938 387866 281174
rect 388102 280938 388186 281174
rect 388422 280938 423866 281174
rect 424102 280938 424186 281174
rect 424422 280938 459866 281174
rect 460102 280938 460186 281174
rect 460422 280938 495866 281174
rect 496102 280938 496186 281174
rect 496422 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 24146 277774
rect 24382 277538 24466 277774
rect 24702 277538 60146 277774
rect 60382 277538 60466 277774
rect 60702 277538 96146 277774
rect 96382 277538 96466 277774
rect 96702 277538 132146 277774
rect 132382 277538 132466 277774
rect 132702 277538 168146 277774
rect 168382 277538 168466 277774
rect 168702 277538 204146 277774
rect 204382 277538 204466 277774
rect 204702 277538 312146 277774
rect 312382 277538 312466 277774
rect 312702 277538 348146 277774
rect 348382 277538 348466 277774
rect 348702 277538 384146 277774
rect 384382 277538 384466 277774
rect 384702 277538 420146 277774
rect 420382 277538 420466 277774
rect 420702 277538 456146 277774
rect 456382 277538 456466 277774
rect 456702 277538 492146 277774
rect 492382 277538 492466 277774
rect 492702 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 592650 277774
rect -8726 277454 592650 277538
rect -8726 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 24146 277454
rect 24382 277218 24466 277454
rect 24702 277218 60146 277454
rect 60382 277218 60466 277454
rect 60702 277218 96146 277454
rect 96382 277218 96466 277454
rect 96702 277218 132146 277454
rect 132382 277218 132466 277454
rect 132702 277218 168146 277454
rect 168382 277218 168466 277454
rect 168702 277218 204146 277454
rect 204382 277218 204466 277454
rect 204702 277218 312146 277454
rect 312382 277218 312466 277454
rect 312702 277218 348146 277454
rect 348382 277218 348466 277454
rect 348702 277218 384146 277454
rect 384382 277218 384466 277454
rect 384702 277218 420146 277454
rect 420382 277218 420466 277454
rect 420702 277218 456146 277454
rect 456382 277218 456466 277454
rect 456702 277218 492146 277454
rect 492382 277218 492466 277454
rect 492702 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 592650 277454
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 56426 274054
rect 56662 273818 56746 274054
rect 56982 273818 92426 274054
rect 92662 273818 92746 274054
rect 92982 273818 128426 274054
rect 128662 273818 128746 274054
rect 128982 273818 164426 274054
rect 164662 273818 164746 274054
rect 164982 273818 200426 274054
rect 200662 273818 200746 274054
rect 200982 273818 236426 274054
rect 236662 273818 236746 274054
rect 236982 273818 308426 274054
rect 308662 273818 308746 274054
rect 308982 273818 344426 274054
rect 344662 273818 344746 274054
rect 344982 273818 380426 274054
rect 380662 273818 380746 274054
rect 380982 273818 416426 274054
rect 416662 273818 416746 274054
rect 416982 273818 452426 274054
rect 452662 273818 452746 274054
rect 452982 273818 488426 274054
rect 488662 273818 488746 274054
rect 488982 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 592650 274054
rect -8726 273734 592650 273818
rect -8726 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 56426 273734
rect 56662 273498 56746 273734
rect 56982 273498 92426 273734
rect 92662 273498 92746 273734
rect 92982 273498 128426 273734
rect 128662 273498 128746 273734
rect 128982 273498 164426 273734
rect 164662 273498 164746 273734
rect 164982 273498 200426 273734
rect 200662 273498 200746 273734
rect 200982 273498 236426 273734
rect 236662 273498 236746 273734
rect 236982 273498 308426 273734
rect 308662 273498 308746 273734
rect 308982 273498 344426 273734
rect 344662 273498 344746 273734
rect 344982 273498 380426 273734
rect 380662 273498 380746 273734
rect 380982 273498 416426 273734
rect 416662 273498 416746 273734
rect 416982 273498 452426 273734
rect 452662 273498 452746 273734
rect 452982 273498 488426 273734
rect 488662 273498 488746 273734
rect 488982 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 592650 273734
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 52706 270334
rect 52942 270098 53026 270334
rect 53262 270098 88706 270334
rect 88942 270098 89026 270334
rect 89262 270098 124706 270334
rect 124942 270098 125026 270334
rect 125262 270098 160706 270334
rect 160942 270098 161026 270334
rect 161262 270098 196706 270334
rect 196942 270098 197026 270334
rect 197262 270098 232706 270334
rect 232942 270098 233026 270334
rect 233262 270098 304706 270334
rect 304942 270098 305026 270334
rect 305262 270098 340706 270334
rect 340942 270098 341026 270334
rect 341262 270098 376706 270334
rect 376942 270098 377026 270334
rect 377262 270098 412706 270334
rect 412942 270098 413026 270334
rect 413262 270098 448706 270334
rect 448942 270098 449026 270334
rect 449262 270098 484706 270334
rect 484942 270098 485026 270334
rect 485262 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 592650 270334
rect -8726 270014 592650 270098
rect -8726 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 52706 270014
rect 52942 269778 53026 270014
rect 53262 269778 88706 270014
rect 88942 269778 89026 270014
rect 89262 269778 124706 270014
rect 124942 269778 125026 270014
rect 125262 269778 160706 270014
rect 160942 269778 161026 270014
rect 161262 269778 196706 270014
rect 196942 269778 197026 270014
rect 197262 269778 232706 270014
rect 232942 269778 233026 270014
rect 233262 269778 304706 270014
rect 304942 269778 305026 270014
rect 305262 269778 340706 270014
rect 340942 269778 341026 270014
rect 341262 269778 376706 270014
rect 376942 269778 377026 270014
rect 377262 269778 412706 270014
rect 412942 269778 413026 270014
rect 413262 269778 448706 270014
rect 448942 269778 449026 270014
rect 449262 269778 484706 270014
rect 484942 269778 485026 270014
rect 485262 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 592650 270014
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 592650 266294
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 592650 262894
rect -8726 262574 592650 262658
rect -8726 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 592650 262574
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 259610 259174
rect 259846 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 592650 259174
rect -8726 258854 592650 258938
rect -8726 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 259610 258854
rect 259846 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 592650 258854
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 244250 255454
rect 244486 255218 274970 255454
rect 275206 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 244250 255134
rect 244486 254898 274970 255134
rect 275206 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 63866 245494
rect 64102 245258 64186 245494
rect 64422 245258 99866 245494
rect 100102 245258 100186 245494
rect 100422 245258 135866 245494
rect 136102 245258 136186 245494
rect 136422 245258 171866 245494
rect 172102 245258 172186 245494
rect 172422 245258 207866 245494
rect 208102 245258 208186 245494
rect 208422 245258 279866 245494
rect 280102 245258 280186 245494
rect 280422 245258 315866 245494
rect 316102 245258 316186 245494
rect 316422 245258 351866 245494
rect 352102 245258 352186 245494
rect 352422 245258 387866 245494
rect 388102 245258 388186 245494
rect 388422 245258 423866 245494
rect 424102 245258 424186 245494
rect 424422 245258 459866 245494
rect 460102 245258 460186 245494
rect 460422 245258 495866 245494
rect 496102 245258 496186 245494
rect 496422 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect -8726 245174 592650 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 63866 245174
rect 64102 244938 64186 245174
rect 64422 244938 99866 245174
rect 100102 244938 100186 245174
rect 100422 244938 135866 245174
rect 136102 244938 136186 245174
rect 136422 244938 171866 245174
rect 172102 244938 172186 245174
rect 172422 244938 207866 245174
rect 208102 244938 208186 245174
rect 208422 244938 279866 245174
rect 280102 244938 280186 245174
rect 280422 244938 315866 245174
rect 316102 244938 316186 245174
rect 316422 244938 351866 245174
rect 352102 244938 352186 245174
rect 352422 244938 387866 245174
rect 388102 244938 388186 245174
rect 388422 244938 423866 245174
rect 424102 244938 424186 245174
rect 424422 244938 459866 245174
rect 460102 244938 460186 245174
rect 460422 244938 495866 245174
rect 496102 244938 496186 245174
rect 496422 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 24146 241774
rect 24382 241538 24466 241774
rect 24702 241538 60146 241774
rect 60382 241538 60466 241774
rect 60702 241538 96146 241774
rect 96382 241538 96466 241774
rect 96702 241538 132146 241774
rect 132382 241538 132466 241774
rect 132702 241538 168146 241774
rect 168382 241538 168466 241774
rect 168702 241538 204146 241774
rect 204382 241538 204466 241774
rect 204702 241538 312146 241774
rect 312382 241538 312466 241774
rect 312702 241538 348146 241774
rect 348382 241538 348466 241774
rect 348702 241538 384146 241774
rect 384382 241538 384466 241774
rect 384702 241538 420146 241774
rect 420382 241538 420466 241774
rect 420702 241538 456146 241774
rect 456382 241538 456466 241774
rect 456702 241538 492146 241774
rect 492382 241538 492466 241774
rect 492702 241538 528146 241774
rect 528382 241538 528466 241774
rect 528702 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 592650 241774
rect -8726 241454 592650 241538
rect -8726 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 24146 241454
rect 24382 241218 24466 241454
rect 24702 241218 60146 241454
rect 60382 241218 60466 241454
rect 60702 241218 96146 241454
rect 96382 241218 96466 241454
rect 96702 241218 132146 241454
rect 132382 241218 132466 241454
rect 132702 241218 168146 241454
rect 168382 241218 168466 241454
rect 168702 241218 204146 241454
rect 204382 241218 204466 241454
rect 204702 241218 312146 241454
rect 312382 241218 312466 241454
rect 312702 241218 348146 241454
rect 348382 241218 348466 241454
rect 348702 241218 384146 241454
rect 384382 241218 384466 241454
rect 384702 241218 420146 241454
rect 420382 241218 420466 241454
rect 420702 241218 456146 241454
rect 456382 241218 456466 241454
rect 456702 241218 492146 241454
rect 492382 241218 492466 241454
rect 492702 241218 528146 241454
rect 528382 241218 528466 241454
rect 528702 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 592650 241454
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 56426 238054
rect 56662 237818 56746 238054
rect 56982 237818 92426 238054
rect 92662 237818 92746 238054
rect 92982 237818 128426 238054
rect 128662 237818 128746 238054
rect 128982 237818 164426 238054
rect 164662 237818 164746 238054
rect 164982 237818 200426 238054
rect 200662 237818 200746 238054
rect 200982 237818 236426 238054
rect 236662 237818 236746 238054
rect 236982 237818 272426 238054
rect 272662 237818 272746 238054
rect 272982 237818 308426 238054
rect 308662 237818 308746 238054
rect 308982 237818 344426 238054
rect 344662 237818 344746 238054
rect 344982 237818 380426 238054
rect 380662 237818 380746 238054
rect 380982 237818 416426 238054
rect 416662 237818 416746 238054
rect 416982 237818 452426 238054
rect 452662 237818 452746 238054
rect 452982 237818 488426 238054
rect 488662 237818 488746 238054
rect 488982 237818 524426 238054
rect 524662 237818 524746 238054
rect 524982 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 592650 238054
rect -8726 237734 592650 237818
rect -8726 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 56426 237734
rect 56662 237498 56746 237734
rect 56982 237498 92426 237734
rect 92662 237498 92746 237734
rect 92982 237498 128426 237734
rect 128662 237498 128746 237734
rect 128982 237498 164426 237734
rect 164662 237498 164746 237734
rect 164982 237498 200426 237734
rect 200662 237498 200746 237734
rect 200982 237498 236426 237734
rect 236662 237498 236746 237734
rect 236982 237498 272426 237734
rect 272662 237498 272746 237734
rect 272982 237498 308426 237734
rect 308662 237498 308746 237734
rect 308982 237498 344426 237734
rect 344662 237498 344746 237734
rect 344982 237498 380426 237734
rect 380662 237498 380746 237734
rect 380982 237498 416426 237734
rect 416662 237498 416746 237734
rect 416982 237498 452426 237734
rect 452662 237498 452746 237734
rect 452982 237498 488426 237734
rect 488662 237498 488746 237734
rect 488982 237498 524426 237734
rect 524662 237498 524746 237734
rect 524982 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 592650 237734
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 52706 234334
rect 52942 234098 53026 234334
rect 53262 234098 88706 234334
rect 88942 234098 89026 234334
rect 89262 234098 124706 234334
rect 124942 234098 125026 234334
rect 125262 234098 160706 234334
rect 160942 234098 161026 234334
rect 161262 234098 196706 234334
rect 196942 234098 197026 234334
rect 197262 234098 232706 234334
rect 232942 234098 233026 234334
rect 233262 234098 268706 234334
rect 268942 234098 269026 234334
rect 269262 234098 304706 234334
rect 304942 234098 305026 234334
rect 305262 234098 340706 234334
rect 340942 234098 341026 234334
rect 341262 234098 376706 234334
rect 376942 234098 377026 234334
rect 377262 234098 412706 234334
rect 412942 234098 413026 234334
rect 413262 234098 448706 234334
rect 448942 234098 449026 234334
rect 449262 234098 484706 234334
rect 484942 234098 485026 234334
rect 485262 234098 520706 234334
rect 520942 234098 521026 234334
rect 521262 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 592650 234334
rect -8726 234014 592650 234098
rect -8726 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 52706 234014
rect 52942 233778 53026 234014
rect 53262 233778 88706 234014
rect 88942 233778 89026 234014
rect 89262 233778 124706 234014
rect 124942 233778 125026 234014
rect 125262 233778 160706 234014
rect 160942 233778 161026 234014
rect 161262 233778 196706 234014
rect 196942 233778 197026 234014
rect 197262 233778 232706 234014
rect 232942 233778 233026 234014
rect 233262 233778 268706 234014
rect 268942 233778 269026 234014
rect 269262 233778 304706 234014
rect 304942 233778 305026 234014
rect 305262 233778 340706 234014
rect 340942 233778 341026 234014
rect 341262 233778 376706 234014
rect 376942 233778 377026 234014
rect 377262 233778 412706 234014
rect 412942 233778 413026 234014
rect 413262 233778 448706 234014
rect 448942 233778 449026 234014
rect 449262 233778 484706 234014
rect 484942 233778 485026 234014
rect 485262 233778 520706 234014
rect 520942 233778 521026 234014
rect 521262 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 592650 234014
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 592650 230294
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 592650 226894
rect -8726 226574 592650 226658
rect -8726 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 592650 226574
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 592650 223174
rect -8726 222854 592650 222938
rect -8726 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 592650 222854
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 63866 209494
rect 64102 209258 64186 209494
rect 64422 209258 99866 209494
rect 100102 209258 100186 209494
rect 100422 209258 135866 209494
rect 136102 209258 136186 209494
rect 136422 209258 171866 209494
rect 172102 209258 172186 209494
rect 172422 209258 207866 209494
rect 208102 209258 208186 209494
rect 208422 209258 243866 209494
rect 244102 209258 244186 209494
rect 244422 209258 279866 209494
rect 280102 209258 280186 209494
rect 280422 209258 315866 209494
rect 316102 209258 316186 209494
rect 316422 209258 351866 209494
rect 352102 209258 352186 209494
rect 352422 209258 387866 209494
rect 388102 209258 388186 209494
rect 388422 209258 423866 209494
rect 424102 209258 424186 209494
rect 424422 209258 459866 209494
rect 460102 209258 460186 209494
rect 460422 209258 495866 209494
rect 496102 209258 496186 209494
rect 496422 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect -8726 209174 592650 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 63866 209174
rect 64102 208938 64186 209174
rect 64422 208938 99866 209174
rect 100102 208938 100186 209174
rect 100422 208938 135866 209174
rect 136102 208938 136186 209174
rect 136422 208938 171866 209174
rect 172102 208938 172186 209174
rect 172422 208938 207866 209174
rect 208102 208938 208186 209174
rect 208422 208938 243866 209174
rect 244102 208938 244186 209174
rect 244422 208938 279866 209174
rect 280102 208938 280186 209174
rect 280422 208938 315866 209174
rect 316102 208938 316186 209174
rect 316422 208938 351866 209174
rect 352102 208938 352186 209174
rect 352422 208938 387866 209174
rect 388102 208938 388186 209174
rect 388422 208938 423866 209174
rect 424102 208938 424186 209174
rect 424422 208938 459866 209174
rect 460102 208938 460186 209174
rect 460422 208938 495866 209174
rect 496102 208938 496186 209174
rect 496422 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 24146 205774
rect 24382 205538 24466 205774
rect 24702 205538 60146 205774
rect 60382 205538 60466 205774
rect 60702 205538 96146 205774
rect 96382 205538 96466 205774
rect 96702 205538 132146 205774
rect 132382 205538 132466 205774
rect 132702 205538 168146 205774
rect 168382 205538 168466 205774
rect 168702 205538 204146 205774
rect 204382 205538 204466 205774
rect 204702 205538 240146 205774
rect 240382 205538 240466 205774
rect 240702 205538 276146 205774
rect 276382 205538 276466 205774
rect 276702 205538 312146 205774
rect 312382 205538 312466 205774
rect 312702 205538 348146 205774
rect 348382 205538 348466 205774
rect 348702 205538 384146 205774
rect 384382 205538 384466 205774
rect 384702 205538 420146 205774
rect 420382 205538 420466 205774
rect 420702 205538 456146 205774
rect 456382 205538 456466 205774
rect 456702 205538 492146 205774
rect 492382 205538 492466 205774
rect 492702 205538 528146 205774
rect 528382 205538 528466 205774
rect 528702 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 592650 205774
rect -8726 205454 592650 205538
rect -8726 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 24146 205454
rect 24382 205218 24466 205454
rect 24702 205218 60146 205454
rect 60382 205218 60466 205454
rect 60702 205218 96146 205454
rect 96382 205218 96466 205454
rect 96702 205218 132146 205454
rect 132382 205218 132466 205454
rect 132702 205218 168146 205454
rect 168382 205218 168466 205454
rect 168702 205218 204146 205454
rect 204382 205218 204466 205454
rect 204702 205218 240146 205454
rect 240382 205218 240466 205454
rect 240702 205218 276146 205454
rect 276382 205218 276466 205454
rect 276702 205218 312146 205454
rect 312382 205218 312466 205454
rect 312702 205218 348146 205454
rect 348382 205218 348466 205454
rect 348702 205218 384146 205454
rect 384382 205218 384466 205454
rect 384702 205218 420146 205454
rect 420382 205218 420466 205454
rect 420702 205218 456146 205454
rect 456382 205218 456466 205454
rect 456702 205218 492146 205454
rect 492382 205218 492466 205454
rect 492702 205218 528146 205454
rect 528382 205218 528466 205454
rect 528702 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 592650 205454
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 56426 202054
rect 56662 201818 56746 202054
rect 56982 201818 92426 202054
rect 92662 201818 92746 202054
rect 92982 201818 128426 202054
rect 128662 201818 128746 202054
rect 128982 201818 164426 202054
rect 164662 201818 164746 202054
rect 164982 201818 200426 202054
rect 200662 201818 200746 202054
rect 200982 201818 236426 202054
rect 236662 201818 236746 202054
rect 236982 201818 272426 202054
rect 272662 201818 272746 202054
rect 272982 201818 308426 202054
rect 308662 201818 308746 202054
rect 308982 201818 344426 202054
rect 344662 201818 344746 202054
rect 344982 201818 380426 202054
rect 380662 201818 380746 202054
rect 380982 201818 416426 202054
rect 416662 201818 416746 202054
rect 416982 201818 452426 202054
rect 452662 201818 452746 202054
rect 452982 201818 488426 202054
rect 488662 201818 488746 202054
rect 488982 201818 524426 202054
rect 524662 201818 524746 202054
rect 524982 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 592650 202054
rect -8726 201734 592650 201818
rect -8726 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 56426 201734
rect 56662 201498 56746 201734
rect 56982 201498 92426 201734
rect 92662 201498 92746 201734
rect 92982 201498 128426 201734
rect 128662 201498 128746 201734
rect 128982 201498 164426 201734
rect 164662 201498 164746 201734
rect 164982 201498 200426 201734
rect 200662 201498 200746 201734
rect 200982 201498 236426 201734
rect 236662 201498 236746 201734
rect 236982 201498 272426 201734
rect 272662 201498 272746 201734
rect 272982 201498 308426 201734
rect 308662 201498 308746 201734
rect 308982 201498 344426 201734
rect 344662 201498 344746 201734
rect 344982 201498 380426 201734
rect 380662 201498 380746 201734
rect 380982 201498 416426 201734
rect 416662 201498 416746 201734
rect 416982 201498 452426 201734
rect 452662 201498 452746 201734
rect 452982 201498 488426 201734
rect 488662 201498 488746 201734
rect 488982 201498 524426 201734
rect 524662 201498 524746 201734
rect 524982 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 592650 201734
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 52706 198334
rect 52942 198098 53026 198334
rect 53262 198098 88706 198334
rect 88942 198098 89026 198334
rect 89262 198098 124706 198334
rect 124942 198098 125026 198334
rect 125262 198098 160706 198334
rect 160942 198098 161026 198334
rect 161262 198098 196706 198334
rect 196942 198098 197026 198334
rect 197262 198098 232706 198334
rect 232942 198098 233026 198334
rect 233262 198098 268706 198334
rect 268942 198098 269026 198334
rect 269262 198098 304706 198334
rect 304942 198098 305026 198334
rect 305262 198098 340706 198334
rect 340942 198098 341026 198334
rect 341262 198098 376706 198334
rect 376942 198098 377026 198334
rect 377262 198098 412706 198334
rect 412942 198098 413026 198334
rect 413262 198098 448706 198334
rect 448942 198098 449026 198334
rect 449262 198098 484706 198334
rect 484942 198098 485026 198334
rect 485262 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 592650 198334
rect -8726 198014 592650 198098
rect -8726 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 52706 198014
rect 52942 197778 53026 198014
rect 53262 197778 88706 198014
rect 88942 197778 89026 198014
rect 89262 197778 124706 198014
rect 124942 197778 125026 198014
rect 125262 197778 160706 198014
rect 160942 197778 161026 198014
rect 161262 197778 196706 198014
rect 196942 197778 197026 198014
rect 197262 197778 232706 198014
rect 232942 197778 233026 198014
rect 233262 197778 268706 198014
rect 268942 197778 269026 198014
rect 269262 197778 304706 198014
rect 304942 197778 305026 198014
rect 305262 197778 340706 198014
rect 340942 197778 341026 198014
rect 341262 197778 376706 198014
rect 376942 197778 377026 198014
rect 377262 197778 412706 198014
rect 412942 197778 413026 198014
rect 413262 197778 448706 198014
rect 448942 197778 449026 198014
rect 449262 197778 484706 198014
rect 484942 197778 485026 198014
rect 485262 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 592650 198014
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 592650 194294
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 592650 190894
rect -8726 190574 592650 190658
rect -8726 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 592650 190574
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 592650 187174
rect -8726 186854 592650 186938
rect -8726 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 592650 186854
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 63866 173494
rect 64102 173258 64186 173494
rect 64422 173258 99866 173494
rect 100102 173258 100186 173494
rect 100422 173258 135866 173494
rect 136102 173258 136186 173494
rect 136422 173258 171866 173494
rect 172102 173258 172186 173494
rect 172422 173258 207866 173494
rect 208102 173258 208186 173494
rect 208422 173258 243866 173494
rect 244102 173258 244186 173494
rect 244422 173258 279866 173494
rect 280102 173258 280186 173494
rect 280422 173258 315866 173494
rect 316102 173258 316186 173494
rect 316422 173258 351866 173494
rect 352102 173258 352186 173494
rect 352422 173258 387866 173494
rect 388102 173258 388186 173494
rect 388422 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 495866 173494
rect 496102 173258 496186 173494
rect 496422 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect -8726 173174 592650 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 63866 173174
rect 64102 172938 64186 173174
rect 64422 172938 99866 173174
rect 100102 172938 100186 173174
rect 100422 172938 135866 173174
rect 136102 172938 136186 173174
rect 136422 172938 171866 173174
rect 172102 172938 172186 173174
rect 172422 172938 207866 173174
rect 208102 172938 208186 173174
rect 208422 172938 243866 173174
rect 244102 172938 244186 173174
rect 244422 172938 279866 173174
rect 280102 172938 280186 173174
rect 280422 172938 315866 173174
rect 316102 172938 316186 173174
rect 316422 172938 351866 173174
rect 352102 172938 352186 173174
rect 352422 172938 387866 173174
rect 388102 172938 388186 173174
rect 388422 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 495866 173174
rect 496102 172938 496186 173174
rect 496422 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 24146 169774
rect 24382 169538 24466 169774
rect 24702 169538 60146 169774
rect 60382 169538 60466 169774
rect 60702 169538 96146 169774
rect 96382 169538 96466 169774
rect 96702 169538 132146 169774
rect 132382 169538 132466 169774
rect 132702 169538 168146 169774
rect 168382 169538 168466 169774
rect 168702 169538 204146 169774
rect 204382 169538 204466 169774
rect 204702 169538 240146 169774
rect 240382 169538 240466 169774
rect 240702 169538 276146 169774
rect 276382 169538 276466 169774
rect 276702 169538 312146 169774
rect 312382 169538 312466 169774
rect 312702 169538 348146 169774
rect 348382 169538 348466 169774
rect 348702 169538 384146 169774
rect 384382 169538 384466 169774
rect 384702 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 492146 169774
rect 492382 169538 492466 169774
rect 492702 169538 528146 169774
rect 528382 169538 528466 169774
rect 528702 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 592650 169774
rect -8726 169454 592650 169538
rect -8726 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 24146 169454
rect 24382 169218 24466 169454
rect 24702 169218 60146 169454
rect 60382 169218 60466 169454
rect 60702 169218 96146 169454
rect 96382 169218 96466 169454
rect 96702 169218 132146 169454
rect 132382 169218 132466 169454
rect 132702 169218 168146 169454
rect 168382 169218 168466 169454
rect 168702 169218 204146 169454
rect 204382 169218 204466 169454
rect 204702 169218 240146 169454
rect 240382 169218 240466 169454
rect 240702 169218 276146 169454
rect 276382 169218 276466 169454
rect 276702 169218 312146 169454
rect 312382 169218 312466 169454
rect 312702 169218 348146 169454
rect 348382 169218 348466 169454
rect 348702 169218 384146 169454
rect 384382 169218 384466 169454
rect 384702 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 492146 169454
rect 492382 169218 492466 169454
rect 492702 169218 528146 169454
rect 528382 169218 528466 169454
rect 528702 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 592650 169454
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 56426 166054
rect 56662 165818 56746 166054
rect 56982 165818 92426 166054
rect 92662 165818 92746 166054
rect 92982 165818 128426 166054
rect 128662 165818 128746 166054
rect 128982 165818 164426 166054
rect 164662 165818 164746 166054
rect 164982 165818 200426 166054
rect 200662 165818 200746 166054
rect 200982 165818 236426 166054
rect 236662 165818 236746 166054
rect 236982 165818 272426 166054
rect 272662 165818 272746 166054
rect 272982 165818 308426 166054
rect 308662 165818 308746 166054
rect 308982 165818 344426 166054
rect 344662 165818 344746 166054
rect 344982 165818 380426 166054
rect 380662 165818 380746 166054
rect 380982 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 592650 166054
rect -8726 165734 592650 165818
rect -8726 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 56426 165734
rect 56662 165498 56746 165734
rect 56982 165498 92426 165734
rect 92662 165498 92746 165734
rect 92982 165498 128426 165734
rect 128662 165498 128746 165734
rect 128982 165498 164426 165734
rect 164662 165498 164746 165734
rect 164982 165498 200426 165734
rect 200662 165498 200746 165734
rect 200982 165498 236426 165734
rect 236662 165498 236746 165734
rect 236982 165498 272426 165734
rect 272662 165498 272746 165734
rect 272982 165498 308426 165734
rect 308662 165498 308746 165734
rect 308982 165498 344426 165734
rect 344662 165498 344746 165734
rect 344982 165498 380426 165734
rect 380662 165498 380746 165734
rect 380982 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 592650 165734
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 52706 162334
rect 52942 162098 53026 162334
rect 53262 162098 88706 162334
rect 88942 162098 89026 162334
rect 89262 162098 124706 162334
rect 124942 162098 125026 162334
rect 125262 162098 160706 162334
rect 160942 162098 161026 162334
rect 161262 162098 196706 162334
rect 196942 162098 197026 162334
rect 197262 162098 232706 162334
rect 232942 162098 233026 162334
rect 233262 162098 268706 162334
rect 268942 162098 269026 162334
rect 269262 162098 304706 162334
rect 304942 162098 305026 162334
rect 305262 162098 340706 162334
rect 340942 162098 341026 162334
rect 341262 162098 376706 162334
rect 376942 162098 377026 162334
rect 377262 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 592650 162334
rect -8726 162014 592650 162098
rect -8726 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 52706 162014
rect 52942 161778 53026 162014
rect 53262 161778 88706 162014
rect 88942 161778 89026 162014
rect 89262 161778 124706 162014
rect 124942 161778 125026 162014
rect 125262 161778 160706 162014
rect 160942 161778 161026 162014
rect 161262 161778 196706 162014
rect 196942 161778 197026 162014
rect 197262 161778 232706 162014
rect 232942 161778 233026 162014
rect 233262 161778 268706 162014
rect 268942 161778 269026 162014
rect 269262 161778 304706 162014
rect 304942 161778 305026 162014
rect 305262 161778 340706 162014
rect 340942 161778 341026 162014
rect 341262 161778 376706 162014
rect 376942 161778 377026 162014
rect 377262 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 592650 162014
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 592650 158294
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 592650 154894
rect -8726 154574 592650 154658
rect -8726 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 592650 154574
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 592650 151174
rect -8726 150854 592650 150938
rect -8726 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 592650 150854
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 63866 137494
rect 64102 137258 64186 137494
rect 64422 137258 99866 137494
rect 100102 137258 100186 137494
rect 100422 137258 135866 137494
rect 136102 137258 136186 137494
rect 136422 137258 171866 137494
rect 172102 137258 172186 137494
rect 172422 137258 207866 137494
rect 208102 137258 208186 137494
rect 208422 137258 243866 137494
rect 244102 137258 244186 137494
rect 244422 137258 279866 137494
rect 280102 137258 280186 137494
rect 280422 137258 315866 137494
rect 316102 137258 316186 137494
rect 316422 137258 351866 137494
rect 352102 137258 352186 137494
rect 352422 137258 387866 137494
rect 388102 137258 388186 137494
rect 388422 137258 423866 137494
rect 424102 137258 424186 137494
rect 424422 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 495866 137494
rect 496102 137258 496186 137494
rect 496422 137258 531866 137494
rect 532102 137258 532186 137494
rect 532422 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect -8726 137174 592650 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 63866 137174
rect 64102 136938 64186 137174
rect 64422 136938 99866 137174
rect 100102 136938 100186 137174
rect 100422 136938 135866 137174
rect 136102 136938 136186 137174
rect 136422 136938 171866 137174
rect 172102 136938 172186 137174
rect 172422 136938 207866 137174
rect 208102 136938 208186 137174
rect 208422 136938 243866 137174
rect 244102 136938 244186 137174
rect 244422 136938 279866 137174
rect 280102 136938 280186 137174
rect 280422 136938 315866 137174
rect 316102 136938 316186 137174
rect 316422 136938 351866 137174
rect 352102 136938 352186 137174
rect 352422 136938 387866 137174
rect 388102 136938 388186 137174
rect 388422 136938 423866 137174
rect 424102 136938 424186 137174
rect 424422 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 495866 137174
rect 496102 136938 496186 137174
rect 496422 136938 531866 137174
rect 532102 136938 532186 137174
rect 532422 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 24146 133774
rect 24382 133538 24466 133774
rect 24702 133538 60146 133774
rect 60382 133538 60466 133774
rect 60702 133538 96146 133774
rect 96382 133538 96466 133774
rect 96702 133538 132146 133774
rect 132382 133538 132466 133774
rect 132702 133538 168146 133774
rect 168382 133538 168466 133774
rect 168702 133538 204146 133774
rect 204382 133538 204466 133774
rect 204702 133538 240146 133774
rect 240382 133538 240466 133774
rect 240702 133538 276146 133774
rect 276382 133538 276466 133774
rect 276702 133538 312146 133774
rect 312382 133538 312466 133774
rect 312702 133538 348146 133774
rect 348382 133538 348466 133774
rect 348702 133538 384146 133774
rect 384382 133538 384466 133774
rect 384702 133538 420146 133774
rect 420382 133538 420466 133774
rect 420702 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 492146 133774
rect 492382 133538 492466 133774
rect 492702 133538 528146 133774
rect 528382 133538 528466 133774
rect 528702 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 592650 133774
rect -8726 133454 592650 133538
rect -8726 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 24146 133454
rect 24382 133218 24466 133454
rect 24702 133218 60146 133454
rect 60382 133218 60466 133454
rect 60702 133218 96146 133454
rect 96382 133218 96466 133454
rect 96702 133218 132146 133454
rect 132382 133218 132466 133454
rect 132702 133218 168146 133454
rect 168382 133218 168466 133454
rect 168702 133218 204146 133454
rect 204382 133218 204466 133454
rect 204702 133218 240146 133454
rect 240382 133218 240466 133454
rect 240702 133218 276146 133454
rect 276382 133218 276466 133454
rect 276702 133218 312146 133454
rect 312382 133218 312466 133454
rect 312702 133218 348146 133454
rect 348382 133218 348466 133454
rect 348702 133218 384146 133454
rect 384382 133218 384466 133454
rect 384702 133218 420146 133454
rect 420382 133218 420466 133454
rect 420702 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 492146 133454
rect 492382 133218 492466 133454
rect 492702 133218 528146 133454
rect 528382 133218 528466 133454
rect 528702 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 592650 133454
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 56426 130054
rect 56662 129818 56746 130054
rect 56982 129818 92426 130054
rect 92662 129818 92746 130054
rect 92982 129818 128426 130054
rect 128662 129818 128746 130054
rect 128982 129818 164426 130054
rect 164662 129818 164746 130054
rect 164982 129818 200426 130054
rect 200662 129818 200746 130054
rect 200982 129818 236426 130054
rect 236662 129818 236746 130054
rect 236982 129818 272426 130054
rect 272662 129818 272746 130054
rect 272982 129818 308426 130054
rect 308662 129818 308746 130054
rect 308982 129818 344426 130054
rect 344662 129818 344746 130054
rect 344982 129818 380426 130054
rect 380662 129818 380746 130054
rect 380982 129818 416426 130054
rect 416662 129818 416746 130054
rect 416982 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 488426 130054
rect 488662 129818 488746 130054
rect 488982 129818 524426 130054
rect 524662 129818 524746 130054
rect 524982 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 592650 130054
rect -8726 129734 592650 129818
rect -8726 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 56426 129734
rect 56662 129498 56746 129734
rect 56982 129498 92426 129734
rect 92662 129498 92746 129734
rect 92982 129498 128426 129734
rect 128662 129498 128746 129734
rect 128982 129498 164426 129734
rect 164662 129498 164746 129734
rect 164982 129498 200426 129734
rect 200662 129498 200746 129734
rect 200982 129498 236426 129734
rect 236662 129498 236746 129734
rect 236982 129498 272426 129734
rect 272662 129498 272746 129734
rect 272982 129498 308426 129734
rect 308662 129498 308746 129734
rect 308982 129498 344426 129734
rect 344662 129498 344746 129734
rect 344982 129498 380426 129734
rect 380662 129498 380746 129734
rect 380982 129498 416426 129734
rect 416662 129498 416746 129734
rect 416982 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 488426 129734
rect 488662 129498 488746 129734
rect 488982 129498 524426 129734
rect 524662 129498 524746 129734
rect 524982 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 592650 129734
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 52706 126334
rect 52942 126098 53026 126334
rect 53262 126098 88706 126334
rect 88942 126098 89026 126334
rect 89262 126098 124706 126334
rect 124942 126098 125026 126334
rect 125262 126098 160706 126334
rect 160942 126098 161026 126334
rect 161262 126098 196706 126334
rect 196942 126098 197026 126334
rect 197262 126098 232706 126334
rect 232942 126098 233026 126334
rect 233262 126098 268706 126334
rect 268942 126098 269026 126334
rect 269262 126098 304706 126334
rect 304942 126098 305026 126334
rect 305262 126098 340706 126334
rect 340942 126098 341026 126334
rect 341262 126098 376706 126334
rect 376942 126098 377026 126334
rect 377262 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 520706 126334
rect 520942 126098 521026 126334
rect 521262 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 592650 126334
rect -8726 126014 592650 126098
rect -8726 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 52706 126014
rect 52942 125778 53026 126014
rect 53262 125778 88706 126014
rect 88942 125778 89026 126014
rect 89262 125778 124706 126014
rect 124942 125778 125026 126014
rect 125262 125778 160706 126014
rect 160942 125778 161026 126014
rect 161262 125778 196706 126014
rect 196942 125778 197026 126014
rect 197262 125778 232706 126014
rect 232942 125778 233026 126014
rect 233262 125778 268706 126014
rect 268942 125778 269026 126014
rect 269262 125778 304706 126014
rect 304942 125778 305026 126014
rect 305262 125778 340706 126014
rect 340942 125778 341026 126014
rect 341262 125778 376706 126014
rect 376942 125778 377026 126014
rect 377262 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 520706 126014
rect 520942 125778 521026 126014
rect 521262 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 592650 126014
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 592650 122294
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 592650 118894
rect -8726 118574 592650 118658
rect -8726 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 592650 118574
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 592650 115174
rect -8726 114854 592650 114938
rect -8726 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 592650 114854
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 63866 101494
rect 64102 101258 64186 101494
rect 64422 101258 99866 101494
rect 100102 101258 100186 101494
rect 100422 101258 135866 101494
rect 136102 101258 136186 101494
rect 136422 101258 171866 101494
rect 172102 101258 172186 101494
rect 172422 101258 207866 101494
rect 208102 101258 208186 101494
rect 208422 101258 243866 101494
rect 244102 101258 244186 101494
rect 244422 101258 279866 101494
rect 280102 101258 280186 101494
rect 280422 101258 315866 101494
rect 316102 101258 316186 101494
rect 316422 101258 351866 101494
rect 352102 101258 352186 101494
rect 352422 101258 387866 101494
rect 388102 101258 388186 101494
rect 388422 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 495866 101494
rect 496102 101258 496186 101494
rect 496422 101258 531866 101494
rect 532102 101258 532186 101494
rect 532422 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect -8726 101174 592650 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 63866 101174
rect 64102 100938 64186 101174
rect 64422 100938 99866 101174
rect 100102 100938 100186 101174
rect 100422 100938 135866 101174
rect 136102 100938 136186 101174
rect 136422 100938 171866 101174
rect 172102 100938 172186 101174
rect 172422 100938 207866 101174
rect 208102 100938 208186 101174
rect 208422 100938 243866 101174
rect 244102 100938 244186 101174
rect 244422 100938 279866 101174
rect 280102 100938 280186 101174
rect 280422 100938 315866 101174
rect 316102 100938 316186 101174
rect 316422 100938 351866 101174
rect 352102 100938 352186 101174
rect 352422 100938 387866 101174
rect 388102 100938 388186 101174
rect 388422 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 495866 101174
rect 496102 100938 496186 101174
rect 496422 100938 531866 101174
rect 532102 100938 532186 101174
rect 532422 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 24146 97774
rect 24382 97538 24466 97774
rect 24702 97538 60146 97774
rect 60382 97538 60466 97774
rect 60702 97538 96146 97774
rect 96382 97538 96466 97774
rect 96702 97538 132146 97774
rect 132382 97538 132466 97774
rect 132702 97538 168146 97774
rect 168382 97538 168466 97774
rect 168702 97538 204146 97774
rect 204382 97538 204466 97774
rect 204702 97538 240146 97774
rect 240382 97538 240466 97774
rect 240702 97538 276146 97774
rect 276382 97538 276466 97774
rect 276702 97538 312146 97774
rect 312382 97538 312466 97774
rect 312702 97538 348146 97774
rect 348382 97538 348466 97774
rect 348702 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 492146 97774
rect 492382 97538 492466 97774
rect 492702 97538 528146 97774
rect 528382 97538 528466 97774
rect 528702 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 592650 97774
rect -8726 97454 592650 97538
rect -8726 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 24146 97454
rect 24382 97218 24466 97454
rect 24702 97218 60146 97454
rect 60382 97218 60466 97454
rect 60702 97218 96146 97454
rect 96382 97218 96466 97454
rect 96702 97218 132146 97454
rect 132382 97218 132466 97454
rect 132702 97218 168146 97454
rect 168382 97218 168466 97454
rect 168702 97218 204146 97454
rect 204382 97218 204466 97454
rect 204702 97218 240146 97454
rect 240382 97218 240466 97454
rect 240702 97218 276146 97454
rect 276382 97218 276466 97454
rect 276702 97218 312146 97454
rect 312382 97218 312466 97454
rect 312702 97218 348146 97454
rect 348382 97218 348466 97454
rect 348702 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 492146 97454
rect 492382 97218 492466 97454
rect 492702 97218 528146 97454
rect 528382 97218 528466 97454
rect 528702 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 592650 97454
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 56426 94054
rect 56662 93818 56746 94054
rect 56982 93818 92426 94054
rect 92662 93818 92746 94054
rect 92982 93818 128426 94054
rect 128662 93818 128746 94054
rect 128982 93818 164426 94054
rect 164662 93818 164746 94054
rect 164982 93818 200426 94054
rect 200662 93818 200746 94054
rect 200982 93818 236426 94054
rect 236662 93818 236746 94054
rect 236982 93818 272426 94054
rect 272662 93818 272746 94054
rect 272982 93818 308426 94054
rect 308662 93818 308746 94054
rect 308982 93818 344426 94054
rect 344662 93818 344746 94054
rect 344982 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 488426 94054
rect 488662 93818 488746 94054
rect 488982 93818 524426 94054
rect 524662 93818 524746 94054
rect 524982 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 592650 94054
rect -8726 93734 592650 93818
rect -8726 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 56426 93734
rect 56662 93498 56746 93734
rect 56982 93498 92426 93734
rect 92662 93498 92746 93734
rect 92982 93498 128426 93734
rect 128662 93498 128746 93734
rect 128982 93498 164426 93734
rect 164662 93498 164746 93734
rect 164982 93498 200426 93734
rect 200662 93498 200746 93734
rect 200982 93498 236426 93734
rect 236662 93498 236746 93734
rect 236982 93498 272426 93734
rect 272662 93498 272746 93734
rect 272982 93498 308426 93734
rect 308662 93498 308746 93734
rect 308982 93498 344426 93734
rect 344662 93498 344746 93734
rect 344982 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 488426 93734
rect 488662 93498 488746 93734
rect 488982 93498 524426 93734
rect 524662 93498 524746 93734
rect 524982 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 592650 93734
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 52706 90334
rect 52942 90098 53026 90334
rect 53262 90098 88706 90334
rect 88942 90098 89026 90334
rect 89262 90098 124706 90334
rect 124942 90098 125026 90334
rect 125262 90098 160706 90334
rect 160942 90098 161026 90334
rect 161262 90098 196706 90334
rect 196942 90098 197026 90334
rect 197262 90098 232706 90334
rect 232942 90098 233026 90334
rect 233262 90098 268706 90334
rect 268942 90098 269026 90334
rect 269262 90098 304706 90334
rect 304942 90098 305026 90334
rect 305262 90098 340706 90334
rect 340942 90098 341026 90334
rect 341262 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 412706 90334
rect 412942 90098 413026 90334
rect 413262 90098 448706 90334
rect 448942 90098 449026 90334
rect 449262 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 520706 90334
rect 520942 90098 521026 90334
rect 521262 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 592650 90334
rect -8726 90014 592650 90098
rect -8726 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 52706 90014
rect 52942 89778 53026 90014
rect 53262 89778 88706 90014
rect 88942 89778 89026 90014
rect 89262 89778 124706 90014
rect 124942 89778 125026 90014
rect 125262 89778 160706 90014
rect 160942 89778 161026 90014
rect 161262 89778 196706 90014
rect 196942 89778 197026 90014
rect 197262 89778 232706 90014
rect 232942 89778 233026 90014
rect 233262 89778 268706 90014
rect 268942 89778 269026 90014
rect 269262 89778 304706 90014
rect 304942 89778 305026 90014
rect 305262 89778 340706 90014
rect 340942 89778 341026 90014
rect 341262 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 412706 90014
rect 412942 89778 413026 90014
rect 413262 89778 448706 90014
rect 448942 89778 449026 90014
rect 449262 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 520706 90014
rect 520942 89778 521026 90014
rect 521262 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 592650 90014
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 592650 86294
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 592650 82894
rect -8726 82574 592650 82658
rect -8726 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 592650 82574
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 59174 79174
rect 59410 78938 67362 79174
rect 67598 78938 75550 79174
rect 75786 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 83738 79174
rect 83974 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 592650 79174
rect -8726 78854 592650 78938
rect -8726 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 59174 78854
rect 59410 78618 67362 78854
rect 67598 78618 75550 78854
rect 75786 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 83738 78854
rect 83974 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 592650 78854
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 55080 75454
rect 55316 75218 63268 75454
rect 63504 75218 71456 75454
rect 71692 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 79644 75454
rect 79880 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 55080 75134
rect 55316 74898 63268 75134
rect 63504 74898 71456 75134
rect 71692 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 79644 75134
rect 79880 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 63866 65494
rect 64102 65258 64186 65494
rect 64422 65258 99866 65494
rect 100102 65258 100186 65494
rect 100422 65258 135866 65494
rect 136102 65258 136186 65494
rect 136422 65258 171866 65494
rect 172102 65258 172186 65494
rect 172422 65258 207866 65494
rect 208102 65258 208186 65494
rect 208422 65258 243866 65494
rect 244102 65258 244186 65494
rect 244422 65258 279866 65494
rect 280102 65258 280186 65494
rect 280422 65258 315866 65494
rect 316102 65258 316186 65494
rect 316422 65258 351866 65494
rect 352102 65258 352186 65494
rect 352422 65258 387866 65494
rect 388102 65258 388186 65494
rect 388422 65258 423866 65494
rect 424102 65258 424186 65494
rect 424422 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect -8726 65174 592650 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 63866 65174
rect 64102 64938 64186 65174
rect 64422 64938 99866 65174
rect 100102 64938 100186 65174
rect 100422 64938 135866 65174
rect 136102 64938 136186 65174
rect 136422 64938 171866 65174
rect 172102 64938 172186 65174
rect 172422 64938 207866 65174
rect 208102 64938 208186 65174
rect 208422 64938 243866 65174
rect 244102 64938 244186 65174
rect 244422 64938 279866 65174
rect 280102 64938 280186 65174
rect 280422 64938 315866 65174
rect 316102 64938 316186 65174
rect 316422 64938 351866 65174
rect 352102 64938 352186 65174
rect 352422 64938 387866 65174
rect 388102 64938 388186 65174
rect 388422 64938 423866 65174
rect 424102 64938 424186 65174
rect 424422 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 24146 61774
rect 24382 61538 24466 61774
rect 24702 61538 60146 61774
rect 60382 61538 60466 61774
rect 60702 61538 96146 61774
rect 96382 61538 96466 61774
rect 96702 61538 132146 61774
rect 132382 61538 132466 61774
rect 132702 61538 168146 61774
rect 168382 61538 168466 61774
rect 168702 61538 204146 61774
rect 204382 61538 204466 61774
rect 204702 61538 240146 61774
rect 240382 61538 240466 61774
rect 240702 61538 276146 61774
rect 276382 61538 276466 61774
rect 276702 61538 312146 61774
rect 312382 61538 312466 61774
rect 312702 61538 348146 61774
rect 348382 61538 348466 61774
rect 348702 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 420146 61774
rect 420382 61538 420466 61774
rect 420702 61538 456146 61774
rect 456382 61538 456466 61774
rect 456702 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 592650 61774
rect -8726 61454 592650 61538
rect -8726 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 24146 61454
rect 24382 61218 24466 61454
rect 24702 61218 60146 61454
rect 60382 61218 60466 61454
rect 60702 61218 96146 61454
rect 96382 61218 96466 61454
rect 96702 61218 132146 61454
rect 132382 61218 132466 61454
rect 132702 61218 168146 61454
rect 168382 61218 168466 61454
rect 168702 61218 204146 61454
rect 204382 61218 204466 61454
rect 204702 61218 240146 61454
rect 240382 61218 240466 61454
rect 240702 61218 276146 61454
rect 276382 61218 276466 61454
rect 276702 61218 312146 61454
rect 312382 61218 312466 61454
rect 312702 61218 348146 61454
rect 348382 61218 348466 61454
rect 348702 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 420146 61454
rect 420382 61218 420466 61454
rect 420702 61218 456146 61454
rect 456382 61218 456466 61454
rect 456702 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 592650 61454
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 56426 58054
rect 56662 57818 56746 58054
rect 56982 57818 92426 58054
rect 92662 57818 92746 58054
rect 92982 57818 128426 58054
rect 128662 57818 128746 58054
rect 128982 57818 164426 58054
rect 164662 57818 164746 58054
rect 164982 57818 200426 58054
rect 200662 57818 200746 58054
rect 200982 57818 236426 58054
rect 236662 57818 236746 58054
rect 236982 57818 272426 58054
rect 272662 57818 272746 58054
rect 272982 57818 308426 58054
rect 308662 57818 308746 58054
rect 308982 57818 344426 58054
rect 344662 57818 344746 58054
rect 344982 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 416426 58054
rect 416662 57818 416746 58054
rect 416982 57818 452426 58054
rect 452662 57818 452746 58054
rect 452982 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 592650 58054
rect -8726 57734 592650 57818
rect -8726 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 56426 57734
rect 56662 57498 56746 57734
rect 56982 57498 92426 57734
rect 92662 57498 92746 57734
rect 92982 57498 128426 57734
rect 128662 57498 128746 57734
rect 128982 57498 164426 57734
rect 164662 57498 164746 57734
rect 164982 57498 200426 57734
rect 200662 57498 200746 57734
rect 200982 57498 236426 57734
rect 236662 57498 236746 57734
rect 236982 57498 272426 57734
rect 272662 57498 272746 57734
rect 272982 57498 308426 57734
rect 308662 57498 308746 57734
rect 308982 57498 344426 57734
rect 344662 57498 344746 57734
rect 344982 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 416426 57734
rect 416662 57498 416746 57734
rect 416982 57498 452426 57734
rect 452662 57498 452746 57734
rect 452982 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 592650 57734
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 52706 54334
rect 52942 54098 53026 54334
rect 53262 54098 88706 54334
rect 88942 54098 89026 54334
rect 89262 54098 124706 54334
rect 124942 54098 125026 54334
rect 125262 54098 160706 54334
rect 160942 54098 161026 54334
rect 161262 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 232706 54334
rect 232942 54098 233026 54334
rect 233262 54098 268706 54334
rect 268942 54098 269026 54334
rect 269262 54098 304706 54334
rect 304942 54098 305026 54334
rect 305262 54098 340706 54334
rect 340942 54098 341026 54334
rect 341262 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 412706 54334
rect 412942 54098 413026 54334
rect 413262 54098 448706 54334
rect 448942 54098 449026 54334
rect 449262 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 592650 54334
rect -8726 54014 592650 54098
rect -8726 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 52706 54014
rect 52942 53778 53026 54014
rect 53262 53778 88706 54014
rect 88942 53778 89026 54014
rect 89262 53778 124706 54014
rect 124942 53778 125026 54014
rect 125262 53778 160706 54014
rect 160942 53778 161026 54014
rect 161262 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 232706 54014
rect 232942 53778 233026 54014
rect 233262 53778 268706 54014
rect 268942 53778 269026 54014
rect 269262 53778 304706 54014
rect 304942 53778 305026 54014
rect 305262 53778 340706 54014
rect 340942 53778 341026 54014
rect 341262 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 412706 54014
rect 412942 53778 413026 54014
rect 413262 53778 448706 54014
rect 448942 53778 449026 54014
rect 449262 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 592650 54014
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 592650 50294
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 592650 46894
rect -8726 46574 592650 46658
rect -8726 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 592650 46574
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 592650 43174
rect -8726 42854 592650 42938
rect -8726 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 592650 42854
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect -8726 29174 592650 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 592650 25774
rect -8726 25454 592650 25538
rect -8726 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 592650 25454
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 592650 22054
rect -8726 21734 592650 21818
rect -8726 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 592650 21734
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 592650 18334
rect -8726 18014 592650 18098
rect -8726 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 592650 18014
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 592650 14294
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 592650 10894
rect -8726 10574 592650 10658
rect -8726 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 592650 10574
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 592650 7174
rect -8726 6854 592650 6938
rect -8726 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 592650 6854
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use ci2406_z80  ci2406_z80
timestamp 0
transform 1 0 50000 0 1 280000
box 0 0 60000 60000
use multiplexer  multiplexer
timestamp 0
transform 1 0 240000 0 1 240000
box 0 0 40000 200000
use scrapcpu  scrapcpu
timestamp 0
transform 1 0 490000 0 1 600000
box 0 0 50000 55000
use unused_tie  unused_tie
timestamp 0
transform 1 0 50000 0 1 50000
box 0 0 35000 35000
use vliw  vliw
timestamp 0
transform 1 0 70000 0 1 480000
box 0 0 220000 150000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 278167 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 340449 74414 478303 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 629612 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 278167 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 340449 110414 478303 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 629257 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 478303 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 629257 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 478303 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 629612 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 478303 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 629257 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 241295 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 402313 254414 478303 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 629257 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 600207 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 654737 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 -7654 45854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 -7654 81854 278167 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 340449 81854 478303 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 629257 81854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 -7654 117854 478303 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 629257 117854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 -7654 153854 478303 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 629257 153854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 -7654 189854 478303 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 629257 189854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 -7654 225854 478303 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 629257 225854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 -7654 261854 241295 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 402313 261854 478303 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 629257 261854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 -7654 297854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 -7654 333854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 -7654 369854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 -7654 405854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 -7654 441854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 -7654 477854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 -7654 513854 600207 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 654737 513854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 -7654 549854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 16674 -7654 17294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 52674 -7654 53294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 -7654 89294 278167 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 340449 89294 478303 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 629257 89294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 -7654 125294 478303 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 629257 125294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 160674 -7654 161294 478303 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 160674 629257 161294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 -7654 197294 478303 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 629612 197294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 -7654 233294 478303 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 629257 233294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 -7654 269294 241295 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 402313 269294 478303 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 629257 269294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 -7654 305294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 -7654 341294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 -7654 377294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 -7654 413294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 -7654 449294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 -7654 485294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 -7654 521294 600207 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 654737 521294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 -7654 557294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 24114 -7654 24734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 -7654 60734 278167 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 340449 60734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 -7654 96734 278167 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 340449 96734 478303 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 629257 96734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132114 -7654 132734 478303 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132114 629257 132734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168114 -7654 168734 478303 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168114 629257 168734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 -7654 204734 478303 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 629257 204734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 -7654 240734 241295 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 402313 240734 478303 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 629257 240734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 -7654 276734 241295 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 402313 276734 478303 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 629257 276734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 -7654 312734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 -7654 348734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 -7654 384734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 -7654 420734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 -7654 456734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 -7654 492734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 -7654 528734 600207 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 654737 528734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 -7654 564734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 20394 -7654 21014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 56394 -7654 57014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 -7654 93014 278167 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 340449 93014 478303 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 629257 93014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 -7654 129014 478303 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 629257 129014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 -7654 165014 478303 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 629257 165014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 -7654 201014 478303 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 629257 201014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 -7654 237014 478303 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 629257 237014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 -7654 273014 241295 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 402313 273014 478303 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 629257 273014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 -7654 309014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 -7654 345014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380394 -7654 381014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 -7654 417014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 -7654 453014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 -7654 489014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 -7654 525014 599988 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 654956 525014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 -7654 561014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 27834 -7654 28454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 -7654 64454 278167 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 340449 64454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 -7654 100454 278167 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 340449 100454 478303 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 629257 100454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 -7654 136454 478303 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 629612 136454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 -7654 172454 478303 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 629257 172454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 -7654 208454 478303 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 629257 208454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 -7654 244454 239988 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 629257 244454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 -7654 280454 478303 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 629257 280454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 -7654 316454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 -7654 352454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 -7654 388454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 -7654 424454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 -7654 460454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 -7654 496454 600207 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 654737 496454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 -7654 532454 600207 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 654737 532454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 567834 -7654 568454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 -7654 42134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 -7654 78134 278167 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 340449 78134 478303 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 629257 78134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 -7654 114134 478303 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 629257 114134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 -7654 150134 478303 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 629257 150134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 -7654 186134 478303 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 629257 186134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 -7654 222134 478303 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 629257 222134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 -7654 258134 241295 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 402313 258134 478303 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 629257 258134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 -7654 294134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 -7654 330134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 -7654 366134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 -7654 402134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 -7654 438134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 -7654 474134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 -7654 510134 599988 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 654956 510134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 -7654 546134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 12954 -7654 13574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 -7654 49574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 -7654 85574 278167 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 340449 85574 478303 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 629257 85574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 -7654 121574 478303 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 629257 121574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 -7654 157574 478303 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 629257 157574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 -7654 193574 478303 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 629257 193574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 -7654 229574 478303 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 629257 229574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 -7654 265574 241295 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 402313 265574 478303 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 629257 265574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 -7654 301574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 -7654 337574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 -7654 373574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 -7654 409574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 -7654 445574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 -7654 481574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 -7654 517574 600207 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 654737 517574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 -7654 553574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
