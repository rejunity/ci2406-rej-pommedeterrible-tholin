// This is the unpowered netlist.
module unused_tie (wb_clk_i,
    wb_rst_i,
    irq,
    la_data_out);
 input wb_clk_i;
 input wb_rst_i;
 output [2:0] irq;
 output [87:0] la_data_out;

 wire net97;
 wire net98;
 wire net99;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0__leaf_wb_clk_i;
 wire clknet_3_1__leaf_wb_clk_i;
 wire clknet_3_2__leaf_wb_clk_i;
 wire clknet_3_3__leaf_wb_clk_i;
 wire clknet_3_4__leaf_wb_clk_i;
 wire clknet_3_5__leaf_wb_clk_i;
 wire clknet_3_6__leaf_wb_clk_i;
 wire clknet_3_7__leaf_wb_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;

 sky130_fd_sc_hd__diode_2 ANTENNA__088__A_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__089__A_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__090__A_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__091__A_N (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__092__A_N (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__093__A_N (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__094__A_N (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__095__A_N (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__096__A_N (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__097__A_N (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__098__A_N (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__099__A_N (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__100__A_N (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__101__A_N (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__102__A_N (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__103__A_N (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__104__A_N (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__105__A_N (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__106__A_N (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__107__A_N (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__108__A_N (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__109__A_N (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__110__A_N (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__111__A_N (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__112__A_N (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__113__A_N (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__114__A_N (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__115__A_N (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__116__A_N (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__117__A_N (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__118__A_N (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__119__A_N (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__120__A_N (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__121__A_N (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__122__A_N (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__123__A_N (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__124__A_N (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__125__A_N (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__126__A_N (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__127__A_N (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__128__A_N (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__129__A_N (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__130__A_N (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__131__A_N (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__131__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__132__A_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__133__A_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__134__A_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__135__A_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__136__A_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__137__A_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__138__A_N (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__139__A_N (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__140__A_N (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__141__A_N (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__151__A_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__152__A_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__153__A_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__154__A_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__155__A_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__156__A_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__157__A_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__158__A_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__161__A_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__162__A_N (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__163__A_N (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__164__A_N (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__165__A_N (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__166__A_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__167__A_N (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__173__A_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__174__A_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__175__A_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__179__CLK (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__180__CLK (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__181__CLK (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__182__CLK (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__183__CLK (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__184__CLK (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__185__CLK (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__189__CLK (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__190__CLK (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__191__CLK (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__192__CLK (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__193__CLK (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__194__CLK (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__195__CLK (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__219__CLK (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__250__CLK (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__251__CLK (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__252__CLK (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout91_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout93_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout94_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout95_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold330_A (.DIODE(net250));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_97 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__and2b_1 _088_ (.A_N(net92),
    .B(net124),
    .X(_000_));
 sky130_fd_sc_hd__and2b_1 _089_ (.A_N(net92),
    .B(net114),
    .X(_001_));
 sky130_fd_sc_hd__and2b_1 _090_ (.A_N(net92),
    .B(net118),
    .X(_002_));
 sky130_fd_sc_hd__and2b_1 _091_ (.A_N(net94),
    .B(net176),
    .X(_003_));
 sky130_fd_sc_hd__and2b_1 _092_ (.A_N(net94),
    .B(net186),
    .X(_004_));
 sky130_fd_sc_hd__and2b_1 _093_ (.A_N(net94),
    .B(net202),
    .X(_005_));
 sky130_fd_sc_hd__and2b_1 _094_ (.A_N(net94),
    .B(net134),
    .X(_006_));
 sky130_fd_sc_hd__and2b_1 _095_ (.A_N(net94),
    .B(net150),
    .X(_007_));
 sky130_fd_sc_hd__and2b_1 _096_ (.A_N(net94),
    .B(net198),
    .X(_008_));
 sky130_fd_sc_hd__and2b_1 _097_ (.A_N(net94),
    .B(net212),
    .X(_009_));
 sky130_fd_sc_hd__and2b_1 _098_ (.A_N(net94),
    .B(net214),
    .X(_010_));
 sky130_fd_sc_hd__and2b_1 _099_ (.A_N(net94),
    .B(net222),
    .X(_011_));
 sky130_fd_sc_hd__and2b_1 _100_ (.A_N(net94),
    .B(net268),
    .X(_012_));
 sky130_fd_sc_hd__and2b_1 _101_ (.A_N(net93),
    .B(net256),
    .X(_013_));
 sky130_fd_sc_hd__and2b_1 _102_ (.A_N(net93),
    .B(net126),
    .X(_014_));
 sky130_fd_sc_hd__and2b_1 _103_ (.A_N(net93),
    .B(net204),
    .X(_015_));
 sky130_fd_sc_hd__and2b_1 _104_ (.A_N(net93),
    .B(net130),
    .X(_016_));
 sky130_fd_sc_hd__and2b_1 _105_ (.A_N(net93),
    .B(net170),
    .X(_017_));
 sky130_fd_sc_hd__and2b_1 _106_ (.A_N(net93),
    .B(net192),
    .X(_018_));
 sky130_fd_sc_hd__and2b_1 _107_ (.A_N(net93),
    .B(net234),
    .X(_019_));
 sky130_fd_sc_hd__and2b_1 _108_ (.A_N(net93),
    .B(net210),
    .X(_020_));
 sky130_fd_sc_hd__and2b_1 _109_ (.A_N(net93),
    .B(net200),
    .X(_021_));
 sky130_fd_sc_hd__and2b_1 _110_ (.A_N(net93),
    .B(net208),
    .X(_022_));
 sky130_fd_sc_hd__and2b_1 _111_ (.A_N(net93),
    .B(net206),
    .X(_023_));
 sky130_fd_sc_hd__and2b_1 _112_ (.A_N(net93),
    .B(net184),
    .X(_024_));
 sky130_fd_sc_hd__and2b_1 _113_ (.A_N(net93),
    .B(net174),
    .X(_025_));
 sky130_fd_sc_hd__and2b_1 _114_ (.A_N(net95),
    .B(net178),
    .X(_026_));
 sky130_fd_sc_hd__and2b_1 _115_ (.A_N(net95),
    .B(net182),
    .X(_027_));
 sky130_fd_sc_hd__and2b_1 _116_ (.A_N(net95),
    .B(net188),
    .X(_028_));
 sky130_fd_sc_hd__and2b_1 _117_ (.A_N(net95),
    .B(net190),
    .X(_029_));
 sky130_fd_sc_hd__and2b_1 _118_ (.A_N(net95),
    .B(net194),
    .X(_030_));
 sky130_fd_sc_hd__and2b_1 _119_ (.A_N(net95),
    .B(net146),
    .X(_031_));
 sky130_fd_sc_hd__and2b_1 _120_ (.A_N(net94),
    .B(net144),
    .X(_032_));
 sky130_fd_sc_hd__and2b_1 _121_ (.A_N(net94),
    .B(net196),
    .X(_033_));
 sky130_fd_sc_hd__and2b_1 _122_ (.A_N(net94),
    .B(net164),
    .X(_034_));
 sky130_fd_sc_hd__and2b_1 _123_ (.A_N(net94),
    .B(net158),
    .X(_035_));
 sky130_fd_sc_hd__and2b_1 _124_ (.A_N(net94),
    .B(net154),
    .X(_036_));
 sky130_fd_sc_hd__and2b_1 _125_ (.A_N(net95),
    .B(net166),
    .X(_037_));
 sky130_fd_sc_hd__and2b_1 _126_ (.A_N(net95),
    .B(net168),
    .X(_038_));
 sky130_fd_sc_hd__and2b_1 _127_ (.A_N(net95),
    .B(net172),
    .X(_039_));
 sky130_fd_sc_hd__and2b_1 _128_ (.A_N(net95),
    .B(net162),
    .X(_040_));
 sky130_fd_sc_hd__and2b_1 _129_ (.A_N(net95),
    .B(net152),
    .X(_041_));
 sky130_fd_sc_hd__and2b_1 _130_ (.A_N(net95),
    .B(net248),
    .X(_042_));
 sky130_fd_sc_hd__and2b_1 _131_ (.A_N(net93),
    .B(net250),
    .X(_043_));
 sky130_fd_sc_hd__and2b_1 _132_ (.A_N(net90),
    .B(net160),
    .X(_044_));
 sky130_fd_sc_hd__and2b_1 _133_ (.A_N(net90),
    .B(net156),
    .X(_045_));
 sky130_fd_sc_hd__and2b_1 _134_ (.A_N(net90),
    .B(net140),
    .X(_046_));
 sky130_fd_sc_hd__and2b_1 _135_ (.A_N(net90),
    .B(net142),
    .X(_047_));
 sky130_fd_sc_hd__and2b_1 _136_ (.A_N(net90),
    .B(net138),
    .X(_048_));
 sky130_fd_sc_hd__and2b_1 _137_ (.A_N(net90),
    .B(net148),
    .X(_049_));
 sky130_fd_sc_hd__and2b_1 _138_ (.A_N(net96),
    .B(net136),
    .X(_050_));
 sky130_fd_sc_hd__and2b_1 _139_ (.A_N(net96),
    .B(net180),
    .X(_051_));
 sky130_fd_sc_hd__and2b_1 _140_ (.A_N(net96),
    .B(net262),
    .X(_052_));
 sky130_fd_sc_hd__and2b_1 _141_ (.A_N(net96),
    .B(net258),
    .X(_053_));
 sky130_fd_sc_hd__and2b_1 _142_ (.A_N(net91),
    .B(net238),
    .X(_054_));
 sky130_fd_sc_hd__and2b_1 _143_ (.A_N(net91),
    .B(net224),
    .X(_055_));
 sky130_fd_sc_hd__and2b_1 _144_ (.A_N(net91),
    .B(net220),
    .X(_056_));
 sky130_fd_sc_hd__and2b_1 _145_ (.A_N(net91),
    .B(net216),
    .X(_057_));
 sky130_fd_sc_hd__and2b_1 _146_ (.A_N(net91),
    .B(net226),
    .X(_058_));
 sky130_fd_sc_hd__and2b_1 _147_ (.A_N(net91),
    .B(net218),
    .X(_059_));
 sky130_fd_sc_hd__and2b_1 _148_ (.A_N(net91),
    .B(net230),
    .X(_060_));
 sky130_fd_sc_hd__and2b_1 _149_ (.A_N(net91),
    .B(net232),
    .X(_061_));
 sky130_fd_sc_hd__and2b_1 _150_ (.A_N(net91),
    .B(net266),
    .X(_062_));
 sky130_fd_sc_hd__and2b_1 _151_ (.A_N(net90),
    .B(net240),
    .X(_063_));
 sky130_fd_sc_hd__and2b_1 _152_ (.A_N(net90),
    .B(net110),
    .X(_064_));
 sky130_fd_sc_hd__and2b_1 _153_ (.A_N(net90),
    .B(net108),
    .X(_065_));
 sky130_fd_sc_hd__and2b_1 _154_ (.A_N(net90),
    .B(net104),
    .X(_066_));
 sky130_fd_sc_hd__and2b_1 _155_ (.A_N(net90),
    .B(net100),
    .X(_067_));
 sky130_fd_sc_hd__and2b_1 _156_ (.A_N(net90),
    .B(net106),
    .X(_068_));
 sky130_fd_sc_hd__and2b_1 _157_ (.A_N(net90),
    .B(net102),
    .X(_069_));
 sky130_fd_sc_hd__and2b_1 _158_ (.A_N(net90),
    .B(net242),
    .X(_070_));
 sky130_fd_sc_hd__and2b_1 _159_ (.A_N(net91),
    .B(net270),
    .X(_071_));
 sky130_fd_sc_hd__or2_1 _160_ (.A(net91),
    .B(net264),
    .X(_072_));
 sky130_fd_sc_hd__and2b_1 _161_ (.A_N(net92),
    .B(net260),
    .X(_073_));
 sky130_fd_sc_hd__and2b_1 _162_ (.A_N(net94),
    .B(net272),
    .X(_074_));
 sky130_fd_sc_hd__and2b_1 _163_ (.A_N(net93),
    .B(net246),
    .X(_075_));
 sky130_fd_sc_hd__and2b_1 _164_ (.A_N(net93),
    .B(net244),
    .X(_076_));
 sky130_fd_sc_hd__and2b_1 _165_ (.A_N(net96),
    .B(net254),
    .X(_077_));
 sky130_fd_sc_hd__and2b_1 _166_ (.A_N(net90),
    .B(net228),
    .X(_078_));
 sky130_fd_sc_hd__and2b_1 _167_ (.A_N(net90),
    .B(net274),
    .X(_079_));
 sky130_fd_sc_hd__and2b_1 _168_ (.A_N(net91),
    .B(net252),
    .X(_080_));
 sky130_fd_sc_hd__and2b_1 _169_ (.A_N(net91),
    .B(net236),
    .X(_081_));
 sky130_fd_sc_hd__and2b_1 _170_ (.A_N(net91),
    .B(net116),
    .X(_082_));
 sky130_fd_sc_hd__and2b_1 _171_ (.A_N(net91),
    .B(net128),
    .X(_083_));
 sky130_fd_sc_hd__and2b_1 _172_ (.A_N(net91),
    .B(net122),
    .X(_084_));
 sky130_fd_sc_hd__and2b_1 _173_ (.A_N(net92),
    .B(net120),
    .X(_085_));
 sky130_fd_sc_hd__and2b_1 _174_ (.A_N(net92),
    .B(net112),
    .X(_086_));
 sky130_fd_sc_hd__and2b_1 _175_ (.A_N(net92),
    .B(net132),
    .X(_087_));
 sky130_fd_sc_hd__dfxtp_1 _176_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_000_),
    .Q(net9));
 sky130_fd_sc_hd__dfxtp_1 _177_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_001_),
    .Q(net10));
 sky130_fd_sc_hd__dfxtp_1 _178_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_002_),
    .Q(net11));
 sky130_fd_sc_hd__dfxtp_1 _179_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_003_),
    .Q(net12));
 sky130_fd_sc_hd__dfxtp_1 _180_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_004_),
    .Q(net14));
 sky130_fd_sc_hd__dfxtp_1 _181_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_005_),
    .Q(net15));
 sky130_fd_sc_hd__dfxtp_1 _182_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_006_),
    .Q(net16));
 sky130_fd_sc_hd__dfxtp_1 _183_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_007_),
    .Q(net17));
 sky130_fd_sc_hd__dfxtp_1 _184_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_008_),
    .Q(net18));
 sky130_fd_sc_hd__dfxtp_1 _185_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_009_),
    .Q(net19));
 sky130_fd_sc_hd__dfxtp_1 _186_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_010_),
    .Q(net20));
 sky130_fd_sc_hd__dfxtp_1 _187_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_011_),
    .Q(net21));
 sky130_fd_sc_hd__dfxtp_1 _188_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_012_),
    .Q(net22));
 sky130_fd_sc_hd__dfxtp_1 _189_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_013_),
    .Q(net23));
 sky130_fd_sc_hd__dfxtp_1 _190_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_014_),
    .Q(net25));
 sky130_fd_sc_hd__dfxtp_1 _191_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_015_),
    .Q(net26));
 sky130_fd_sc_hd__dfxtp_1 _192_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_016_),
    .Q(net27));
 sky130_fd_sc_hd__dfxtp_1 _193_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_017_),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_1 _194_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_018_),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_1 _195_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_019_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_1 _196_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_020_),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_1 _197_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_021_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_1 _198_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_022_),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_1 _199_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_023_),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_1 _200_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_024_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_1 _201_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_025_),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_1 _202_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_026_),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_1 _203_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_027_),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_1 _204_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_028_),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_1 _205_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_029_),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_1 _206_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_030_),
    .Q(net42));
 sky130_fd_sc_hd__dfxtp_1 _207_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_031_),
    .Q(net43));
 sky130_fd_sc_hd__dfxtp_1 _208_ (.CLK(clknet_3_5__leaf_wb_clk_i),
    .D(_032_),
    .Q(net44));
 sky130_fd_sc_hd__dfxtp_1 _209_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_033_),
    .Q(net45));
 sky130_fd_sc_hd__dfxtp_1 _210_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_034_),
    .Q(net47));
 sky130_fd_sc_hd__dfxtp_1 _211_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_035_),
    .Q(net48));
 sky130_fd_sc_hd__dfxtp_1 _212_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_036_),
    .Q(net49));
 sky130_fd_sc_hd__dfxtp_1 _213_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_037_),
    .Q(net50));
 sky130_fd_sc_hd__dfxtp_1 _214_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_038_),
    .Q(net51));
 sky130_fd_sc_hd__dfxtp_1 _215_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_039_),
    .Q(net52));
 sky130_fd_sc_hd__dfxtp_1 _216_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_040_),
    .Q(net53));
 sky130_fd_sc_hd__dfxtp_1 _217_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_041_),
    .Q(net54));
 sky130_fd_sc_hd__dfxtp_1 _218_ (.CLK(clknet_3_7__leaf_wb_clk_i),
    .D(_042_),
    .Q(net55));
 sky130_fd_sc_hd__dfxtp_1 _219_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_043_),
    .Q(net56));
 sky130_fd_sc_hd__dfxtp_1 _220_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_044_),
    .Q(net58));
 sky130_fd_sc_hd__dfxtp_1 _221_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_045_),
    .Q(net59));
 sky130_fd_sc_hd__dfxtp_1 _222_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_046_),
    .Q(net60));
 sky130_fd_sc_hd__dfxtp_1 _223_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_047_),
    .Q(net61));
 sky130_fd_sc_hd__dfxtp_1 _224_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_048_),
    .Q(net62));
 sky130_fd_sc_hd__dfxtp_1 _225_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_049_),
    .Q(net63));
 sky130_fd_sc_hd__dfxtp_1 _226_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_050_),
    .Q(net64));
 sky130_fd_sc_hd__dfxtp_1 _227_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_051_),
    .Q(net65));
 sky130_fd_sc_hd__dfxtp_1 _228_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_052_),
    .Q(net66));
 sky130_fd_sc_hd__dfxtp_1 _229_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_053_),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_1 _230_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_054_),
    .Q(net69));
 sky130_fd_sc_hd__dfxtp_1 _231_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_055_),
    .Q(net70));
 sky130_fd_sc_hd__dfxtp_1 _232_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_056_),
    .Q(net71));
 sky130_fd_sc_hd__dfxtp_1 _233_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_057_),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_1 _234_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_058_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_1 _235_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_059_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_1 _236_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_060_),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_1 _237_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_061_),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_1 _238_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_062_),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_1 _239_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_063_),
    .Q(net78));
 sky130_fd_sc_hd__dfxtp_1 _240_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_064_),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_1 _241_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_065_),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_1 _242_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_066_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_1 _243_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_067_),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_1 _244_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_068_),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_1 _245_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_069_),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_1 _246_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_070_),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_1 _247_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_071_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_1 _248_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_072_),
    .Q(net2));
 sky130_fd_sc_hd__dfxtp_1 _249_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_073_),
    .Q(net13));
 sky130_fd_sc_hd__dfxtp_1 _250_ (.CLK(clknet_3_6__leaf_wb_clk_i),
    .D(_074_),
    .Q(net24));
 sky130_fd_sc_hd__dfxtp_1 _251_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_075_),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_1 _252_ (.CLK(clknet_3_4__leaf_wb_clk_i),
    .D(_076_),
    .Q(net46));
 sky130_fd_sc_hd__dfxtp_1 _253_ (.CLK(clknet_3_1__leaf_wb_clk_i),
    .D(_077_),
    .Q(net57));
 sky130_fd_sc_hd__dfxtp_1 _254_ (.CLK(clknet_3_0__leaf_wb_clk_i),
    .D(_078_),
    .Q(net68));
 sky130_fd_sc_hd__dfxtp_1 _255_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_079_),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_1 _256_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_080_),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_1 _257_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_081_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_1 _258_ (.CLK(clknet_3_2__leaf_wb_clk_i),
    .D(_082_),
    .Q(net3));
 sky130_fd_sc_hd__dfxtp_1 _259_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_083_),
    .Q(net4));
 sky130_fd_sc_hd__dfxtp_1 _260_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_084_),
    .Q(net5));
 sky130_fd_sc_hd__dfxtp_1 _261_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_085_),
    .Q(net6));
 sky130_fd_sc_hd__dfxtp_1 _262_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_086_),
    .Q(net7));
 sky130_fd_sc_hd__dfxtp_1 _263_ (.CLK(clknet_3_3__leaf_wb_clk_i),
    .D(_087_),
    .Q(net8));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_4 fanout90 (.A(net96),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_4 fanout91 (.A(net92),
    .X(net91));
 sky130_fd_sc_hd__buf_2 fanout92 (.A(net96),
    .X(net92));
 sky130_fd_sc_hd__buf_4 fanout93 (.A(net95),
    .X(net93));
 sky130_fd_sc_hd__buf_4 fanout94 (.A(net95),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_4 fanout95 (.A(net96),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_4 fanout96 (.A(net1),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net302),
    .X(net100));
 sky130_fd_sc_hd__buf_12 hold10 (.A(net109),
    .X(la_data_out[82]));
 sky130_fd_sc_hd__buf_12 hold100 (.A(net199),
    .X(la_data_out[25]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(net346),
    .X(net200));
 sky130_fd_sc_hd__buf_12 hold102 (.A(net201),
    .X(la_data_out[38]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(net406),
    .X(net202));
 sky130_fd_sc_hd__buf_12 hold104 (.A(net203),
    .X(la_data_out[22]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(net420),
    .X(net204));
 sky130_fd_sc_hd__buf_12 hold106 (.A(net205),
    .X(la_data_out[32]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(net410),
    .X(net206));
 sky130_fd_sc_hd__buf_12 hold108 (.A(net207),
    .X(la_data_out[40]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(net364),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net380),
    .X(net110));
 sky130_fd_sc_hd__buf_12 hold110 (.A(net209),
    .X(la_data_out[39]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(net376),
    .X(net210));
 sky130_fd_sc_hd__buf_12 hold112 (.A(net211),
    .X(la_data_out[37]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(net284),
    .X(net212));
 sky130_fd_sc_hd__buf_12 hold114 (.A(net213),
    .X(la_data_out[26]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(net412),
    .X(net214));
 sky130_fd_sc_hd__buf_12 hold116 (.A(net215),
    .X(la_data_out[27]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(net370),
    .X(net216));
 sky130_fd_sc_hd__buf_12 hold118 (.A(net217),
    .X(la_data_out[74]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(net386),
    .X(net218));
 sky130_fd_sc_hd__buf_12 hold12 (.A(net111),
    .X(la_data_out[81]));
 sky130_fd_sc_hd__buf_12 hold120 (.A(net219),
    .X(la_data_out[76]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(net362),
    .X(net220));
 sky130_fd_sc_hd__buf_12 hold122 (.A(net221),
    .X(la_data_out[73]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(net416),
    .X(net222));
 sky130_fd_sc_hd__buf_12 hold124 (.A(net223),
    .X(la_data_out[28]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(net360),
    .X(net224));
 sky130_fd_sc_hd__buf_12 hold126 (.A(net225),
    .X(la_data_out[72]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(net378),
    .X(net226));
 sky130_fd_sc_hd__buf_12 hold128 (.A(net227),
    .X(la_data_out[75]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(net374),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net290),
    .X(net112));
 sky130_fd_sc_hd__buf_12 hold130 (.A(net229),
    .X(la_data_out[7]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(net382),
    .X(net230));
 sky130_fd_sc_hd__buf_12 hold132 (.A(net231),
    .X(la_data_out[77]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(net398),
    .X(net232));
 sky130_fd_sc_hd__buf_12 hold134 (.A(net233),
    .X(la_data_out[78]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(net292),
    .X(net234));
 sky130_fd_sc_hd__buf_12 hold136 (.A(net235),
    .X(la_data_out[36]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(net394),
    .X(net236));
 sky130_fd_sc_hd__buf_12 hold138 (.A(net237),
    .X(la_data_out[10]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(net400),
    .X(net238));
 sky130_fd_sc_hd__buf_12 hold14 (.A(net113),
    .X(la_data_out[15]));
 sky130_fd_sc_hd__buf_12 hold140 (.A(net239),
    .X(la_data_out[71]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(net422),
    .X(net240));
 sky130_fd_sc_hd__buf_12 hold142 (.A(net241),
    .X(la_data_out[80]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(net426),
    .X(net242));
 sky130_fd_sc_hd__buf_12 hold144 (.A(net243),
    .X(la_data_out[87]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(net282),
    .X(net244));
 sky130_fd_sc_hd__buf_12 hold146 (.A(net245),
    .X(la_data_out[5]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(net418),
    .X(net246));
 sky130_fd_sc_hd__buf_12 hold148 (.A(net247),
    .X(la_data_out[4]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(net286),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net288),
    .X(net114));
 sky130_fd_sc_hd__buf_12 hold150 (.A(net249),
    .X(la_data_out[59]));
 sky130_fd_sc_hd__buf_1 hold151 (.A(net428),
    .X(net250));
 sky130_fd_sc_hd__buf_12 hold152 (.A(net251),
    .X(la_data_out[60]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(net434),
    .X(net252));
 sky130_fd_sc_hd__buf_12 hold154 (.A(net253),
    .X(la_data_out[9]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(net432),
    .X(net254));
 sky130_fd_sc_hd__buf_12 hold156 (.A(net255),
    .X(la_data_out[6]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(net444),
    .X(net256));
 sky130_fd_sc_hd__buf_12 hold158 (.A(net257),
    .X(la_data_out[30]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(net438),
    .X(net258));
 sky130_fd_sc_hd__buf_12 hold16 (.A(net115),
    .X(la_data_out[18]));
 sky130_fd_sc_hd__buf_12 hold160 (.A(net259),
    .X(la_data_out[70]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(net436),
    .X(net260));
 sky130_fd_sc_hd__buf_12 hold162 (.A(net261),
    .X(la_data_out[2]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(net446),
    .X(net262));
 sky130_fd_sc_hd__buf_12 hold164 (.A(net263),
    .X(la_data_out[69]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(net424),
    .X(net264));
 sky130_fd_sc_hd__buf_12 hold166 (.A(net265),
    .X(la_data_out[1]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(net440),
    .X(net266));
 sky130_fd_sc_hd__buf_12 hold168 (.A(net267),
    .X(la_data_out[79]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(net430),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net276),
    .X(net116));
 sky130_fd_sc_hd__buf_12 hold170 (.A(net269),
    .X(la_data_out[29]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(net448),
    .X(net270));
 sky130_fd_sc_hd__buf_12 hold172 (.A(net271),
    .X(la_data_out[0]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(net442),
    .X(net272));
 sky130_fd_sc_hd__buf_12 hold174 (.A(net273),
    .X(la_data_out[3]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(net450),
    .X(net274));
 sky130_fd_sc_hd__buf_12 hold176 (.A(net275),
    .X(la_data_out[8]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(net4),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(net116),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(net12),
    .X(net278));
 sky130_fd_sc_hd__buf_12 hold18 (.A(net117),
    .X(la_data_out[11]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(net118),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(net45),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(net144),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(net57),
    .X(net282));
 sky130_fd_sc_hd__buf_1 hold184 (.A(net244),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(net20),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(net212),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(net56),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(net248),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(net11),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net278),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(net114),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(net8),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(net112),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(net31),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(net234),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(net44),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(net146),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(net55),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(net152),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(net83),
    .X(net298));
 sky130_fd_sc_hd__buf_12 hold2 (.A(net101),
    .X(la_data_out[84]));
 sky130_fd_sc_hd__buf_12 hold20 (.A(net119),
    .X(la_data_out[19]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(net104),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(net86),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(net102),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(net84),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(net100),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(net26),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(net126),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(net7),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(net120),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(net85),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net306),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(net106),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(net62),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(net142),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(net10),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(net124),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(net82),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(net108),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(net65),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(net136),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(net28),
    .X(net318));
 sky130_fd_sc_hd__buf_12 hold22 (.A(net121),
    .X(la_data_out[14]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(net130),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(net54),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(net162),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(net50),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(net154),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(net5),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(net128),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(net48),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(net164),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(net37),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net342),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(net184),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(net52),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(net168),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(net43),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(net194),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(net39),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(net178),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(net41),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(net188),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(net53),
    .X(net338));
 sky130_fd_sc_hd__buf_12 hold24 (.A(net123),
    .X(la_data_out[13]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(net172),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(net49),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(net158),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(net6),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(net122),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(net38),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(net174),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(net33),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(net200),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(net63),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net312),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(net138),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(net42),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(net190),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(net51),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(net166),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(net40),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(net182),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(net60),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(net156),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(net17),
    .X(net358));
 sky130_fd_sc_hd__buf_12 hold26 (.A(net125),
    .X(la_data_out[17]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(net134),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(net71),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(net224),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(net72),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(net220),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(net34),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(net208),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(net64),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(net148),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(net9),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net304),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(net132),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(net73),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(net216),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(net66),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(net180),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(net79),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(net228),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(net32),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(net210),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(net74),
    .X(net378));
 sky130_fd_sc_hd__buf_12 hold28 (.A(net127),
    .X(la_data_out[31]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(net226),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(net81),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(net110),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(net76),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(net230),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(net59),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(net160),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(net75),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(net218),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(net47),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net324),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(net196),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(net61),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(net140),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(net18),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(net150),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(net3),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(net236),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(net15),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(net186),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(net77),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net300),
    .X(net102));
 sky130_fd_sc_hd__buf_12 hold30 (.A(net129),
    .X(la_data_out[12]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(net232),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(net70),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(net238),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(net14),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(net176),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(net30),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(net192),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(net16),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(net202),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(net19),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(net318),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(net198),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(net36),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(net206),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(net21),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(net214),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(net29),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(net170),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(net22),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(net222),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(net46),
    .X(net418));
 sky130_fd_sc_hd__buf_12 hold32 (.A(net131),
    .X(la_data_out[33]));
 sky130_fd_sc_hd__buf_1 hold320 (.A(net246),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(net27),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(net204),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(net80),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(net240),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(net13),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(net264),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(net87),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(net242),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(net452),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net368),
    .X(net132));
 sky130_fd_sc_hd__buf_1 hold330 (.A(net250),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(net23),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(net268),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(net68),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(net254),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(net89),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(net252),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(net24),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(net260),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(net69),
    .X(net438));
 sky130_fd_sc_hd__buf_12 hold34 (.A(net133),
    .X(la_data_out[16]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(net258),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(net78),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(net266),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(net35),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(net272),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(net25),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(net256),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(net67),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(net262),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(net2),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net358),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(net270),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(net88),
    .X(net450));
 sky130_fd_sc_hd__buf_1 hold352 (.A(net274),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(net58),
    .X(net452));
 sky130_fd_sc_hd__buf_12 hold36 (.A(net135),
    .X(la_data_out[23]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net316),
    .X(net136));
 sky130_fd_sc_hd__buf_12 hold38 (.A(net137),
    .X(la_data_out[67]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(net348),
    .X(net138));
 sky130_fd_sc_hd__buf_12 hold4 (.A(net103),
    .X(la_data_out[86]));
 sky130_fd_sc_hd__buf_12 hold40 (.A(net139),
    .X(la_data_out[65]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net390),
    .X(net140));
 sky130_fd_sc_hd__buf_12 hold42 (.A(net141),
    .X(la_data_out[63]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net310),
    .X(net142));
 sky130_fd_sc_hd__buf_12 hold44 (.A(net143),
    .X(la_data_out[64]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net280),
    .X(net144));
 sky130_fd_sc_hd__buf_12 hold46 (.A(net145),
    .X(la_data_out[49]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net294),
    .X(net146));
 sky130_fd_sc_hd__buf_12 hold48 (.A(net147),
    .X(la_data_out[48]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net366),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net298),
    .X(net104));
 sky130_fd_sc_hd__buf_12 hold50 (.A(net149),
    .X(la_data_out[66]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(net392),
    .X(net150));
 sky130_fd_sc_hd__buf_12 hold52 (.A(net151),
    .X(la_data_out[24]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net296),
    .X(net152));
 sky130_fd_sc_hd__buf_12 hold54 (.A(net153),
    .X(la_data_out[58]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net322),
    .X(net154));
 sky130_fd_sc_hd__buf_12 hold56 (.A(net155),
    .X(la_data_out[53]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net356),
    .X(net156));
 sky130_fd_sc_hd__buf_12 hold58 (.A(net157),
    .X(la_data_out[62]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net340),
    .X(net158));
 sky130_fd_sc_hd__buf_12 hold6 (.A(net105),
    .X(la_data_out[83]));
 sky130_fd_sc_hd__buf_12 hold60 (.A(net159),
    .X(la_data_out[52]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net384),
    .X(net160));
 sky130_fd_sc_hd__buf_12 hold62 (.A(net161),
    .X(la_data_out[61]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net320),
    .X(net162));
 sky130_fd_sc_hd__buf_12 hold64 (.A(net163),
    .X(la_data_out[57]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net326),
    .X(net164));
 sky130_fd_sc_hd__buf_12 hold66 (.A(net165),
    .X(la_data_out[51]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net352),
    .X(net166));
 sky130_fd_sc_hd__buf_12 hold68 (.A(net167),
    .X(la_data_out[54]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(net330),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net308),
    .X(net106));
 sky130_fd_sc_hd__buf_12 hold70 (.A(net169),
    .X(la_data_out[55]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net414),
    .X(net170));
 sky130_fd_sc_hd__buf_12 hold72 (.A(net171),
    .X(la_data_out[34]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net338),
    .X(net172));
 sky130_fd_sc_hd__buf_12 hold74 (.A(net173),
    .X(la_data_out[56]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net344),
    .X(net174));
 sky130_fd_sc_hd__buf_12 hold76 (.A(net175),
    .X(la_data_out[42]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net402),
    .X(net176));
 sky130_fd_sc_hd__buf_12 hold78 (.A(net177),
    .X(la_data_out[20]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net334),
    .X(net178));
 sky130_fd_sc_hd__buf_12 hold8 (.A(net107),
    .X(la_data_out[85]));
 sky130_fd_sc_hd__buf_12 hold80 (.A(net179),
    .X(la_data_out[43]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(net372),
    .X(net180));
 sky130_fd_sc_hd__buf_12 hold82 (.A(net181),
    .X(la_data_out[68]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net354),
    .X(net182));
 sky130_fd_sc_hd__buf_12 hold84 (.A(net183),
    .X(la_data_out[44]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(net328),
    .X(net184));
 sky130_fd_sc_hd__buf_12 hold86 (.A(net185),
    .X(la_data_out[41]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(net396),
    .X(net186));
 sky130_fd_sc_hd__buf_12 hold88 (.A(net187),
    .X(la_data_out[21]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(net336),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net314),
    .X(net108));
 sky130_fd_sc_hd__buf_12 hold90 (.A(net189),
    .X(la_data_out[45]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(net350),
    .X(net190));
 sky130_fd_sc_hd__buf_12 hold92 (.A(net191),
    .X(la_data_out[46]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(net404),
    .X(net192));
 sky130_fd_sc_hd__buf_12 hold94 (.A(net193),
    .X(la_data_out[35]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(net332),
    .X(net194));
 sky130_fd_sc_hd__buf_12 hold96 (.A(net195),
    .X(la_data_out[47]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(net388),
    .X(net196));
 sky130_fd_sc_hd__buf_12 hold98 (.A(net197),
    .X(la_data_out[50]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(net408),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(wb_rst_i),
    .X(net1));
 sky130_fd_sc_hd__buf_6 output10 (.A(net313),
    .X(net125));
 sky130_fd_sc_hd__buf_6 output11 (.A(net289),
    .X(net115));
 sky130_fd_sc_hd__buf_6 output12 (.A(net279),
    .X(net119));
 sky130_fd_sc_hd__buf_6 output13 (.A(net425),
    .X(net265));
 sky130_fd_sc_hd__buf_6 output14 (.A(net403),
    .X(net177));
 sky130_fd_sc_hd__buf_6 output15 (.A(net397),
    .X(net187));
 sky130_fd_sc_hd__buf_6 output16 (.A(net407),
    .X(net203));
 sky130_fd_sc_hd__buf_6 output17 (.A(net359),
    .X(net135));
 sky130_fd_sc_hd__buf_6 output18 (.A(net393),
    .X(net151));
 sky130_fd_sc_hd__buf_6 output19 (.A(net409),
    .X(net199));
 sky130_fd_sc_hd__buf_6 output2 (.A(net449),
    .X(net271));
 sky130_fd_sc_hd__buf_6 output20 (.A(net285),
    .X(net213));
 sky130_fd_sc_hd__buf_6 output21 (.A(net413),
    .X(net215));
 sky130_fd_sc_hd__buf_6 output22 (.A(net417),
    .X(net223));
 sky130_fd_sc_hd__buf_6 output23 (.A(net431),
    .X(net269));
 sky130_fd_sc_hd__buf_6 output24 (.A(net437),
    .X(net261));
 sky130_fd_sc_hd__buf_6 output25 (.A(net445),
    .X(net257));
 sky130_fd_sc_hd__buf_6 output26 (.A(net305),
    .X(net127));
 sky130_fd_sc_hd__buf_6 output27 (.A(net421),
    .X(net205));
 sky130_fd_sc_hd__buf_6 output28 (.A(net319),
    .X(net131));
 sky130_fd_sc_hd__buf_6 output29 (.A(net415),
    .X(net171));
 sky130_fd_sc_hd__buf_6 output3 (.A(net395),
    .X(net237));
 sky130_fd_sc_hd__buf_6 output30 (.A(net405),
    .X(net193));
 sky130_fd_sc_hd__buf_6 output31 (.A(net293),
    .X(net235));
 sky130_fd_sc_hd__buf_6 output32 (.A(net377),
    .X(net211));
 sky130_fd_sc_hd__buf_6 output33 (.A(net347),
    .X(net201));
 sky130_fd_sc_hd__buf_6 output34 (.A(net365),
    .X(net209));
 sky130_fd_sc_hd__buf_6 output35 (.A(net443),
    .X(net273));
 sky130_fd_sc_hd__buf_6 output36 (.A(net411),
    .X(net207));
 sky130_fd_sc_hd__buf_6 output37 (.A(net329),
    .X(net185));
 sky130_fd_sc_hd__buf_6 output38 (.A(net345),
    .X(net175));
 sky130_fd_sc_hd__buf_6 output39 (.A(net335),
    .X(net179));
 sky130_fd_sc_hd__buf_6 output4 (.A(net277),
    .X(net117));
 sky130_fd_sc_hd__buf_6 output40 (.A(net355),
    .X(net183));
 sky130_fd_sc_hd__buf_6 output41 (.A(net337),
    .X(net189));
 sky130_fd_sc_hd__buf_6 output42 (.A(net351),
    .X(net191));
 sky130_fd_sc_hd__buf_6 output43 (.A(net333),
    .X(net195));
 sky130_fd_sc_hd__buf_6 output44 (.A(net295),
    .X(net147));
 sky130_fd_sc_hd__buf_6 output45 (.A(net281),
    .X(net145));
 sky130_fd_sc_hd__buf_6 output46 (.A(net419),
    .X(net247));
 sky130_fd_sc_hd__buf_6 output47 (.A(net389),
    .X(net197));
 sky130_fd_sc_hd__buf_6 output48 (.A(net327),
    .X(net165));
 sky130_fd_sc_hd__buf_6 output49 (.A(net341),
    .X(net159));
 sky130_fd_sc_hd__buf_6 output5 (.A(net325),
    .X(net129));
 sky130_fd_sc_hd__buf_6 output50 (.A(net323),
    .X(net155));
 sky130_fd_sc_hd__buf_6 output51 (.A(net353),
    .X(net167));
 sky130_fd_sc_hd__buf_6 output52 (.A(net331),
    .X(net169));
 sky130_fd_sc_hd__buf_6 output53 (.A(net339),
    .X(net173));
 sky130_fd_sc_hd__buf_6 output54 (.A(net321),
    .X(net163));
 sky130_fd_sc_hd__buf_6 output55 (.A(net297),
    .X(net153));
 sky130_fd_sc_hd__buf_6 output56 (.A(net287),
    .X(net249));
 sky130_fd_sc_hd__buf_6 output57 (.A(net283),
    .X(net245));
 sky130_fd_sc_hd__buf_6 output58 (.A(net429),
    .X(net251));
 sky130_fd_sc_hd__buf_6 output59 (.A(net385),
    .X(net161));
 sky130_fd_sc_hd__buf_6 output6 (.A(net343),
    .X(net123));
 sky130_fd_sc_hd__buf_6 output60 (.A(net357),
    .X(net157));
 sky130_fd_sc_hd__buf_6 output61 (.A(net391),
    .X(net141));
 sky130_fd_sc_hd__buf_6 output62 (.A(net311),
    .X(net143));
 sky130_fd_sc_hd__buf_6 output63 (.A(net349),
    .X(net139));
 sky130_fd_sc_hd__buf_6 output64 (.A(net367),
    .X(net149));
 sky130_fd_sc_hd__buf_6 output65 (.A(net317),
    .X(net137));
 sky130_fd_sc_hd__buf_6 output66 (.A(net373),
    .X(net181));
 sky130_fd_sc_hd__buf_6 output67 (.A(net447),
    .X(net263));
 sky130_fd_sc_hd__buf_6 output68 (.A(net433),
    .X(net255));
 sky130_fd_sc_hd__buf_6 output69 (.A(net439),
    .X(net259));
 sky130_fd_sc_hd__buf_6 output7 (.A(net307),
    .X(net121));
 sky130_fd_sc_hd__buf_6 output70 (.A(net401),
    .X(net239));
 sky130_fd_sc_hd__buf_6 output71 (.A(net361),
    .X(net225));
 sky130_fd_sc_hd__buf_6 output72 (.A(net363),
    .X(net221));
 sky130_fd_sc_hd__buf_6 output73 (.A(net371),
    .X(net217));
 sky130_fd_sc_hd__buf_6 output74 (.A(net379),
    .X(net227));
 sky130_fd_sc_hd__buf_6 output75 (.A(net387),
    .X(net219));
 sky130_fd_sc_hd__buf_6 output76 (.A(net383),
    .X(net231));
 sky130_fd_sc_hd__buf_6 output77 (.A(net399),
    .X(net233));
 sky130_fd_sc_hd__buf_6 output78 (.A(net441),
    .X(net267));
 sky130_fd_sc_hd__buf_6 output79 (.A(net375),
    .X(net229));
 sky130_fd_sc_hd__buf_6 output8 (.A(net291),
    .X(net113));
 sky130_fd_sc_hd__buf_6 output80 (.A(net423),
    .X(net241));
 sky130_fd_sc_hd__buf_6 output81 (.A(net381),
    .X(net111));
 sky130_fd_sc_hd__buf_6 output82 (.A(net315),
    .X(net109));
 sky130_fd_sc_hd__buf_6 output83 (.A(net299),
    .X(net105));
 sky130_fd_sc_hd__buf_6 output84 (.A(net303),
    .X(net101));
 sky130_fd_sc_hd__buf_6 output85 (.A(net309),
    .X(net107));
 sky130_fd_sc_hd__buf_6 output86 (.A(net301),
    .X(net103));
 sky130_fd_sc_hd__buf_6 output87 (.A(net427),
    .X(net243));
 sky130_fd_sc_hd__buf_6 output88 (.A(net451),
    .X(net275));
 sky130_fd_sc_hd__buf_6 output89 (.A(net435),
    .X(net253));
 sky130_fd_sc_hd__buf_6 output9 (.A(net369),
    .X(net133));
 sky130_fd_sc_hd__conb_1 unused_tie_97 (.LO(net97));
 sky130_fd_sc_hd__conb_1 unused_tie_98 (.LO(net98));
 sky130_fd_sc_hd__conb_1 unused_tie_99 (.LO(net99));
 assign irq[0] = net97;
 assign irq[1] = net98;
 assign irq[2] = net99;
endmodule

