// This is the unpowered netlist.
module wrapped_8x305 (rst_n,
    wb_clk_i,
    custom_settings,
    io_in,
    io_oeb,
    io_out);
 input rst_n;
 input wb_clk_i;
 input [1:0] custom_settings;
 input [35:0] io_in;
 output [4:0] io_oeb;
 output [35:0] io_out;

 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire ROM_OEB;
 wire \ROM_addr_buff[10] ;
 wire \ROM_addr_buff[11] ;
 wire \ROM_addr_buff[12] ;
 wire \ROM_addr_buff[13] ;
 wire \ROM_addr_buff[1] ;
 wire \ROM_addr_buff[2] ;
 wire \ROM_addr_buff[3] ;
 wire \ROM_addr_buff[4] ;
 wire \ROM_addr_buff[5] ;
 wire \ROM_addr_buff[6] ;
 wire \ROM_addr_buff[7] ;
 wire \ROM_addr_buff[8] ;
 wire \ROM_addr_buff[9] ;
 wire \ROM_spi_cycle[0] ;
 wire \ROM_spi_cycle[1] ;
 wire \ROM_spi_cycle[2] ;
 wire \ROM_spi_cycle[3] ;
 wire \ROM_spi_cycle[4] ;
 wire \ROM_spi_dat_out[0] ;
 wire \ROM_spi_dat_out[1] ;
 wire \ROM_spi_dat_out[2] ;
 wire \ROM_spi_dat_out[3] ;
 wire \ROM_spi_dat_out[4] ;
 wire \ROM_spi_dat_out[5] ;
 wire \ROM_spi_dat_out[6] ;
 wire \ROM_spi_dat_out[7] ;
 wire ROM_spi_mode;
 wire \S8x305.ALU_in1[0] ;
 wire \S8x305.ALU_in1[1] ;
 wire \S8x305.ALU_in1[2] ;
 wire \S8x305.ALU_in1[3] ;
 wire \S8x305.ALU_in1[4] ;
 wire \S8x305.ALU_in1[5] ;
 wire \S8x305.ALU_in1[6] ;
 wire \S8x305.ALU_in1[7] ;
 wire \S8x305.A[0] ;
 wire \S8x305.A[10] ;
 wire \S8x305.A[11] ;
 wire \S8x305.A[12] ;
 wire \S8x305.A[1] ;
 wire \S8x305.A[2] ;
 wire \S8x305.A[3] ;
 wire \S8x305.A[4] ;
 wire \S8x305.A[5] ;
 wire \S8x305.A[6] ;
 wire \S8x305.A[7] ;
 wire \S8x305.A[8] ;
 wire \S8x305.A[9] ;
 wire \S8x305.I[0] ;
 wire \S8x305.I[10] ;
 wire \S8x305.I[11] ;
 wire \S8x305.I[12] ;
 wire \S8x305.I[13] ;
 wire \S8x305.I[14] ;
 wire \S8x305.I[15] ;
 wire \S8x305.I[1] ;
 wire \S8x305.I[2] ;
 wire \S8x305.I[3] ;
 wire \S8x305.I[4] ;
 wire \S8x305.I[5] ;
 wire \S8x305.I[6] ;
 wire \S8x305.I[7] ;
 wire \S8x305.I[8] ;
 wire \S8x305.I[9] ;
 wire \S8x305.PC[0] ;
 wire \S8x305.PC[10] ;
 wire \S8x305.PC[11] ;
 wire \S8x305.PC[12] ;
 wire \S8x305.PC[1] ;
 wire \S8x305.PC[2] ;
 wire \S8x305.PC[3] ;
 wire \S8x305.PC[4] ;
 wire \S8x305.PC[5] ;
 wire \S8x305.PC[6] ;
 wire \S8x305.PC[7] ;
 wire \S8x305.PC[8] ;
 wire \S8x305.PC[9] ;
 wire \S8x305.cycle[0] ;
 wire \S8x305.cycle[1] ;
 wire \S8x305.i_latch[0] ;
 wire \S8x305.i_latch[10] ;
 wire \S8x305.i_latch[11] ;
 wire \S8x305.i_latch[12] ;
 wire \S8x305.i_latch[13] ;
 wire \S8x305.i_latch[14] ;
 wire \S8x305.i_latch[15] ;
 wire \S8x305.i_latch[1] ;
 wire \S8x305.i_latch[2] ;
 wire \S8x305.i_latch[3] ;
 wire \S8x305.i_latch[4] ;
 wire \S8x305.i_latch[5] ;
 wire \S8x305.i_latch[6] ;
 wire \S8x305.i_latch[7] ;
 wire \S8x305.i_latch[8] ;
 wire \S8x305.i_latch[9] ;
 wire \S8x305.iv_latch[0] ;
 wire \S8x305.iv_latch[1] ;
 wire \S8x305.iv_latch[2] ;
 wire \S8x305.iv_latch[3] ;
 wire \S8x305.iv_latch[4] ;
 wire \S8x305.iv_latch[5] ;
 wire \S8x305.iv_latch[6] ;
 wire \S8x305.iv_latch[7] ;
 wire \S8x305.regs[10][0] ;
 wire \S8x305.regs[10][1] ;
 wire \S8x305.regs[10][2] ;
 wire \S8x305.regs[10][3] ;
 wire \S8x305.regs[10][4] ;
 wire \S8x305.regs[10][5] ;
 wire \S8x305.regs[10][6] ;
 wire \S8x305.regs[10][7] ;
 wire \S8x305.regs[11][0] ;
 wire \S8x305.regs[11][1] ;
 wire \S8x305.regs[11][2] ;
 wire \S8x305.regs[11][3] ;
 wire \S8x305.regs[11][4] ;
 wire \S8x305.regs[11][5] ;
 wire \S8x305.regs[11][6] ;
 wire \S8x305.regs[11][7] ;
 wire \S8x305.regs[12][0] ;
 wire \S8x305.regs[12][1] ;
 wire \S8x305.regs[12][2] ;
 wire \S8x305.regs[12][3] ;
 wire \S8x305.regs[12][4] ;
 wire \S8x305.regs[12][5] ;
 wire \S8x305.regs[12][6] ;
 wire \S8x305.regs[12][7] ;
 wire \S8x305.regs[13][0] ;
 wire \S8x305.regs[13][1] ;
 wire \S8x305.regs[13][2] ;
 wire \S8x305.regs[13][3] ;
 wire \S8x305.regs[13][4] ;
 wire \S8x305.regs[13][5] ;
 wire \S8x305.regs[13][6] ;
 wire \S8x305.regs[13][7] ;
 wire \S8x305.regs[14][0] ;
 wire \S8x305.regs[14][1] ;
 wire \S8x305.regs[14][2] ;
 wire \S8x305.regs[14][3] ;
 wire \S8x305.regs[14][4] ;
 wire \S8x305.regs[14][5] ;
 wire \S8x305.regs[14][6] ;
 wire \S8x305.regs[14][7] ;
 wire \S8x305.regs[15][0] ;
 wire \S8x305.regs[15][1] ;
 wire \S8x305.regs[15][2] ;
 wire \S8x305.regs[15][3] ;
 wire \S8x305.regs[15][4] ;
 wire \S8x305.regs[15][5] ;
 wire \S8x305.regs[15][6] ;
 wire \S8x305.regs[15][7] ;
 wire \S8x305.regs[1][0] ;
 wire \S8x305.regs[1][1] ;
 wire \S8x305.regs[1][2] ;
 wire \S8x305.regs[1][3] ;
 wire \S8x305.regs[1][4] ;
 wire \S8x305.regs[1][5] ;
 wire \S8x305.regs[1][6] ;
 wire \S8x305.regs[1][7] ;
 wire \S8x305.regs[2][0] ;
 wire \S8x305.regs[2][1] ;
 wire \S8x305.regs[2][2] ;
 wire \S8x305.regs[2][3] ;
 wire \S8x305.regs[2][4] ;
 wire \S8x305.regs[2][5] ;
 wire \S8x305.regs[2][6] ;
 wire \S8x305.regs[2][7] ;
 wire \S8x305.regs[3][0] ;
 wire \S8x305.regs[3][1] ;
 wire \S8x305.regs[3][2] ;
 wire \S8x305.regs[3][3] ;
 wire \S8x305.regs[3][4] ;
 wire \S8x305.regs[3][5] ;
 wire \S8x305.regs[3][6] ;
 wire \S8x305.regs[3][7] ;
 wire \S8x305.regs[4][0] ;
 wire \S8x305.regs[4][1] ;
 wire \S8x305.regs[4][2] ;
 wire \S8x305.regs[4][3] ;
 wire \S8x305.regs[4][4] ;
 wire \S8x305.regs[4][5] ;
 wire \S8x305.regs[4][6] ;
 wire \S8x305.regs[4][7] ;
 wire \S8x305.regs[5][0] ;
 wire \S8x305.regs[5][1] ;
 wire \S8x305.regs[5][2] ;
 wire \S8x305.regs[5][3] ;
 wire \S8x305.regs[5][4] ;
 wire \S8x305.regs[5][5] ;
 wire \S8x305.regs[5][6] ;
 wire \S8x305.regs[5][7] ;
 wire \S8x305.regs[6][0] ;
 wire \S8x305.regs[6][1] ;
 wire \S8x305.regs[6][2] ;
 wire \S8x305.regs[6][3] ;
 wire \S8x305.regs[6][4] ;
 wire \S8x305.regs[6][5] ;
 wire \S8x305.regs[6][6] ;
 wire \S8x305.regs[6][7] ;
 wire \S8x305.regs[7][0] ;
 wire \S8x305.regs[7][1] ;
 wire \S8x305.regs[7][2] ;
 wire \S8x305.regs[7][3] ;
 wire \S8x305.regs[7][4] ;
 wire \S8x305.regs[7][5] ;
 wire \S8x305.regs[7][6] ;
 wire \S8x305.regs[7][7] ;
 wire \S8x305.regs[8][0] ;
 wire \S8x305.regs[8][1] ;
 wire \S8x305.regs[8][2] ;
 wire \S8x305.regs[8][3] ;
 wire \S8x305.regs[8][4] ;
 wire \S8x305.regs[8][5] ;
 wire \S8x305.regs[8][6] ;
 wire \S8x305.regs[8][7] ;
 wire \S8x305.regs[9][0] ;
 wire \S8x305.regs[9][1] ;
 wire \S8x305.regs[9][2] ;
 wire \S8x305.regs[9][3] ;
 wire \S8x305.regs[9][4] ;
 wire \S8x305.regs[9][5] ;
 wire \S8x305.regs[9][6] ;
 wire \S8x305.regs[9][7] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire clknet_0_wb_clk_i;
 wire clknet_2_0__leaf_wb_clk_i;
 wire clknet_2_1__leaf_wb_clk_i;
 wire clknet_2_2__leaf_wb_clk_i;
 wire clknet_2_3__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire \cmdl[0] ;
 wire \cmdl[1] ;
 wire \cmdl[2] ;
 wire \cmdl[3] ;
 wire \cmdl[4] ;
 wire \cmdl[5] ;
 wire \cmdl[6] ;
 wire \cmdl[7] ;
 wire \cmdr[0] ;
 wire \cmdr[1] ;
 wire \cmdr[2] ;
 wire \cmdr[3] ;
 wire \cmdr[4] ;
 wire \cmdr[5] ;
 wire \cmdr[6] ;
 wire \cmdr[7] ;
 wire \last_A[10] ;
 wire \last_A[11] ;
 wire \last_A[12] ;
 wire \last_A[1] ;
 wire \last_A[2] ;
 wire \last_A[3] ;
 wire \last_A[4] ;
 wire \last_A[5] ;
 wire \last_A[6] ;
 wire \last_A[7] ;
 wire \last_A[9] ;
 wire \last_addr[0] ;
 wire \last_addr[10] ;
 wire \last_addr[11] ;
 wire \last_addr[12] ;
 wire \last_addr[13] ;
 wire \last_addr[1] ;
 wire \last_addr[2] ;
 wire \last_addr[3] ;
 wire \last_addr[4] ;
 wire \last_addr[5] ;
 wire \last_addr[6] ;
 wire \last_addr[7] ;
 wire \last_addr[8] ;
 wire \last_addr[9] ;
 wire \mem_cycle[0] ;
 wire \mem_cycle[1] ;
 wire \mem_cycle[2] ;
 wire \mem_cycle[3] ;
 wire \mem_cycle[4] ;
 wire \mem_cycle[5] ;
 wire \memory[0][0] ;
 wire \memory[0][1] ;
 wire \memory[0][2] ;
 wire \memory[0][3] ;
 wire \memory[0][4] ;
 wire \memory[0][5] ;
 wire \memory[0][6] ;
 wire \memory[0][7] ;
 wire \memory[10][0] ;
 wire \memory[10][1] ;
 wire \memory[10][2] ;
 wire \memory[10][3] ;
 wire \memory[10][4] ;
 wire \memory[10][5] ;
 wire \memory[10][6] ;
 wire \memory[10][7] ;
 wire \memory[11][0] ;
 wire \memory[11][1] ;
 wire \memory[11][2] ;
 wire \memory[11][3] ;
 wire \memory[11][4] ;
 wire \memory[11][5] ;
 wire \memory[11][6] ;
 wire \memory[11][7] ;
 wire \memory[12][0] ;
 wire \memory[12][1] ;
 wire \memory[12][2] ;
 wire \memory[12][3] ;
 wire \memory[12][4] ;
 wire \memory[12][5] ;
 wire \memory[12][6] ;
 wire \memory[12][7] ;
 wire \memory[13][0] ;
 wire \memory[13][1] ;
 wire \memory[13][2] ;
 wire \memory[13][3] ;
 wire \memory[13][4] ;
 wire \memory[13][5] ;
 wire \memory[13][6] ;
 wire \memory[13][7] ;
 wire \memory[14][0] ;
 wire \memory[14][1] ;
 wire \memory[14][2] ;
 wire \memory[14][3] ;
 wire \memory[14][4] ;
 wire \memory[14][5] ;
 wire \memory[14][6] ;
 wire \memory[14][7] ;
 wire \memory[15][0] ;
 wire \memory[15][1] ;
 wire \memory[15][2] ;
 wire \memory[15][3] ;
 wire \memory[15][4] ;
 wire \memory[15][5] ;
 wire \memory[15][6] ;
 wire \memory[15][7] ;
 wire \memory[1][0] ;
 wire \memory[1][1] ;
 wire \memory[1][2] ;
 wire \memory[1][3] ;
 wire \memory[1][4] ;
 wire \memory[1][5] ;
 wire \memory[1][6] ;
 wire \memory[1][7] ;
 wire \memory[2][0] ;
 wire \memory[2][1] ;
 wire \memory[2][2] ;
 wire \memory[2][3] ;
 wire \memory[2][4] ;
 wire \memory[2][5] ;
 wire \memory[2][6] ;
 wire \memory[2][7] ;
 wire \memory[3][0] ;
 wire \memory[3][1] ;
 wire \memory[3][2] ;
 wire \memory[3][3] ;
 wire \memory[3][4] ;
 wire \memory[3][5] ;
 wire \memory[3][6] ;
 wire \memory[3][7] ;
 wire \memory[4][0] ;
 wire \memory[4][1] ;
 wire \memory[4][2] ;
 wire \memory[4][3] ;
 wire \memory[4][4] ;
 wire \memory[4][5] ;
 wire \memory[4][6] ;
 wire \memory[4][7] ;
 wire \memory[5][0] ;
 wire \memory[5][1] ;
 wire \memory[5][2] ;
 wire \memory[5][3] ;
 wire \memory[5][4] ;
 wire \memory[5][5] ;
 wire \memory[5][6] ;
 wire \memory[5][7] ;
 wire \memory[6][0] ;
 wire \memory[6][1] ;
 wire \memory[6][2] ;
 wire \memory[6][3] ;
 wire \memory[6][4] ;
 wire \memory[6][5] ;
 wire \memory[6][6] ;
 wire \memory[6][7] ;
 wire \memory[7][0] ;
 wire \memory[7][1] ;
 wire \memory[7][2] ;
 wire \memory[7][3] ;
 wire \memory[7][4] ;
 wire \memory[7][5] ;
 wire \memory[7][6] ;
 wire \memory[7][7] ;
 wire \memory[8][0] ;
 wire \memory[8][1] ;
 wire \memory[8][2] ;
 wire \memory[8][3] ;
 wire \memory[8][4] ;
 wire \memory[8][5] ;
 wire \memory[8][6] ;
 wire \memory[8][7] ;
 wire \memory[9][0] ;
 wire \memory[9][1] ;
 wire \memory[9][2] ;
 wire \memory[9][3] ;
 wire \memory[9][4] ;
 wire \memory[9][5] ;
 wire \memory[9][6] ;
 wire \memory[9][7] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net12;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire spi_clkdiv;
 wire \startup_cycle[0] ;
 wire \startup_cycle[1] ;
 wire \startup_cycle[2] ;
 wire \startup_cycle[3] ;
 wire \startup_cycle[4] ;
 wire \startup_cycle[5] ;
 wire \startup_cycle[6] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\memory[11][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_0300_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_1004_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net351));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA__1862__A (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__1863__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__1864__A (.DIODE(\S8x305.iv_latch[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1865__A (.DIODE(\S8x305.iv_latch[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1866__A (.DIODE(\S8x305.iv_latch[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1868__A (.DIODE(\S8x305.iv_latch[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1906__B (.DIODE(_1796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1910__C (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__1912__A2 (.DIODE(_1796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1912__B1 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1915__A (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1920__C (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__1921__A2 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1922__A2 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1923__A2 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1928__A2 (.DIODE(_1796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1932__A2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__1937__A0 (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1937__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__1938__B (.DIODE(_1796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1939__A (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1940__A (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1943__A (.DIODE(_1816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1943__B (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1945__A (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1945__B (.DIODE(_1796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1946__A2 (.DIODE(_1837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1948__A (.DIODE(_1816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1948__B (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1953__A1 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1956__A (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1959__B (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__1959__C (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1962__D (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1969__A2 (.DIODE(_1796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1969__A3 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__1969__B1 (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1970__A2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__1970__A3 (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1975__A1 (.DIODE(_1816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1975__A2 (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1982__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__1985__B (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1985__C (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1987__B (.DIODE(_1796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1992__A1 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1993__A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1993__S (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__1994__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__1998__S (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__2000__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2007__B (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2010__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2010__C (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2011__A3 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2015__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2018__S (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__2019__S (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__2020__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__2022__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2023__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__2024__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__2025__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__2026__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2026__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__2027__A1 (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2029__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2032__S (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__2033__S (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__2034__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2035__S (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__2036__S (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__2037__S (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__2038__S (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__2039__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__2041__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2042__S (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__2043__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__2044__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__2044__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__2045__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2046__A1 (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2048__A1 (.DIODE(\S8x305.iv_latch[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2052__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2053__S (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__2054__S (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__2055__S (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__2056__S (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__2059__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2060__S (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__2061__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__2062__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__2063__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2063__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__2064__A1 (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2067__A1 (.DIODE(\S8x305.iv_latch[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2068__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2070__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2071__S (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__2073__S (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__2074__S (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__2075__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__2077__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2078__S (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__2079__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__2080__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__2081__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2081__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__2082__A1 (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2085__A1 (.DIODE(\S8x305.iv_latch[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2088__A1 (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2089__A0 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__2089__S (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__2090__A1 (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2091__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__2095__S (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__2096__S (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__2097__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2098__S (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__2099__S (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__2100__S (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__2101__S (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__2104__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2105__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__2106__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__2107__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__2108__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2108__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__2109__A1 (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2113__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2115__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2117__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2118__S (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__2119__S (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__2122__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2123__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__2124__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__2125__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__2126__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2126__B1 (.DIODE(_1829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2127__A1 (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2129__C (.DIODE(_0606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2131__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2133__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2136__S (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__2137__S (.DIODE(_1829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2140__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2141__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__2142__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__2143__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__2144__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2144__B1 (.DIODE(_1829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2145__A1 (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2148__A1 (.DIODE(\S8x305.iv_latch[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2151__S (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2153__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2154__S (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2155__S (.DIODE(_1829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2156__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__2158__S (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2159__S (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__2160__A (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2161__S (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__2162__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2162__B1 (.DIODE(_1829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2163__A1 (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2173__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__2176__S (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__2180__A (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2180__B (.DIODE(_1796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2182__A1 (.DIODE(_1837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2182__B2 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2183__A1 (.DIODE(\S8x305.iv_latch[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2184__A1 (.DIODE(\S8x305.iv_latch[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2193__A1 (.DIODE(\S8x305.iv_latch[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2202__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__2204__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__2212__B (.DIODE(_0606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2216__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2217__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__2231__A1 (.DIODE(\S8x305.iv_latch[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2232__S (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2242__C1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__2243__A1 (.DIODE(\S8x305.iv_latch[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2244__A1 (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2253__B2 (.DIODE(\S8x305.iv_latch[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2254__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__2267__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__2270__B2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__2271__A1_N (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__2277__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__2278__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__2292__B1 (.DIODE(_1796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2296__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__2296__B (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2297__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__2297__B1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2309__A1 (.DIODE(_1837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2309__B2 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2311__B1 (.DIODE(_1796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2315__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__2322__A1 (.DIODE(_1837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2322__B2 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2325__C1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2327__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__2328__B (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2330__A1 (.DIODE(_1837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2330__B2 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2331__A1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2333__B1 (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2334__C1 (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2340__A1 (.DIODE(_1837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2340__B2 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2343__A0 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2344__B1 (.DIODE(_1837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2345__A1 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2346__A0 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2349__A (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2351__A1_N (.DIODE(_1837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2353__B1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2354__A1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2357__A1 (.DIODE(_1837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2357__B2 (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2362__A0 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2368__A2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__2383__A2 (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2384__A2 (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2392__B (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2396__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__2396__C_N (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2397__S0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2397__S1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__2399__S0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2399__S1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2401__S0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2401__S1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2403__S0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2403__S1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__2410__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__2411__S (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2433__A1 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__2438__C1 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2440__S0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2440__S1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__2442__S0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2442__S1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2444__S0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2444__S1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2446__S0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2446__S1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__2450__S (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2452__A1 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__2452__C1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2461__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2462__B1 (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2463__A1 (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2463__B1 (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2467__S0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2467__S1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2469__S0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2469__S1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2471__S0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2473__S0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2473__S1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__2477__S (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2479__A1 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2480__A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__2480__C1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2488__B1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__2489__A1 (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2492__C1 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2494__S0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2494__S1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__2496__S0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2496__S1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2498__S0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2498__S1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2500__S0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2500__S1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__2504__S (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2506__C1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__2510__A2 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2513__C1 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2515__S0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2515__S1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__2517__S0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2517__S1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2519__S0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2519__S1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2521__S0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2521__S1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__2525__S (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2527__C1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__2530__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2531__A2 (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2534__C1 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2536__S0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2536__S1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__2538__S0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2540__S0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2540__S1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2542__S0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2542__S1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__2546__S (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2553__A1 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2555__C1 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2557__S0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2557__S1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__2559__S0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2559__S1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2561__S0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2561__S1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2563__S0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2563__S1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__2567__S (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2569__C1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__2572__A0 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA__2573__A0 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2576__C1 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2578__S0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2578__S1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2580__S0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__2580__S1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2582__S0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2582__S1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2584__S0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2584__S1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__2588__S (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2590__A1 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA__2590__C1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__2591__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__2592__C (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__2596__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__2597__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__2598__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2599__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2600__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2601__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2602__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2603__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2607__B (.DIODE(_0606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2610__B (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2612__B (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2616__A (.DIODE(_1787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2631__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__2635__A1 (.DIODE(_1828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2643__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__2646__A (.DIODE(_1771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2646__C (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__2646__D (.DIODE(_0487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2648__A (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2649__A1 (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2649__B1 (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2650__A1 (.DIODE(_1825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2650__B1 (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2655__S (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2656__A2 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2658__S (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2659__A2 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2661__S (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2662__A2 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2664__S (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2665__A2 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2667__S (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2668__A2 (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2670__B (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2671__A2 (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2672__A2 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2673__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2674__S (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2675__A2 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2676__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2677__B (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2679__A2 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2683__A1 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA__2693__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2695__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2696__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2697__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2698__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2699__A1 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2701__A1 (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2703__A1 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2704__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2705__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2706__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2707__A1 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2708__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__2713__B2 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2714__B2 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2715__B2 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2716__B2 (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2717__B2 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2718__B2 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2719__B2 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2721__A1 (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2722__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__2725__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2731__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2736__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2737__C (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2738__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2741__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2744__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2745__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2747__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2749__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2751__A1 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2753__A1 (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2754__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2755__A1 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2756__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2757__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2758__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2759__A1 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2761__A (.DIODE(_1816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2762__A (.DIODE(_1816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2763__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2764__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2766__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2768__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2770__A1 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2772__A1 (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2774__A1 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2776__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2777__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2778__A1 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2779__A (.DIODE(_1816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2780__A (.DIODE(_1816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2781__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2782__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2784__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2786__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2788__A1 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2790__A1 (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2791__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2792__A1 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2794__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2795__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2796__A1 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2799__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2800__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2802__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2804__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2806__A1 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2808__A1 (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2810__A1 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2812__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2813__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2814__A1 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2818__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2820__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2822__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2824__A1 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2826__A1 (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2828__A1 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2830__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2832__A1 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2838__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2840__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2842__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2844__A1 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2846__A1 (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2848__A1 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2850__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2852__A1 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2856__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2858__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2860__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2862__A1 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2864__A1 (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2866__A1 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2868__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2870__A1 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2873__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2874__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2875__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2876__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2877__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2878__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2879__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2880__A1 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2881__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2882__A1 (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2883__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2884__A1 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2885__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2886__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2887__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2888__A1 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2926__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__2928__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__2930__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__2932__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__2939__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__2941__A2 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2941__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__2942__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2942__A2 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2943__A1 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__2943__A2 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2943__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__2944__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2944__A2 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2945__A2 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2945__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__2946__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2946__A2 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2947__A1 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA__2947__A2 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2947__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__2948__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2948__A2 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2949__A2 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2949__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__2950__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2950__A2 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2951__A2 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2951__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__2952__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2952__A2 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2953__A2 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2953__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__2954__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__2954__A2 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2955__A2 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2956__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__2956__A2 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2979__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__2999__C1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3002__D1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3007__C1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3062__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3071__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3091__C1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3139__C1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3141__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3172__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3184__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3186__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3188__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3190__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3202__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__3203__A1 (.DIODE(\S8x305.iv_latch[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3204__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__3206__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__3207__A1 (.DIODE(\S8x305.iv_latch[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3208__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__A1 (.DIODE(\S8x305.iv_latch[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3210__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__3211__A1 (.DIODE(\S8x305.iv_latch[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3212__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__3213__A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__3214__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__3215__A1 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__3216__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__3219__A1 (.DIODE(\S8x305.iv_latch[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3221__A1 (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__3223__A1 (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__3249__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3250__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3251__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3252__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3253__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3254__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3255__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3256__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3260__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3262__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3264__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3266__A1 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3268__A1 (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3270__A1 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3272__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3274__A1 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3277__A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__3281__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__A0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__3286__A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__3288__A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__3290__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__3291__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3292__A0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__3293__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3295__A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__3297__A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__3299__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__3301__A0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__3315__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3320__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3322__A (.DIODE(_1816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3325__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3327__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3329__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3331__A1 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3333__A1 (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3335__A1 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3337__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3339__A1 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3343__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3345__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3347__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3349__A1 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3351__A1 (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3353__A1 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3355__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3357__A1 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3361__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3363__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3365__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3367__A1 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3369__A1 (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3371__A1 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3373__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3375__A1 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3377__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3378__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3380__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3381__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3382__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3383__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3384__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3389__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3390__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3391__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3393__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3394__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3396__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3399__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3399__S (.DIODE(_1607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3400__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3400__S (.DIODE(_1607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3401__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3401__S (.DIODE(_1607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__S (.DIODE(_1607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3403__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3403__S (.DIODE(_1607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3404__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3404__S (.DIODE(_1607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3405__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3405__S (.DIODE(_1607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3406__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3406__S (.DIODE(_1607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3409__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3410__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3411__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3412__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3413__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3414__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3415__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3416__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3418__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3419__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3420__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3421__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3423__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3425__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3430__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3431__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3432__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3433__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3438__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3440__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3442__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3443__A0 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__3444__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3448__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3450__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3452__A0 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__3453__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3456__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3457__A (.DIODE(_1771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__A (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__C1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA__3461__C1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3462__A (.DIODE(\S8x305.iv_latch[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3463__C1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__A (.DIODE(\S8x305.iv_latch[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3465__C1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3467__A (.DIODE(_1771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3469__C1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__A (.DIODE(\S8x305.iv_latch[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3471__C1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__A (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__A (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3503__A1 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__A1 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__A (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3507__A (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3508__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__3513__A (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3514__A (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3516__A1 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__A (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3519__A1 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3519__B2 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__S (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__A (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3526__A1 (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__A1 (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__A (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__S (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__A1 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__A1 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__A (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3540__A (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3541__A1 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3542__A1 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3544__S (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__3548__A1 (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3549__A1 (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__A (.DIODE(_0606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__B (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__A (.DIODE(_0606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__B (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__C1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__C1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__B (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3573__B (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__A2 (.DIODE(_0487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__B (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__B (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__A2 (.DIODE(_0487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__B (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__A2 (.DIODE(_0487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3585__B2 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3590__A1 (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3594__A1 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__C1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__B1 (.DIODE(_1771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3606__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3607__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3608__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3609__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3611__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__A0 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__3617__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3620__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3623__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__A0 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__3625__A0 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3627__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3630__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3634__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3636__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3639__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3643__A1 (.DIODE(_1112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3645__A1 (.DIODE(_1114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__A1 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3649__A1 (.DIODE(_1118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__A1 (.DIODE(_1120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3653__A1 (.DIODE(_1123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__A1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3657__A1 (.DIODE(_1128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3659__A0 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3660__A0 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3661__A0 (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3662__A0 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3663__A0 (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3667__A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3669__A0 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__A0 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__A0 (.DIODE(_1796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__S (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__A0 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__S (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__A0 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__S (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__S (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3680__S (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__S (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3682__S (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__S (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__A1 (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__D (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__D (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout101_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout102_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout103_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_A (.DIODE(_1829_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout62_A (.DIODE(_1802_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout65_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_A (.DIODE(_1824_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout67_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout69_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout87_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout89_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout91_A (.DIODE(_1771_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_A (.DIODE(_1771_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout94_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout95_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout97_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold368_A (.DIODE(_0487_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold478_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold479_A (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold499_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold536_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold547_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold559_A (.DIODE(\S8x305.iv_latch[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold609_A (.DIODE(\S8x305.iv_latch[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold638_A (.DIODE(\S8x305.iv_latch[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold688_A (.DIODE(\S8x305.iv_latch[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_output24_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_output30_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_output31_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_output32_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_output35_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_output40_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_output44_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_output46_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_output47_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_output50_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_output51_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_output52_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_output53_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_output54_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_output55_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_output56_A (.DIODE(net75));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__inv_2 _1838_ (.A(net599),
    .Y(_1740_));
 sky130_fd_sc_hd__inv_2 _1839_ (.A(net453),
    .Y(_1741_));
 sky130_fd_sc_hd__inv_2 _1840_ (.A(net494),
    .Y(_1742_));
 sky130_fd_sc_hd__inv_2 _1841_ (.A(net672),
    .Y(_1743_));
 sky130_fd_sc_hd__inv_2 _1842_ (.A(net753),
    .Y(_1744_));
 sky130_fd_sc_hd__inv_2 _1843_ (.A(net639),
    .Y(_1745_));
 sky130_fd_sc_hd__inv_2 _1844_ (.A(net483),
    .Y(_1746_));
 sky130_fd_sc_hd__inv_2 _1845_ (.A(net543),
    .Y(_1747_));
 sky130_fd_sc_hd__inv_2 _1846_ (.A(net455),
    .Y(_1748_));
 sky130_fd_sc_hd__inv_2 _1847_ (.A(\S8x305.A[1] ),
    .Y(_1749_));
 sky130_fd_sc_hd__inv_2 _1848_ (.A(\S8x305.A[0] ),
    .Y(_1750_));
 sky130_fd_sc_hd__inv_2 _1849_ (.A(\ROM_addr_buff[9] ),
    .Y(_1751_));
 sky130_fd_sc_hd__inv_2 _1850_ (.A(\ROM_addr_buff[1] ),
    .Y(_1752_));
 sky130_fd_sc_hd__inv_2 _1851_ (.A(\S8x305.I[12] ),
    .Y(_1753_));
 sky130_fd_sc_hd__inv_2 _1852_ (.A(net708),
    .Y(_1754_));
 sky130_fd_sc_hd__inv_2 _1853_ (.A(net724),
    .Y(_1755_));
 sky130_fd_sc_hd__inv_2 _1854_ (.A(net836),
    .Y(_1756_));
 sky130_fd_sc_hd__inv_2 _1855_ (.A(\last_A[9] ),
    .Y(_1757_));
 sky130_fd_sc_hd__inv_2 _1856_ (.A(\last_A[5] ),
    .Y(_1758_));
 sky130_fd_sc_hd__inv_2 _1857_ (.A(\last_A[4] ),
    .Y(_1759_));
 sky130_fd_sc_hd__inv_2 _1858_ (.A(\last_A[3] ),
    .Y(_1760_));
 sky130_fd_sc_hd__inv_2 _1859_ (.A(\last_A[2] ),
    .Y(_1761_));
 sky130_fd_sc_hd__inv_2 _1860_ (.A(net751),
    .Y(_1762_));
 sky130_fd_sc_hd__inv_2 _1861_ (.A(\S8x305.iv_latch[7] ),
    .Y(net50));
 sky130_fd_sc_hd__inv_2 _1862_ (.A(net400),
    .Y(net51));
 sky130_fd_sc_hd__inv_2 _1863_ (.A(net429),
    .Y(net52));
 sky130_fd_sc_hd__inv_2 _1864_ (.A(\S8x305.iv_latch[4] ),
    .Y(net53));
 sky130_fd_sc_hd__inv_2 _1865_ (.A(\S8x305.iv_latch[3] ),
    .Y(net54));
 sky130_fd_sc_hd__inv_2 _1866_ (.A(\S8x305.iv_latch[2] ),
    .Y(net55));
 sky130_fd_sc_hd__inv_2 _1867_ (.A(\S8x305.iv_latch[1] ),
    .Y(net56));
 sky130_fd_sc_hd__inv_2 _1868_ (.A(\S8x305.iv_latch[0] ),
    .Y(net30));
 sky130_fd_sc_hd__inv_2 _1869_ (.A(net826),
    .Y(_1763_));
 sky130_fd_sc_hd__inv_2 _1870_ (.A(net822),
    .Y(_1764_));
 sky130_fd_sc_hd__inv_2 _1871_ (.A(net443),
    .Y(_1765_));
 sky130_fd_sc_hd__inv_2 _1872_ (.A(\mem_cycle[0] ),
    .Y(_1766_));
 sky130_fd_sc_hd__inv_2 _1873_ (.A(net720),
    .Y(_1767_));
 sky130_fd_sc_hd__inv_2 _1874_ (.A(net661),
    .Y(_1768_));
 sky130_fd_sc_hd__inv_2 _1875_ (.A(net768),
    .Y(_1769_));
 sky130_fd_sc_hd__inv_2 _1876_ (.A(net688),
    .Y(_1770_));
 sky130_fd_sc_hd__inv_2 _1877_ (.A(net99),
    .Y(_1771_));
 sky130_fd_sc_hd__inv_2 _1878_ (.A(\S8x305.ALU_in1[1] ),
    .Y(_1772_));
 sky130_fd_sc_hd__inv_2 _1879_ (.A(net771),
    .Y(_1773_));
 sky130_fd_sc_hd__inv_2 _1880_ (.A(net3),
    .Y(_1774_));
 sky130_fd_sc_hd__inv_2 _1881_ (.A(net22),
    .Y(_1775_));
 sky130_fd_sc_hd__inv_2 _1882_ (.A(net21),
    .Y(_1776_));
 sky130_fd_sc_hd__inv_2 _1883_ (.A(net20),
    .Y(_1777_));
 sky130_fd_sc_hd__inv_2 _1884_ (.A(net19),
    .Y(_1778_));
 sky130_fd_sc_hd__inv_2 _1885_ (.A(net18),
    .Y(_1779_));
 sky130_fd_sc_hd__inv_2 _1886_ (.A(net17),
    .Y(_1780_));
 sky130_fd_sc_hd__inv_2 _1887_ (.A(net16),
    .Y(_1781_));
 sky130_fd_sc_hd__nand2_2 _1888_ (.A(net82),
    .B(net84),
    .Y(_1782_));
 sky130_fd_sc_hd__clkinv_4 _1889_ (.A(_1782_),
    .Y(net35));
 sky130_fd_sc_hd__nor2_8 _1890_ (.A(net82),
    .B(net84),
    .Y(_1783_));
 sky130_fd_sc_hd__or2_4 _1891_ (.A(net82),
    .B(net84),
    .X(_1784_));
 sky130_fd_sc_hd__o21bai_4 _1892_ (.A1(net83),
    .A2(net84),
    .B1_N(net459),
    .Y(_1785_));
 sky130_fd_sc_hd__or3_4 _1893_ (.A(net83),
    .B(net84),
    .C(\S8x305.I[13] ),
    .X(_1786_));
 sky130_fd_sc_hd__nand2_4 _1894_ (.A(_1785_),
    .B(_1786_),
    .Y(_1787_));
 sky130_fd_sc_hd__and2_2 _1895_ (.A(_1785_),
    .B(_1786_),
    .X(_1788_));
 sky130_fd_sc_hd__o21ba_2 _1896_ (.A1(net82),
    .A2(net84),
    .B1_N(net158),
    .X(_1789_));
 sky130_fd_sc_hd__nor3_2 _1897_ (.A(net82),
    .B(net84),
    .C(\S8x305.I[15] ),
    .Y(_1790_));
 sky130_fd_sc_hd__or2_2 _1898_ (.A(_1789_),
    .B(_1790_),
    .X(_1791_));
 sky130_fd_sc_hd__nor2_2 _1899_ (.A(_1789_),
    .B(_1790_),
    .Y(_1792_));
 sky130_fd_sc_hd__a211oi_4 _1900_ (.A1(_1785_),
    .A2(_1786_),
    .B1(_1789_),
    .C1(_1790_),
    .Y(_1793_));
 sky130_fd_sc_hd__a211o_2 _1901_ (.A1(_1785_),
    .A2(_1786_),
    .B1(_1789_),
    .C1(_1790_),
    .X(_1794_));
 sky130_fd_sc_hd__or3_2 _1902_ (.A(net82),
    .B(net84),
    .C(net663),
    .X(_1795_));
 sky130_fd_sc_hd__o21a_4 _1903_ (.A1(net760),
    .A2(_1783_),
    .B1(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__o21ai_4 _1904_ (.A1(\S8x305.i_latch[14] ),
    .A2(_1783_),
    .B1(_1795_),
    .Y(_1797_));
 sky130_fd_sc_hd__nor2_1 _1905_ (.A(_1794_),
    .B(_1797_),
    .Y(_1798_));
 sky130_fd_sc_hd__nand2_8 _1906_ (.A(_1793_),
    .B(_1796_),
    .Y(_1799_));
 sky130_fd_sc_hd__or2_1 _1907_ (.A(\S8x305.I[9] ),
    .B(_1784_),
    .X(_1800_));
 sky130_fd_sc_hd__mux2_1 _1908_ (.A0(\S8x305.I[9] ),
    .A1(net686),
    .S(_1784_),
    .X(_1801_));
 sky130_fd_sc_hd__o21ai_4 _1909_ (.A1(\S8x305.i_latch[9] ),
    .A2(_1783_),
    .B1(_1800_),
    .Y(_1802_));
 sky130_fd_sc_hd__or3_2 _1910_ (.A(_1794_),
    .B(_1797_),
    .C(net72),
    .X(_1803_));
 sky130_fd_sc_hd__mux2_8 _1911_ (.A0(net746),
    .A1(net390),
    .S(_1784_),
    .X(_1804_));
 sky130_fd_sc_hd__a21o_1 _1912_ (.A1(_1793_),
    .A2(_1796_),
    .B1(_1804_),
    .X(_1805_));
 sky130_fd_sc_hd__and2_2 _1913_ (.A(_1803_),
    .B(_1805_),
    .X(_1806_));
 sky130_fd_sc_hd__mux2_8 _1914_ (.A0(net772),
    .A1(net437),
    .S(_1784_),
    .X(_1807_));
 sky130_fd_sc_hd__inv_2 _1915_ (.A(_1807_),
    .Y(_1808_));
 sky130_fd_sc_hd__or3b_1 _1916_ (.A(net83),
    .B(net84),
    .C_N(\S8x305.I[8] ),
    .X(_1809_));
 sky130_fd_sc_hd__o21ai_1 _1917_ (.A1(net82),
    .A2(net84),
    .B1(net407),
    .Y(_1810_));
 sky130_fd_sc_hd__and2_1 _1918_ (.A(_1809_),
    .B(_1810_),
    .X(_1811_));
 sky130_fd_sc_hd__nand2_1 _1919_ (.A(_1809_),
    .B(_1810_),
    .Y(_1812_));
 sky130_fd_sc_hd__or3_2 _1920_ (.A(_1794_),
    .B(_1797_),
    .C(net71),
    .X(_1813_));
 sky130_fd_sc_hd__o21a_2 _1921_ (.A1(net63),
    .A2(_1807_),
    .B1(_1813_),
    .X(_1814_));
 sky130_fd_sc_hd__o21ai_2 _1922_ (.A1(net63),
    .A2(_1807_),
    .B1(_1813_),
    .Y(_1815_));
 sky130_fd_sc_hd__o2111a_4 _1923_ (.A1(net63),
    .A2(_1807_),
    .B1(_1813_),
    .C1(_1803_),
    .D1(_1805_),
    .X(_1816_));
 sky130_fd_sc_hd__nand2_1 _1924_ (.A(_1806_),
    .B(_1814_),
    .Y(_1817_));
 sky130_fd_sc_hd__or3_2 _1925_ (.A(net82),
    .B(net84),
    .C(net425),
    .X(_1818_));
 sky130_fd_sc_hd__o21ai_4 _1926_ (.A1(\S8x305.i_latch[4] ),
    .A2(_1783_),
    .B1(_1818_),
    .Y(_1819_));
 sky130_fd_sc_hd__o21a_4 _1927_ (.A1(net757),
    .A2(_1783_),
    .B1(_1818_),
    .X(_1820_));
 sky130_fd_sc_hd__a21oi_4 _1928_ (.A1(net853),
    .A2(_1796_),
    .B1(_1819_),
    .Y(_1821_));
 sky130_fd_sc_hd__nor2_1 _1929_ (.A(_1753_),
    .B(_1784_),
    .Y(_1822_));
 sky130_fd_sc_hd__a21oi_2 _1930_ (.A1(net449),
    .A2(_1784_),
    .B1(_1822_),
    .Y(_1823_));
 sky130_fd_sc_hd__mux2_4 _1931_ (.A0(net804),
    .A1(net449),
    .S(_1784_),
    .X(_1824_));
 sky130_fd_sc_hd__a21oi_4 _1932_ (.A1(net63),
    .A2(net66),
    .B1(_1821_),
    .Y(_1825_));
 sky130_fd_sc_hd__mux2_8 _1933_ (.A0(net732),
    .A1(net378),
    .S(_1784_),
    .X(_1826_));
 sky130_fd_sc_hd__or2_2 _1934_ (.A(net676),
    .B(_1784_),
    .X(_1827_));
 sky130_fd_sc_hd__o21ai_4 _1935_ (.A1(net713),
    .A2(_1783_),
    .B1(_1827_),
    .Y(_1828_));
 sky130_fd_sc_hd__o21a_4 _1936_ (.A1(\S8x305.i_latch[10] ),
    .A2(_1783_),
    .B1(_1827_),
    .X(_1829_));
 sky130_fd_sc_hd__mux2_4 _1937_ (.A0(_1826_),
    .A1(net60),
    .S(net63),
    .X(_1830_));
 sky130_fd_sc_hd__nor2_2 _1938_ (.A(_1788_),
    .B(_1796_),
    .Y(_1831_));
 sky130_fd_sc_hd__nand2_1 _1939_ (.A(_1787_),
    .B(_1797_),
    .Y(_1832_));
 sky130_fd_sc_hd__and3_2 _1940_ (.A(_1787_),
    .B(_1791_),
    .C(_1797_),
    .X(_1833_));
 sky130_fd_sc_hd__nand2_1 _1941_ (.A(_1791_),
    .B(_1831_),
    .Y(_1834_));
 sky130_fd_sc_hd__or2_1 _1942_ (.A(net63),
    .B(_1833_),
    .X(_1835_));
 sky130_fd_sc_hd__and4_4 _1943_ (.A(_1816_),
    .B(_1825_),
    .C(_1830_),
    .D(_1835_),
    .X(_1836_));
 sky130_fd_sc_hd__and2_1 _1944_ (.A(net82),
    .B(_1836_),
    .X(net33));
 sky130_fd_sc_hd__nand2_4 _1945_ (.A(_1787_),
    .B(_1796_),
    .Y(_1837_));
 sky130_fd_sc_hd__a21bo_1 _1946_ (.A1(_1792_),
    .A2(_1837_),
    .B1_N(net82),
    .X(_0430_));
 sky130_fd_sc_hd__inv_2 _1947_ (.A(_0430_),
    .Y(_0431_));
 sky130_fd_sc_hd__and3_1 _1948_ (.A(_1816_),
    .B(_1825_),
    .C(_0431_),
    .X(_0432_));
 sky130_fd_sc_hd__or2_2 _1949_ (.A(net776),
    .B(_1784_),
    .X(_0433_));
 sky130_fd_sc_hd__o21a_2 _1950_ (.A1(net684),
    .A2(_1783_),
    .B1(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__o21ai_4 _1951_ (.A1(net684),
    .A2(_1783_),
    .B1(_0433_),
    .Y(_0435_));
 sky130_fd_sc_hd__mux2_8 _1952_ (.A0(net794),
    .A1(net433),
    .S(_1784_),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_4 _1953_ (.A0(_0434_),
    .A1(_0436_),
    .S(_1799_),
    .X(_0437_));
 sky130_fd_sc_hd__inv_2 _1954_ (.A(_0437_),
    .Y(_0438_));
 sky130_fd_sc_hd__o31a_1 _1955_ (.A1(\S8x305.I[12] ),
    .A2(_1784_),
    .A3(_1834_),
    .B1(_0430_),
    .X(_0439_));
 sky130_fd_sc_hd__or2_1 _1956_ (.A(_1825_),
    .B(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__inv_2 _1957_ (.A(_0440_),
    .Y(_0441_));
 sky130_fd_sc_hd__a2bb2o_1 _1958_ (.A1_N(_1753_),
    .A2_N(_0433_),
    .B1(_0438_),
    .B2(_0441_),
    .X(_0442_));
 sky130_fd_sc_hd__and4_2 _1959_ (.A(net63),
    .B(net72),
    .C(_1828_),
    .D(_0434_),
    .X(_0443_));
 sky130_fd_sc_hd__and2_2 _1960_ (.A(_1806_),
    .B(_1815_),
    .X(_0444_));
 sky130_fd_sc_hd__nand2_1 _1961_ (.A(_1806_),
    .B(_1815_),
    .Y(_0445_));
 sky130_fd_sc_hd__and4b_1 _1962_ (.A_N(_1830_),
    .B(_0437_),
    .C(_0444_),
    .D(_1825_),
    .X(_0446_));
 sky130_fd_sc_hd__a31o_1 _1963_ (.A1(net82),
    .A2(_0443_),
    .A3(_0446_),
    .B1(_0442_),
    .X(_0447_));
 sky130_fd_sc_hd__a31o_4 _1964_ (.A1(_1830_),
    .A2(_0432_),
    .A3(_0438_),
    .B1(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__inv_2 _1965_ (.A(_0448_),
    .Y(net32));
 sky130_fd_sc_hd__and3_1 _1966_ (.A(net82),
    .B(\S8x305.i_latch[8] ),
    .C(_0443_),
    .X(_0449_));
 sky130_fd_sc_hd__a221o_1 _1967_ (.A1(\S8x305.I[11] ),
    .A2(_1822_),
    .B1(_0437_),
    .B2(_0441_),
    .C1(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__a31oi_4 _1968_ (.A1(_1830_),
    .A2(_0432_),
    .A3(_0437_),
    .B1(_0450_),
    .Y(net31));
 sky130_fd_sc_hd__a32o_1 _1969_ (.A1(net853),
    .A2(_1796_),
    .A3(net66),
    .B1(_1820_),
    .B2(_1791_),
    .X(_0451_));
 sky130_fd_sc_hd__a41o_1 _1970_ (.A1(net63),
    .A2(net72),
    .A3(_1828_),
    .A4(_0434_),
    .B1(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__and2_2 _1971_ (.A(net82),
    .B(_0452_),
    .X(net34));
 sky130_fd_sc_hd__and2b_1 _1972_ (.A_N(ROM_spi_mode),
    .B(ROM_OEB),
    .X(net28));
 sky130_fd_sc_hd__or2_1 _1973_ (.A(ROM_spi_mode),
    .B(ROM_OEB),
    .X(net26));
 sky130_fd_sc_hd__nor2_1 _1974_ (.A(_1836_),
    .B(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__a41o_2 _1975_ (.A1(_1816_),
    .A2(_1825_),
    .A3(_1830_),
    .A4(_1835_),
    .B1(_0452_),
    .X(_0454_));
 sky130_fd_sc_hd__nand2_2 _1976_ (.A(net82),
    .B(_0454_),
    .Y(net24));
 sky130_fd_sc_hd__nor2_2 _1977_ (.A(_1799_),
    .B(_0453_),
    .Y(_0455_));
 sky130_fd_sc_hd__nand2_4 _1978_ (.A(net63),
    .B(_0454_),
    .Y(_0456_));
 sky130_fd_sc_hd__or2_1 _1979_ (.A(net427),
    .B(_1784_),
    .X(_0457_));
 sky130_fd_sc_hd__o21ai_4 _1980_ (.A1(net710),
    .A2(_1783_),
    .B1(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__o21a_2 _1981_ (.A1(net710),
    .A2(_1783_),
    .B1(_0457_),
    .X(_0459_));
 sky130_fd_sc_hd__nor2_2 _1982_ (.A(net66),
    .B(_0458_),
    .Y(_0460_));
 sky130_fd_sc_hd__and2b_4 _1983_ (.A_N(net83),
    .B(net84),
    .X(_0461_));
 sky130_fd_sc_hd__nand2b_4 _1984_ (.A_N(net83),
    .B(net84),
    .Y(_0462_));
 sky130_fd_sc_hd__and3_4 _1985_ (.A(_1791_),
    .B(_1820_),
    .C(_0461_),
    .X(_0463_));
 sky130_fd_sc_hd__or3_4 _1986_ (.A(_1792_),
    .B(_1819_),
    .C(_0462_),
    .X(_0464_));
 sky130_fd_sc_hd__nor2_1 _1987_ (.A(_1794_),
    .B(_1796_),
    .Y(_0465_));
 sky130_fd_sc_hd__nand2_1 _1988_ (.A(net853),
    .B(_1797_),
    .Y(_0466_));
 sky130_fd_sc_hd__or2_1 _1989_ (.A(net405),
    .B(_1784_),
    .X(_0467_));
 sky130_fd_sc_hd__o21ai_2 _1990_ (.A1(net701),
    .A2(_1783_),
    .B1(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__o21a_2 _1991_ (.A1(net451),
    .A2(_1783_),
    .B1(_0467_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _1992_ (.A0(_0468_),
    .A1(_1804_),
    .S(_1821_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _1993_ (.A0(net73),
    .A1(_0470_),
    .S(net61),
    .X(_0471_));
 sky130_fd_sc_hd__o22a_4 _1994_ (.A1(net62),
    .A2(net59),
    .B1(_0471_),
    .B2(net853),
    .X(_0472_));
 sky130_fd_sc_hd__inv_2 _1995_ (.A(_0472_),
    .Y(_0473_));
 sky130_fd_sc_hd__mux2_4 _1996_ (.A0(net421),
    .A1(net386),
    .S(_1784_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _1997_ (.A0(_0474_),
    .A1(_1808_),
    .S(_1821_),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _1998_ (.A0(_1811_),
    .A1(_0475_),
    .S(net61),
    .X(_0476_));
 sky130_fd_sc_hd__o2bb2a_4 _1999_ (.A1_N(_1794_),
    .A2_N(_0476_),
    .B1(net59),
    .B2(_1811_),
    .X(_0477_));
 sky130_fd_sc_hd__a22o_2 _2000_ (.A1(net71),
    .A2(_0465_),
    .B1(_0476_),
    .B2(_1794_),
    .X(_0478_));
 sky130_fd_sc_hd__and2_1 _2001_ (.A(_0472_),
    .B(_0477_),
    .X(_0479_));
 sky130_fd_sc_hd__nand2_1 _2002_ (.A(_0472_),
    .B(_0477_),
    .Y(_0480_));
 sky130_fd_sc_hd__nor2_1 _2003_ (.A(_0472_),
    .B(_0477_),
    .Y(_0481_));
 sky130_fd_sc_hd__nor2_1 _2004_ (.A(_0479_),
    .B(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__or2_2 _2005_ (.A(_0479_),
    .B(_0481_),
    .X(_0483_));
 sky130_fd_sc_hd__nor2_8 _2006_ (.A(_1821_),
    .B(net65),
    .Y(_0484_));
 sky130_fd_sc_hd__or2_2 _2007_ (.A(_1821_),
    .B(_1824_),
    .X(_0485_));
 sky130_fd_sc_hd__and3b_2 _2008_ (.A_N(net84),
    .B(net599),
    .C(net83),
    .X(_0486_));
 sky130_fd_sc_hd__or3b_4 _2009_ (.A(net488),
    .B(_1740_),
    .C_N(net83),
    .X(_0487_));
 sky130_fd_sc_hd__and3_2 _2010_ (.A(net113),
    .B(_1791_),
    .C(_0486_),
    .X(_0488_));
 sky130_fd_sc_hd__a31o_2 _2011_ (.A1(_1799_),
    .A2(_0454_),
    .A3(_0461_),
    .B1(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__nand2_4 _2012_ (.A(_0484_),
    .B(_0489_),
    .Y(_0490_));
 sky130_fd_sc_hd__mux2_1 _2013_ (.A0(\S8x305.regs[8][1] ),
    .A1(\S8x305.regs[9][1] ),
    .S(net67),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_1 _2014_ (.A0(\S8x305.regs[10][1] ),
    .A1(\S8x305.regs[11][1] ),
    .S(net67),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_1 _2015_ (.A0(_0491_),
    .A1(_0492_),
    .S(net73),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _2016_ (.A0(\S8x305.regs[14][1] ),
    .A1(\S8x305.regs[15][1] ),
    .S(net67),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _2017_ (.A0(\S8x305.regs[12][1] ),
    .A1(\S8x305.regs[13][1] ),
    .S(net67),
    .X(_0495_));
 sky130_fd_sc_hd__mux2_1 _2018_ (.A0(_0494_),
    .A1(_0495_),
    .S(net62),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_1 _2019_ (.A0(_0493_),
    .A1(_0496_),
    .S(net60),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _2020_ (.A0(\S8x305.ALU_in1[1] ),
    .A1(\S8x305.regs[1][1] ),
    .S(net69),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _2021_ (.A0(\S8x305.regs[2][1] ),
    .A1(\S8x305.regs[3][1] ),
    .S(net70),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _2022_ (.A0(_0498_),
    .A1(_0499_),
    .S(net72),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _2023_ (.A0(\S8x305.regs[6][1] ),
    .A1(\S8x305.regs[7][1] ),
    .S(net69),
    .X(_0501_));
 sky130_fd_sc_hd__or2_1 _2024_ (.A(net62),
    .B(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _2025_ (.A0(\S8x305.regs[4][1] ),
    .A1(\S8x305.regs[5][1] ),
    .S(net69),
    .X(_0503_));
 sky130_fd_sc_hd__o21a_1 _2026_ (.A1(net72),
    .A2(_0503_),
    .B1(net60),
    .X(_0504_));
 sky130_fd_sc_hd__a22o_1 _2027_ (.A1(_1828_),
    .A2(_0500_),
    .B1(_0502_),
    .B2(_0504_),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_2 _2028_ (.A0(_0497_),
    .A1(_0505_),
    .S(_0435_),
    .X(_0506_));
 sky130_fd_sc_hd__a21oi_1 _2029_ (.A1(_0484_),
    .A2(_0489_),
    .B1(net75),
    .Y(_0507_));
 sky130_fd_sc_hd__and3_1 _2030_ (.A(_0484_),
    .B(_0489_),
    .C(_0506_),
    .X(_0508_));
 sky130_fd_sc_hd__or3_1 _2031_ (.A(_0478_),
    .B(_0507_),
    .C(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _2032_ (.A0(\S8x305.regs[8][0] ),
    .A1(\S8x305.regs[9][0] ),
    .S(net68),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _2033_ (.A0(\S8x305.regs[10][0] ),
    .A1(\S8x305.regs[11][0] ),
    .S(net68),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _2034_ (.A0(_0510_),
    .A1(_0511_),
    .S(net73),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _2035_ (.A0(\S8x305.regs[14][0] ),
    .A1(\S8x305.regs[15][0] ),
    .S(net68),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _2036_ (.A0(\S8x305.regs[12][0] ),
    .A1(\S8x305.regs[13][0] ),
    .S(net68),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _2037_ (.A0(_0513_),
    .A1(_0514_),
    .S(net62),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _2038_ (.A0(_0512_),
    .A1(_0515_),
    .S(net60),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _2039_ (.A0(\S8x305.ALU_in1[0] ),
    .A1(\S8x305.regs[1][0] ),
    .S(net69),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_1 _2040_ (.A0(\S8x305.regs[2][0] ),
    .A1(\S8x305.regs[3][0] ),
    .S(net70),
    .X(_0518_));
 sky130_fd_sc_hd__mux2_1 _2041_ (.A0(_0517_),
    .A1(_0518_),
    .S(net72),
    .X(_0519_));
 sky130_fd_sc_hd__mux2_1 _2042_ (.A0(\S8x305.regs[6][0] ),
    .A1(\S8x305.regs[7][0] ),
    .S(net68),
    .X(_0520_));
 sky130_fd_sc_hd__mux2_1 _2043_ (.A0(\S8x305.regs[4][0] ),
    .A1(\S8x305.regs[5][0] ),
    .S(net69),
    .X(_0521_));
 sky130_fd_sc_hd__o21a_1 _2044_ (.A1(net62),
    .A2(_0520_),
    .B1(net60),
    .X(_0522_));
 sky130_fd_sc_hd__o21ai_1 _2045_ (.A1(net73),
    .A2(_0521_),
    .B1(_0522_),
    .Y(_0523_));
 sky130_fd_sc_hd__a21oi_1 _2046_ (.A1(_1828_),
    .A2(_0519_),
    .B1(_0434_),
    .Y(_0524_));
 sky130_fd_sc_hd__o2bb2a_2 _2047_ (.A1_N(_0523_),
    .A2_N(_0524_),
    .B1(_0435_),
    .B2(_0516_),
    .X(_0525_));
 sky130_fd_sc_hd__mux2_2 _2048_ (.A0(_0525_),
    .A1(\S8x305.iv_latch[0] ),
    .S(_0490_),
    .X(_0526_));
 sky130_fd_sc_hd__o21a_1 _2049_ (.A1(_0477_),
    .A2(_0526_),
    .B1(_0509_),
    .X(_0527_));
 sky130_fd_sc_hd__mux2_1 _2050_ (.A0(\S8x305.regs[8][3] ),
    .A1(\S8x305.regs[9][3] ),
    .S(net67),
    .X(_0528_));
 sky130_fd_sc_hd__mux2_1 _2051_ (.A0(\S8x305.regs[10][3] ),
    .A1(\S8x305.regs[11][3] ),
    .S(net67),
    .X(_0529_));
 sky130_fd_sc_hd__mux2_1 _2052_ (.A0(_0528_),
    .A1(_0529_),
    .S(net73),
    .X(_0530_));
 sky130_fd_sc_hd__mux2_1 _2053_ (.A0(\S8x305.regs[14][3] ),
    .A1(\S8x305.regs[15][3] ),
    .S(net68),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_1 _2054_ (.A0(\S8x305.regs[12][3] ),
    .A1(\S8x305.regs[13][3] ),
    .S(net68),
    .X(_0532_));
 sky130_fd_sc_hd__mux2_1 _2055_ (.A0(_0531_),
    .A1(_0532_),
    .S(net62),
    .X(_0533_));
 sky130_fd_sc_hd__mux2_1 _2056_ (.A0(_0530_),
    .A1(_0533_),
    .S(net60),
    .X(_0534_));
 sky130_fd_sc_hd__mux2_1 _2057_ (.A0(\S8x305.ALU_in1[3] ),
    .A1(\S8x305.regs[1][3] ),
    .S(net70),
    .X(_0535_));
 sky130_fd_sc_hd__mux2_1 _2058_ (.A0(\S8x305.regs[2][3] ),
    .A1(\S8x305.regs[3][3] ),
    .S(net70),
    .X(_0536_));
 sky130_fd_sc_hd__mux2_1 _2059_ (.A0(_0535_),
    .A1(_0536_),
    .S(net72),
    .X(_0537_));
 sky130_fd_sc_hd__mux2_1 _2060_ (.A0(\S8x305.regs[6][3] ),
    .A1(\S8x305.regs[7][3] ),
    .S(net68),
    .X(_0538_));
 sky130_fd_sc_hd__or2_1 _2061_ (.A(net62),
    .B(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__mux2_1 _2062_ (.A0(\S8x305.regs[4][3] ),
    .A1(\S8x305.regs[5][3] ),
    .S(net69),
    .X(_0540_));
 sky130_fd_sc_hd__o21a_1 _2063_ (.A1(net72),
    .A2(_0540_),
    .B1(net60),
    .X(_0541_));
 sky130_fd_sc_hd__a22o_1 _2064_ (.A1(_1828_),
    .A2(_0537_),
    .B1(_0539_),
    .B2(_0541_),
    .X(_0542_));
 sky130_fd_sc_hd__mux2_2 _2065_ (.A0(_0534_),
    .A1(_0542_),
    .S(_0435_),
    .X(_0543_));
 sky130_fd_sc_hd__and3_1 _2066_ (.A(_0484_),
    .B(_0489_),
    .C(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__a211o_1 _2067_ (.A1(\S8x305.iv_latch[3] ),
    .A2(_0490_),
    .B1(_0544_),
    .C1(_0478_),
    .X(_0545_));
 sky130_fd_sc_hd__mux2_1 _2068_ (.A0(\S8x305.regs[8][2] ),
    .A1(\S8x305.regs[9][2] ),
    .S(net71),
    .X(_0546_));
 sky130_fd_sc_hd__mux2_1 _2069_ (.A0(\S8x305.regs[10][2] ),
    .A1(\S8x305.regs[11][2] ),
    .S(net67),
    .X(_0547_));
 sky130_fd_sc_hd__mux2_1 _2070_ (.A0(_0546_),
    .A1(_0547_),
    .S(net73),
    .X(_0548_));
 sky130_fd_sc_hd__mux2_1 _2071_ (.A0(\S8x305.regs[14][2] ),
    .A1(\S8x305.regs[15][2] ),
    .S(net68),
    .X(_0549_));
 sky130_fd_sc_hd__mux2_1 _2072_ (.A0(\S8x305.regs[12][2] ),
    .A1(\S8x305.regs[13][2] ),
    .S(net67),
    .X(_0550_));
 sky130_fd_sc_hd__mux2_1 _2073_ (.A0(_0549_),
    .A1(_0550_),
    .S(net62),
    .X(_0551_));
 sky130_fd_sc_hd__mux2_1 _2074_ (.A0(_0548_),
    .A1(_0551_),
    .S(net60),
    .X(_0552_));
 sky130_fd_sc_hd__mux2_1 _2075_ (.A0(\S8x305.ALU_in1[2] ),
    .A1(\S8x305.regs[1][2] ),
    .S(net69),
    .X(_0553_));
 sky130_fd_sc_hd__mux2_1 _2076_ (.A0(\S8x305.regs[2][2] ),
    .A1(\S8x305.regs[3][2] ),
    .S(net70),
    .X(_0554_));
 sky130_fd_sc_hd__mux2_1 _2077_ (.A0(_0553_),
    .A1(_0554_),
    .S(net72),
    .X(_0555_));
 sky130_fd_sc_hd__mux2_1 _2078_ (.A0(\S8x305.regs[6][2] ),
    .A1(\S8x305.regs[7][2] ),
    .S(net68),
    .X(_0556_));
 sky130_fd_sc_hd__or2_1 _2079_ (.A(net62),
    .B(_0556_),
    .X(_0557_));
 sky130_fd_sc_hd__mux2_1 _2080_ (.A0(\S8x305.regs[4][2] ),
    .A1(\S8x305.regs[5][2] ),
    .S(net69),
    .X(_0558_));
 sky130_fd_sc_hd__o21a_1 _2081_ (.A1(net72),
    .A2(_0558_),
    .B1(net60),
    .X(_0559_));
 sky130_fd_sc_hd__a22o_1 _2082_ (.A1(_1828_),
    .A2(_0555_),
    .B1(_0557_),
    .B2(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__mux2_2 _2083_ (.A0(_0552_),
    .A1(_0560_),
    .S(_0435_),
    .X(_0561_));
 sky130_fd_sc_hd__and3_1 _2084_ (.A(_0484_),
    .B(_0489_),
    .C(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__a211o_1 _2085_ (.A1(\S8x305.iv_latch[2] ),
    .A2(_0490_),
    .B1(_0562_),
    .C1(_0477_),
    .X(_0563_));
 sky130_fd_sc_hd__and3_1 _2086_ (.A(_0483_),
    .B(_0545_),
    .C(_0563_),
    .X(_0564_));
 sky130_fd_sc_hd__a21o_1 _2087_ (.A1(_0482_),
    .A2(_0527_),
    .B1(_0564_),
    .X(_0565_));
 sky130_fd_sc_hd__mux2_1 _2088_ (.A0(_0458_),
    .A1(_1826_),
    .S(_1821_),
    .X(_0566_));
 sky130_fd_sc_hd__mux2_1 _2089_ (.A0(net60),
    .A1(_0566_),
    .S(net61),
    .X(_0567_));
 sky130_fd_sc_hd__o22a_4 _2090_ (.A1(_1828_),
    .A2(_0466_),
    .B1(_0567_),
    .B2(net853),
    .X(_0568_));
 sky130_fd_sc_hd__a2bb2o_2 _2091_ (.A1_N(net853),
    .A2_N(_0567_),
    .B1(_0465_),
    .B2(net60),
    .X(_0569_));
 sky130_fd_sc_hd__nor2_1 _2092_ (.A(_0480_),
    .B(_0569_),
    .Y(_0570_));
 sky130_fd_sc_hd__nor2_1 _2093_ (.A(_0479_),
    .B(_0568_),
    .Y(_0571_));
 sky130_fd_sc_hd__nor2_1 _2094_ (.A(_0570_),
    .B(_0571_),
    .Y(_0572_));
 sky130_fd_sc_hd__mux2_1 _2095_ (.A0(\S8x305.regs[8][7] ),
    .A1(\S8x305.regs[9][7] ),
    .S(net68),
    .X(_0573_));
 sky130_fd_sc_hd__mux2_1 _2096_ (.A0(\S8x305.regs[10][7] ),
    .A1(\S8x305.regs[11][7] ),
    .S(net68),
    .X(_0574_));
 sky130_fd_sc_hd__mux2_1 _2097_ (.A0(_0573_),
    .A1(_0574_),
    .S(net73),
    .X(_0575_));
 sky130_fd_sc_hd__mux2_1 _2098_ (.A0(\S8x305.regs[14][7] ),
    .A1(\S8x305.regs[15][7] ),
    .S(net68),
    .X(_0576_));
 sky130_fd_sc_hd__mux2_1 _2099_ (.A0(\S8x305.regs[12][7] ),
    .A1(\S8x305.regs[13][7] ),
    .S(net68),
    .X(_0577_));
 sky130_fd_sc_hd__mux2_1 _2100_ (.A0(_0576_),
    .A1(_0577_),
    .S(net62),
    .X(_0578_));
 sky130_fd_sc_hd__mux2_1 _2101_ (.A0(_0575_),
    .A1(_0578_),
    .S(net60),
    .X(_0579_));
 sky130_fd_sc_hd__mux2_1 _2102_ (.A0(\S8x305.ALU_in1[7] ),
    .A1(\S8x305.regs[1][7] ),
    .S(net70),
    .X(_0580_));
 sky130_fd_sc_hd__mux2_1 _2103_ (.A0(\S8x305.regs[2][7] ),
    .A1(\S8x305.regs[3][7] ),
    .S(net70),
    .X(_0581_));
 sky130_fd_sc_hd__mux2_1 _2104_ (.A0(_0580_),
    .A1(_0581_),
    .S(net72),
    .X(_0582_));
 sky130_fd_sc_hd__mux2_1 _2105_ (.A0(\S8x305.regs[6][7] ),
    .A1(\S8x305.regs[7][7] ),
    .S(net69),
    .X(_0583_));
 sky130_fd_sc_hd__or2_1 _2106_ (.A(net62),
    .B(_0583_),
    .X(_0584_));
 sky130_fd_sc_hd__mux2_1 _2107_ (.A0(\S8x305.regs[4][7] ),
    .A1(\S8x305.regs[5][7] ),
    .S(net69),
    .X(_0585_));
 sky130_fd_sc_hd__o21a_1 _2108_ (.A1(net72),
    .A2(_0585_),
    .B1(net60),
    .X(_0586_));
 sky130_fd_sc_hd__a22o_1 _2109_ (.A1(_1828_),
    .A2(_0582_),
    .B1(_0584_),
    .B2(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__mux2_2 _2110_ (.A0(_0579_),
    .A1(_0587_),
    .S(_0435_),
    .X(_0588_));
 sky130_fd_sc_hd__and3_1 _2111_ (.A(_0484_),
    .B(_0489_),
    .C(_0588_),
    .X(_0589_));
 sky130_fd_sc_hd__a21o_1 _2112_ (.A1(\S8x305.iv_latch[7] ),
    .A2(_0490_),
    .B1(_0589_),
    .X(_0590_));
 sky130_fd_sc_hd__mux2_1 _2113_ (.A0(\S8x305.regs[8][5] ),
    .A1(\S8x305.regs[9][5] ),
    .S(net71),
    .X(_0591_));
 sky130_fd_sc_hd__mux2_1 _2114_ (.A0(\S8x305.regs[10][5] ),
    .A1(\S8x305.regs[11][5] ),
    .S(net67),
    .X(_0592_));
 sky130_fd_sc_hd__mux2_1 _2115_ (.A0(_0591_),
    .A1(_0592_),
    .S(net73),
    .X(_0593_));
 sky130_fd_sc_hd__mux2_1 _2116_ (.A0(\S8x305.regs[14][5] ),
    .A1(\S8x305.regs[15][5] ),
    .S(net67),
    .X(_0594_));
 sky130_fd_sc_hd__mux2_1 _2117_ (.A0(\S8x305.regs[12][5] ),
    .A1(\S8x305.regs[13][5] ),
    .S(net71),
    .X(_0595_));
 sky130_fd_sc_hd__mux2_1 _2118_ (.A0(_0594_),
    .A1(_0595_),
    .S(net62),
    .X(_0596_));
 sky130_fd_sc_hd__mux2_1 _2119_ (.A0(_0593_),
    .A1(_0596_),
    .S(net60),
    .X(_0597_));
 sky130_fd_sc_hd__mux2_1 _2120_ (.A0(\S8x305.ALU_in1[5] ),
    .A1(\S8x305.regs[1][5] ),
    .S(net70),
    .X(_0598_));
 sky130_fd_sc_hd__mux2_1 _2121_ (.A0(\S8x305.regs[2][5] ),
    .A1(\S8x305.regs[3][5] ),
    .S(net70),
    .X(_0599_));
 sky130_fd_sc_hd__mux2_1 _2122_ (.A0(_0598_),
    .A1(_0599_),
    .S(net73),
    .X(_0600_));
 sky130_fd_sc_hd__mux2_1 _2123_ (.A0(\S8x305.regs[6][5] ),
    .A1(\S8x305.regs[7][5] ),
    .S(net69),
    .X(_0601_));
 sky130_fd_sc_hd__or2_1 _2124_ (.A(net62),
    .B(_0601_),
    .X(_0602_));
 sky130_fd_sc_hd__mux2_1 _2125_ (.A0(\S8x305.regs[4][5] ),
    .A1(\S8x305.regs[5][5] ),
    .S(net69),
    .X(_0603_));
 sky130_fd_sc_hd__o21a_1 _2126_ (.A1(net73),
    .A2(_0603_),
    .B1(_1829_),
    .X(_0604_));
 sky130_fd_sc_hd__a22o_1 _2127_ (.A1(_1828_),
    .A2(_0600_),
    .B1(_0602_),
    .B2(_0604_),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_2 _2128_ (.A0(_0597_),
    .A1(_0605_),
    .S(_0435_),
    .X(_0606_));
 sky130_fd_sc_hd__and3_1 _2129_ (.A(_0484_),
    .B(_0489_),
    .C(_0606_),
    .X(_0607_));
 sky130_fd_sc_hd__a211o_1 _2130_ (.A1(\S8x305.iv_latch[5] ),
    .A2(_0490_),
    .B1(_0607_),
    .C1(_0478_),
    .X(_0608_));
 sky130_fd_sc_hd__mux2_1 _2131_ (.A0(\S8x305.regs[8][4] ),
    .A1(\S8x305.regs[9][4] ),
    .S(net71),
    .X(_0609_));
 sky130_fd_sc_hd__mux2_1 _2132_ (.A0(\S8x305.regs[10][4] ),
    .A1(\S8x305.regs[11][4] ),
    .S(net67),
    .X(_0610_));
 sky130_fd_sc_hd__mux2_1 _2133_ (.A0(_0609_),
    .A1(_0610_),
    .S(net73),
    .X(_0611_));
 sky130_fd_sc_hd__mux2_1 _2134_ (.A0(\S8x305.regs[14][4] ),
    .A1(\S8x305.regs[15][4] ),
    .S(net67),
    .X(_0612_));
 sky130_fd_sc_hd__mux2_1 _2135_ (.A0(\S8x305.regs[12][4] ),
    .A1(\S8x305.regs[13][4] ),
    .S(net67),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_1 _2136_ (.A0(_0612_),
    .A1(_0613_),
    .S(net62),
    .X(_0614_));
 sky130_fd_sc_hd__mux2_1 _2137_ (.A0(_0611_),
    .A1(_0614_),
    .S(_1829_),
    .X(_0615_));
 sky130_fd_sc_hd__mux2_1 _2138_ (.A0(\S8x305.ALU_in1[4] ),
    .A1(\S8x305.regs[1][4] ),
    .S(net70),
    .X(_0616_));
 sky130_fd_sc_hd__mux2_1 _2139_ (.A0(\S8x305.regs[2][4] ),
    .A1(\S8x305.regs[3][4] ),
    .S(net70),
    .X(_0617_));
 sky130_fd_sc_hd__mux2_1 _2140_ (.A0(_0616_),
    .A1(_0617_),
    .S(net72),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_1 _2141_ (.A0(\S8x305.regs[6][4] ),
    .A1(\S8x305.regs[7][4] ),
    .S(net69),
    .X(_0619_));
 sky130_fd_sc_hd__or2_1 _2142_ (.A(net62),
    .B(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__mux2_1 _2143_ (.A0(\S8x305.regs[4][4] ),
    .A1(\S8x305.regs[5][4] ),
    .S(net69),
    .X(_0621_));
 sky130_fd_sc_hd__o21a_1 _2144_ (.A1(net72),
    .A2(_0621_),
    .B1(_1829_),
    .X(_0622_));
 sky130_fd_sc_hd__a22o_1 _2145_ (.A1(_1828_),
    .A2(_0618_),
    .B1(_0620_),
    .B2(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__mux2_2 _2146_ (.A0(_0615_),
    .A1(_0623_),
    .S(_0435_),
    .X(_0624_));
 sky130_fd_sc_hd__and3_1 _2147_ (.A(_0484_),
    .B(_0489_),
    .C(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__a211o_1 _2148_ (.A1(\S8x305.iv_latch[4] ),
    .A2(_0490_),
    .B1(_0625_),
    .C1(_0477_),
    .X(_0626_));
 sky130_fd_sc_hd__mux2_1 _2149_ (.A0(\S8x305.regs[8][6] ),
    .A1(\S8x305.regs[9][6] ),
    .S(net67),
    .X(_0627_));
 sky130_fd_sc_hd__mux2_1 _2150_ (.A0(\S8x305.regs[10][6] ),
    .A1(\S8x305.regs[11][6] ),
    .S(net67),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_1 _2151_ (.A0(_0627_),
    .A1(_0628_),
    .S(net73),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_1 _2152_ (.A0(\S8x305.regs[14][6] ),
    .A1(\S8x305.regs[15][6] ),
    .S(net67),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_1 _2153_ (.A0(\S8x305.regs[12][6] ),
    .A1(\S8x305.regs[13][6] ),
    .S(net71),
    .X(_0631_));
 sky130_fd_sc_hd__mux2_1 _2154_ (.A0(_0630_),
    .A1(_0631_),
    .S(_1802_),
    .X(_0632_));
 sky130_fd_sc_hd__mux2_1 _2155_ (.A0(_0629_),
    .A1(_0632_),
    .S(_1829_),
    .X(_0633_));
 sky130_fd_sc_hd__mux2_1 _2156_ (.A0(\S8x305.ALU_in1[6] ),
    .A1(\S8x305.regs[1][6] ),
    .S(net69),
    .X(_0634_));
 sky130_fd_sc_hd__mux2_1 _2157_ (.A0(\S8x305.regs[2][6] ),
    .A1(\S8x305.regs[3][6] ),
    .S(net70),
    .X(_0635_));
 sky130_fd_sc_hd__mux2_1 _2158_ (.A0(_0634_),
    .A1(_0635_),
    .S(net72),
    .X(_0636_));
 sky130_fd_sc_hd__mux2_1 _2159_ (.A0(\S8x305.regs[6][6] ),
    .A1(\S8x305.regs[7][6] ),
    .S(net68),
    .X(_0637_));
 sky130_fd_sc_hd__or2_1 _2160_ (.A(_1802_),
    .B(_0637_),
    .X(_0638_));
 sky130_fd_sc_hd__mux2_1 _2161_ (.A0(\S8x305.regs[4][6] ),
    .A1(\S8x305.regs[5][6] ),
    .S(net69),
    .X(_0639_));
 sky130_fd_sc_hd__o21a_1 _2162_ (.A1(net72),
    .A2(_0639_),
    .B1(_1829_),
    .X(_0640_));
 sky130_fd_sc_hd__a22o_1 _2163_ (.A1(_1828_),
    .A2(_0636_),
    .B1(_0638_),
    .B2(_0640_),
    .X(_0641_));
 sky130_fd_sc_hd__mux2_2 _2164_ (.A0(_0633_),
    .A1(_0641_),
    .S(_0435_),
    .X(_0642_));
 sky130_fd_sc_hd__and3_1 _2165_ (.A(_0484_),
    .B(_0489_),
    .C(_0642_),
    .X(_0643_));
 sky130_fd_sc_hd__a211o_1 _2166_ (.A1(\S8x305.iv_latch[6] ),
    .A2(_0490_),
    .B1(_0643_),
    .C1(_0477_),
    .X(_0644_));
 sky130_fd_sc_hd__o211a_1 _2167_ (.A1(_0478_),
    .A2(_0590_),
    .B1(_0644_),
    .C1(_0483_),
    .X(_0645_));
 sky130_fd_sc_hd__a31o_1 _2168_ (.A1(_0482_),
    .A2(_0608_),
    .A3(_0626_),
    .B1(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__a22o_1 _2169_ (.A1(_0570_),
    .A2(_0590_),
    .B1(_0646_),
    .B2(_0571_),
    .X(_0647_));
 sky130_fd_sc_hd__a21o_1 _2170_ (.A1(_0565_),
    .A2(_0572_),
    .B1(_0647_),
    .X(_0648_));
 sky130_fd_sc_hd__nor2_1 _2171_ (.A(_0469_),
    .B(_0474_),
    .Y(_0649_));
 sky130_fd_sc_hd__and3_1 _2172_ (.A(_1799_),
    .B(_0458_),
    .C(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__o2bb2a_1 _2173_ (.A1_N(_0648_),
    .A2_N(_0650_),
    .B1(net81),
    .B2(_1799_),
    .X(_0651_));
 sky130_fd_sc_hd__mux2_1 _2174_ (.A0(_0648_),
    .A1(_0588_),
    .S(_1821_),
    .X(_0652_));
 sky130_fd_sc_hd__inv_2 _2175_ (.A(_0652_),
    .Y(_0653_));
 sky130_fd_sc_hd__mux2_1 _2176_ (.A0(_0651_),
    .A1(_0653_),
    .S(net61),
    .X(_0654_));
 sky130_fd_sc_hd__nor2_1 _2177_ (.A(_1773_),
    .B(_0654_),
    .Y(_0655_));
 sky130_fd_sc_hd__nand2_1 _2178_ (.A(_1773_),
    .B(_0654_),
    .Y(_0656_));
 sky130_fd_sc_hd__and2b_1 _2179_ (.A_N(_0655_),
    .B(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__nor2_2 _2180_ (.A(_1787_),
    .B(_1796_),
    .Y(_0658_));
 sky130_fd_sc_hd__nand2_2 _2181_ (.A(_1788_),
    .B(_1797_),
    .Y(_0659_));
 sky130_fd_sc_hd__o221a_1 _2182_ (.A1(_1837_),
    .A2(_0655_),
    .B1(_0657_),
    .B2(_1787_),
    .C1(_0659_),
    .X(_0660_));
 sky130_fd_sc_hd__a211o_1 _2183_ (.A1(\S8x305.iv_latch[4] ),
    .A2(_0490_),
    .B1(_0625_),
    .C1(_0478_),
    .X(_0661_));
 sky130_fd_sc_hd__a211o_1 _2184_ (.A1(\S8x305.iv_latch[3] ),
    .A2(_0490_),
    .B1(_0544_),
    .C1(_0477_),
    .X(_0662_));
 sky130_fd_sc_hd__a21o_1 _2185_ (.A1(_0661_),
    .A2(_0662_),
    .B1(_0483_),
    .X(_0663_));
 sky130_fd_sc_hd__a211o_1 _2186_ (.A1(\S8x305.iv_latch[6] ),
    .A2(_0490_),
    .B1(_0643_),
    .C1(_0478_),
    .X(_0664_));
 sky130_fd_sc_hd__a211o_1 _2187_ (.A1(\S8x305.iv_latch[5] ),
    .A2(_0490_),
    .B1(_0607_),
    .C1(_0477_),
    .X(_0665_));
 sky130_fd_sc_hd__a21o_1 _2188_ (.A1(_0664_),
    .A2(_0665_),
    .B1(_0482_),
    .X(_0666_));
 sky130_fd_sc_hd__and3_1 _2189_ (.A(_0571_),
    .B(_0663_),
    .C(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__a211o_1 _2190_ (.A1(\S8x305.iv_latch[7] ),
    .A2(_0490_),
    .B1(_0589_),
    .C1(_0477_),
    .X(_0668_));
 sky130_fd_sc_hd__and3_1 _2191_ (.A(_0472_),
    .B(_0664_),
    .C(_0668_),
    .X(_0669_));
 sky130_fd_sc_hd__or3_1 _2192_ (.A(_0477_),
    .B(_0507_),
    .C(_0508_),
    .X(_0670_));
 sky130_fd_sc_hd__a211o_1 _2193_ (.A1(\S8x305.iv_latch[2] ),
    .A2(_0490_),
    .B1(_0562_),
    .C1(_0478_),
    .X(_0671_));
 sky130_fd_sc_hd__nor2_1 _2194_ (.A(_0472_),
    .B(_0478_),
    .Y(_0672_));
 sky130_fd_sc_hd__a32o_1 _2195_ (.A1(_0483_),
    .A2(_0670_),
    .A3(_0671_),
    .B1(_0672_),
    .B2(_0526_),
    .X(_0673_));
 sky130_fd_sc_hd__a22o_1 _2196_ (.A1(_0568_),
    .A2(_0669_),
    .B1(_0673_),
    .B2(_0572_),
    .X(_0674_));
 sky130_fd_sc_hd__nor2_1 _2197_ (.A(_0667_),
    .B(_0674_),
    .Y(_0675_));
 sky130_fd_sc_hd__nand2_2 _2198_ (.A(_0469_),
    .B(_0474_),
    .Y(_0676_));
 sky130_fd_sc_hd__nor2_2 _2199_ (.A(_0459_),
    .B(_0649_),
    .Y(_0677_));
 sky130_fd_sc_hd__nor2_1 _2200_ (.A(net63),
    .B(_0677_),
    .Y(_0678_));
 sky130_fd_sc_hd__a211o_1 _2201_ (.A1(_0459_),
    .A2(_0676_),
    .B1(_0677_),
    .C1(net63),
    .X(_0679_));
 sky130_fd_sc_hd__o221a_1 _2202_ (.A1(net80),
    .A2(_1799_),
    .B1(_0675_),
    .B2(_0679_),
    .C1(net65),
    .X(_0680_));
 sky130_fd_sc_hd__o2bb2a_1 _2203_ (.A1_N(_1821_),
    .A2_N(_0642_),
    .B1(_0675_),
    .B2(_0485_),
    .X(_0681_));
 sky130_fd_sc_hd__a21oi_1 _2204_ (.A1(net61),
    .A2(_0681_),
    .B1(_0680_),
    .Y(_0682_));
 sky130_fd_sc_hd__and2_1 _2205_ (.A(net788),
    .B(_0682_),
    .X(_0683_));
 sky130_fd_sc_hd__or2_1 _2206_ (.A(net788),
    .B(_0682_),
    .X(_0684_));
 sky130_fd_sc_hd__a32o_1 _2207_ (.A1(_0472_),
    .A2(_0608_),
    .A3(_0644_),
    .B1(_0672_),
    .B2(_0590_),
    .X(_0685_));
 sky130_fd_sc_hd__and3_1 _2208_ (.A(_0482_),
    .B(_0545_),
    .C(_0563_),
    .X(_0686_));
 sky130_fd_sc_hd__a31o_1 _2209_ (.A1(_0483_),
    .A2(_0608_),
    .A3(_0626_),
    .B1(_0686_),
    .X(_0687_));
 sky130_fd_sc_hd__a32o_1 _2210_ (.A1(_0483_),
    .A2(_0527_),
    .A3(_0572_),
    .B1(_0685_),
    .B2(_0568_),
    .X(_0688_));
 sky130_fd_sc_hd__a21oi_1 _2211_ (.A1(_0571_),
    .A2(_0687_),
    .B1(_0688_),
    .Y(_0689_));
 sky130_fd_sc_hd__nor2_1 _2212_ (.A(_0484_),
    .B(_0606_),
    .Y(_0690_));
 sky130_fd_sc_hd__a211o_1 _2213_ (.A1(_0484_),
    .A2(_0689_),
    .B1(_0690_),
    .C1(net65),
    .X(_0691_));
 sky130_fd_sc_hd__nor2_1 _2214_ (.A(_0458_),
    .B(_0469_),
    .Y(_0692_));
 sky130_fd_sc_hd__or3_1 _2215_ (.A(net63),
    .B(_0677_),
    .C(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__o22a_1 _2216_ (.A1(net79),
    .A2(_1799_),
    .B1(_0689_),
    .B2(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__o21a_1 _2217_ (.A1(net61),
    .A2(_0694_),
    .B1(_0691_),
    .X(_0695_));
 sky130_fd_sc_hd__and2b_1 _2218_ (.A_N(\S8x305.ALU_in1[5] ),
    .B(_0695_),
    .X(_0696_));
 sky130_fd_sc_hd__nand2b_1 _2219_ (.A_N(net812),
    .B(_0695_),
    .Y(_0697_));
 sky130_fd_sc_hd__or2_1 _2220_ (.A(_0480_),
    .B(_0526_),
    .X(_0698_));
 sky130_fd_sc_hd__and3_1 _2221_ (.A(_0482_),
    .B(_0670_),
    .C(_0671_),
    .X(_0699_));
 sky130_fd_sc_hd__and3_1 _2222_ (.A(_0483_),
    .B(_0661_),
    .C(_0662_),
    .X(_0700_));
 sky130_fd_sc_hd__a21o_1 _2223_ (.A1(_0661_),
    .A2(_0665_),
    .B1(_0473_),
    .X(_0701_));
 sky130_fd_sc_hd__a21o_1 _2224_ (.A1(_0664_),
    .A2(_0668_),
    .B1(_0472_),
    .X(_0702_));
 sky130_fd_sc_hd__o311a_1 _2225_ (.A1(_0572_),
    .A2(_0699_),
    .A3(_0700_),
    .B1(_0698_),
    .C1(_0569_),
    .X(_0703_));
 sky130_fd_sc_hd__a31o_1 _2226_ (.A1(_0568_),
    .A2(_0701_),
    .A3(_0702_),
    .B1(_0703_),
    .X(_0704_));
 sky130_fd_sc_hd__mux2_1 _2227_ (.A0(_0704_),
    .A1(_0624_),
    .S(_1821_),
    .X(_0705_));
 sky130_fd_sc_hd__and2_1 _2228_ (.A(_0459_),
    .B(_0649_),
    .X(_0706_));
 sky130_fd_sc_hd__or2_1 _2229_ (.A(_0677_),
    .B(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__nor2_1 _2230_ (.A(net63),
    .B(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__a22o_1 _2231_ (.A1(\S8x305.iv_latch[4] ),
    .A2(net63),
    .B1(_0704_),
    .B2(_0708_),
    .X(_0709_));
 sky130_fd_sc_hd__mux2_1 _2232_ (.A0(_0705_),
    .A1(_0709_),
    .S(_1824_),
    .X(_0710_));
 sky130_fd_sc_hd__and2_1 _2233_ (.A(\S8x305.ALU_in1[4] ),
    .B(_0710_),
    .X(_0711_));
 sky130_fd_sc_hd__xnor2_1 _2234_ (.A(\S8x305.ALU_in1[4] ),
    .B(_0710_),
    .Y(_0712_));
 sky130_fd_sc_hd__inv_2 _2235_ (.A(_0712_),
    .Y(_0713_));
 sky130_fd_sc_hd__a21o_1 _2236_ (.A1(_0608_),
    .A2(_0644_),
    .B1(_0472_),
    .X(_0714_));
 sky130_fd_sc_hd__a21o_1 _2237_ (.A1(_0545_),
    .A2(_0626_),
    .B1(_0473_),
    .X(_0715_));
 sky130_fd_sc_hd__and3_1 _2238_ (.A(_0479_),
    .B(_0569_),
    .C(_0590_),
    .X(_0716_));
 sky130_fd_sc_hd__a31o_1 _2239_ (.A1(_0568_),
    .A2(_0714_),
    .A3(_0715_),
    .B1(_0716_),
    .X(_0717_));
 sky130_fd_sc_hd__a21o_1 _2240_ (.A1(_0565_),
    .A2(_0571_),
    .B1(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__or2_1 _2241_ (.A(_0484_),
    .B(_0543_),
    .X(_0719_));
 sky130_fd_sc_hd__o211a_1 _2242_ (.A1(_0485_),
    .A2(_0718_),
    .B1(_0719_),
    .C1(net61),
    .X(_0720_));
 sky130_fd_sc_hd__a22o_2 _2243_ (.A1(\S8x305.iv_latch[3] ),
    .A2(_1798_),
    .B1(_0678_),
    .B2(_0718_),
    .X(_0721_));
 sky130_fd_sc_hd__a21oi_2 _2244_ (.A1(_1824_),
    .A2(_0721_),
    .B1(_0720_),
    .Y(_0722_));
 sky130_fd_sc_hd__and2b_1 _2245_ (.A_N(\S8x305.ALU_in1[3] ),
    .B(_0722_),
    .X(_0723_));
 sky130_fd_sc_hd__inv_2 _2246_ (.A(_0723_),
    .Y(_0724_));
 sky130_fd_sc_hd__and2b_1 _2247_ (.A_N(_0722_),
    .B(\S8x305.ALU_in1[3] ),
    .X(_0725_));
 sky130_fd_sc_hd__a21o_1 _2248_ (.A1(_0662_),
    .A2(_0671_),
    .B1(_0473_),
    .X(_0726_));
 sky130_fd_sc_hd__a21o_1 _2249_ (.A1(_0661_),
    .A2(_0665_),
    .B1(_0472_),
    .X(_0727_));
 sky130_fd_sc_hd__a21o_1 _2250_ (.A1(_0726_),
    .A2(_0727_),
    .B1(_0569_),
    .X(_0728_));
 sky130_fd_sc_hd__a211o_1 _2251_ (.A1(_0480_),
    .A2(_0673_),
    .B1(_0669_),
    .C1(_0568_),
    .X(_0729_));
 sky130_fd_sc_hd__a21oi_1 _2252_ (.A1(_0676_),
    .A2(_0677_),
    .B1(net63),
    .Y(_0730_));
 sky130_fd_sc_hd__a32o_1 _2253_ (.A1(_0728_),
    .A2(_0729_),
    .A3(_0730_),
    .B1(net63),
    .B2(\S8x305.iv_latch[2] ),
    .X(_0731_));
 sky130_fd_sc_hd__or2_2 _2254_ (.A(net61),
    .B(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__a21o_1 _2255_ (.A1(_0728_),
    .A2(_0729_),
    .B1(_0485_),
    .X(_0733_));
 sky130_fd_sc_hd__or2_1 _2256_ (.A(_0484_),
    .B(_0561_),
    .X(_0734_));
 sky130_fd_sc_hd__a21o_1 _2257_ (.A1(_0733_),
    .A2(_0734_),
    .B1(net65),
    .X(_0735_));
 sky130_fd_sc_hd__nand2_1 _2258_ (.A(_0732_),
    .B(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__a21oi_1 _2259_ (.A1(_0732_),
    .A2(_0735_),
    .B1(\S8x305.ALU_in1[2] ),
    .Y(_0737_));
 sky130_fd_sc_hd__a21o_1 _2260_ (.A1(_0732_),
    .A2(_0735_),
    .B1(\S8x305.ALU_in1[2] ),
    .X(_0738_));
 sky130_fd_sc_hd__and3_1 _2261_ (.A(\S8x305.ALU_in1[2] ),
    .B(_0732_),
    .C(_0735_),
    .X(_0739_));
 sky130_fd_sc_hd__a211oi_2 _2262_ (.A1(_0481_),
    .A2(_0526_),
    .B1(_0568_),
    .C1(_0685_),
    .Y(_0740_));
 sky130_fd_sc_hd__a21o_1 _2263_ (.A1(_0509_),
    .A2(_0563_),
    .B1(_0473_),
    .X(_0741_));
 sky130_fd_sc_hd__a21o_1 _2264_ (.A1(_0545_),
    .A2(_0626_),
    .B1(_0472_),
    .X(_0742_));
 sky130_fd_sc_hd__a21oi_2 _2265_ (.A1(_0741_),
    .A2(_0742_),
    .B1(_0569_),
    .Y(_0743_));
 sky130_fd_sc_hd__or3_1 _2266_ (.A(_0485_),
    .B(_0740_),
    .C(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__a21oi_1 _2267_ (.A1(_1821_),
    .A2(_0506_),
    .B1(net66),
    .Y(_0745_));
 sky130_fd_sc_hd__and3_1 _2268_ (.A(_0458_),
    .B(_0468_),
    .C(_0474_),
    .X(_0746_));
 sky130_fd_sc_hd__or2_1 _2269_ (.A(_1798_),
    .B(_0746_),
    .X(_0747_));
 sky130_fd_sc_hd__o32ai_4 _2270_ (.A1(_0740_),
    .A2(_0743_),
    .A3(_0747_),
    .B1(_1799_),
    .B2(net56),
    .Y(_0748_));
 sky130_fd_sc_hd__a2bb2o_2 _2271_ (.A1_N(net61),
    .A2_N(_0748_),
    .B1(_0744_),
    .B2(_0745_),
    .X(_0749_));
 sky130_fd_sc_hd__nor2_1 _2272_ (.A(_1772_),
    .B(_0749_),
    .Y(_0750_));
 sky130_fd_sc_hd__o31a_1 _2273_ (.A1(_0477_),
    .A2(_0507_),
    .A3(_0508_),
    .B1(_0472_),
    .X(_0751_));
 sky130_fd_sc_hd__a31o_1 _2274_ (.A1(_0473_),
    .A2(_0662_),
    .A3(_0671_),
    .B1(_0751_),
    .X(_0752_));
 sky130_fd_sc_hd__o21a_1 _2275_ (.A1(_0480_),
    .A2(_0526_),
    .B1(_0568_),
    .X(_0753_));
 sky130_fd_sc_hd__a32o_1 _2276_ (.A1(_0569_),
    .A2(_0701_),
    .A3(_0702_),
    .B1(_0752_),
    .B2(_0753_),
    .X(_0754_));
 sky130_fd_sc_hd__or2_1 _2277_ (.A(net66),
    .B(_0525_),
    .X(_0755_));
 sky130_fd_sc_hd__o21a_1 _2278_ (.A1(net61),
    .A2(_0754_),
    .B1(_0755_),
    .X(_0756_));
 sky130_fd_sc_hd__mux2_1 _2279_ (.A0(_0754_),
    .A1(_0756_),
    .S(_0485_),
    .X(_0757_));
 sky130_fd_sc_hd__and2_1 _2280_ (.A(\S8x305.ALU_in1[0] ),
    .B(_0757_),
    .X(_0758_));
 sky130_fd_sc_hd__xnor2_2 _2281_ (.A(\S8x305.ALU_in1[1] ),
    .B(_0749_),
    .Y(_0759_));
 sky130_fd_sc_hd__a21oi_1 _2282_ (.A1(_0758_),
    .A2(_0759_),
    .B1(_0750_),
    .Y(_0760_));
 sky130_fd_sc_hd__a211o_1 _2283_ (.A1(_0758_),
    .A2(_0759_),
    .B1(_0739_),
    .C1(_0750_),
    .X(_0761_));
 sky130_fd_sc_hd__a21o_1 _2284_ (.A1(_0738_),
    .A2(_0761_),
    .B1(_0725_),
    .X(_0762_));
 sky130_fd_sc_hd__or3b_1 _2285_ (.A(_0712_),
    .B(_0723_),
    .C_N(_0762_),
    .X(_0763_));
 sky130_fd_sc_hd__and2b_1 _2286_ (.A_N(_0695_),
    .B(\S8x305.ALU_in1[5] ),
    .X(_0764_));
 sky130_fd_sc_hd__a311o_1 _2287_ (.A1(_0713_),
    .A2(_0724_),
    .A3(_0762_),
    .B1(_0764_),
    .C1(_0711_),
    .X(_0765_));
 sky130_fd_sc_hd__nor2_1 _2288_ (.A(_0696_),
    .B(_0764_),
    .Y(_0766_));
 sky130_fd_sc_hd__inv_2 _2289_ (.A(_0766_),
    .Y(_0767_));
 sky130_fd_sc_hd__a31o_1 _2290_ (.A1(_0684_),
    .A2(_0697_),
    .A3(_0765_),
    .B1(_0683_),
    .X(_0768_));
 sky130_fd_sc_hd__or2_1 _2291_ (.A(_0657_),
    .B(_0768_),
    .X(_0769_));
 sky130_fd_sc_hd__a21oi_1 _2292_ (.A1(_0657_),
    .A2(_0768_),
    .B1(_1796_),
    .Y(_0770_));
 sky130_fd_sc_hd__a21oi_1 _2293_ (.A1(_0769_),
    .A2(_0770_),
    .B1(_0660_),
    .Y(_0771_));
 sky130_fd_sc_hd__a21oi_1 _2294_ (.A1(_1831_),
    .A2(_0654_),
    .B1(_0771_),
    .Y(_0772_));
 sky130_fd_sc_hd__a211o_1 _2295_ (.A1(_1831_),
    .A2(_0654_),
    .B1(_0771_),
    .C1(_0464_),
    .X(_0773_));
 sky130_fd_sc_hd__or3_1 _2296_ (.A(net61),
    .B(_1825_),
    .C(_1834_),
    .X(_0774_));
 sky130_fd_sc_hd__a22o_1 _2297_ (.A1(net66),
    .A2(_1833_),
    .B1(_0658_),
    .B2(_1792_),
    .X(_0775_));
 sky130_fd_sc_hd__o22a_1 _2298_ (.A1(_1814_),
    .A2(_0774_),
    .B1(_0775_),
    .B2(_0477_),
    .X(_0776_));
 sky130_fd_sc_hd__mux2_4 _2299_ (.A0(_1814_),
    .A1(_0776_),
    .S(_0463_),
    .X(_0777_));
 sky130_fd_sc_hd__inv_2 _2300_ (.A(_0777_),
    .Y(_0778_));
 sky130_fd_sc_hd__nand2_1 _2301_ (.A(_0460_),
    .B(_0464_),
    .Y(_0779_));
 sky130_fd_sc_hd__o22a_2 _2302_ (.A1(_1806_),
    .A2(_0774_),
    .B1(_0775_),
    .B2(_0472_),
    .X(_0780_));
 sky130_fd_sc_hd__or2_1 _2303_ (.A(_1806_),
    .B(_0463_),
    .X(_0781_));
 sky130_fd_sc_hd__o21ai_2 _2304_ (.A1(_0464_),
    .A2(_0780_),
    .B1(_0781_),
    .Y(_0782_));
 sky130_fd_sc_hd__o21a_2 _2305_ (.A1(_0464_),
    .A2(_0780_),
    .B1(_0781_),
    .X(_0783_));
 sky130_fd_sc_hd__or2_1 _2306_ (.A(_1832_),
    .B(_0682_),
    .X(_0784_));
 sky130_fd_sc_hd__nand2b_1 _2307_ (.A_N(_0683_),
    .B(_0684_),
    .Y(_0785_));
 sky130_fd_sc_hd__inv_2 _2308_ (.A(_0785_),
    .Y(_0786_));
 sky130_fd_sc_hd__o221a_1 _2309_ (.A1(_1837_),
    .A2(_0683_),
    .B1(_0786_),
    .B2(_1787_),
    .C1(_0659_),
    .X(_0787_));
 sky130_fd_sc_hd__a21oi_1 _2310_ (.A1(_0697_),
    .A2(_0765_),
    .B1(_0786_),
    .Y(_0788_));
 sky130_fd_sc_hd__a31o_1 _2311_ (.A1(_0697_),
    .A2(_0765_),
    .A3(_0786_),
    .B1(_1796_),
    .X(_0789_));
 sky130_fd_sc_hd__o21bai_1 _2312_ (.A1(_0788_),
    .A2(_0789_),
    .B1_N(_0787_),
    .Y(_0790_));
 sky130_fd_sc_hd__and2_1 _2313_ (.A(_0784_),
    .B(_0790_),
    .X(_0791_));
 sky130_fd_sc_hd__a21o_1 _2314_ (.A1(_0784_),
    .A2(_0790_),
    .B1(_0464_),
    .X(_0792_));
 sky130_fd_sc_hd__nor2_2 _2315_ (.A(net66),
    .B(_0468_),
    .Y(_0793_));
 sky130_fd_sc_hd__or2_1 _2316_ (.A(_0463_),
    .B(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__a21oi_1 _2317_ (.A1(_0792_),
    .A2(_0794_),
    .B1(_0777_),
    .Y(_0795_));
 sky130_fd_sc_hd__a311o_1 _2318_ (.A1(_0773_),
    .A2(_0777_),
    .A3(_0779_),
    .B1(_0782_),
    .C1(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__o22a_1 _2319_ (.A1(_1830_),
    .A2(_0774_),
    .B1(_0775_),
    .B2(_0568_),
    .X(_0797_));
 sky130_fd_sc_hd__mux2_2 _2320_ (.A0(_1830_),
    .A1(_0797_),
    .S(_0463_),
    .X(_0798_));
 sky130_fd_sc_hd__inv_2 _2321_ (.A(_0798_),
    .Y(_0799_));
 sky130_fd_sc_hd__o221a_1 _2322_ (.A1(_1837_),
    .A2(_0764_),
    .B1(_0766_),
    .B2(_1787_),
    .C1(_0659_),
    .X(_0800_));
 sky130_fd_sc_hd__a31oi_1 _2323_ (.A1(_0713_),
    .A2(_0724_),
    .A3(_0762_),
    .B1(_0711_),
    .Y(_0801_));
 sky130_fd_sc_hd__a311o_1 _2324_ (.A1(_0713_),
    .A2(_0724_),
    .A3(_0762_),
    .B1(_0766_),
    .C1(_0711_),
    .X(_0802_));
 sky130_fd_sc_hd__o211a_1 _2325_ (.A1(_0767_),
    .A2(_0801_),
    .B1(_0802_),
    .C1(_0658_),
    .X(_0803_));
 sky130_fd_sc_hd__a2bb2o_1 _2326_ (.A1_N(_0800_),
    .A2_N(_0803_),
    .B1(_1831_),
    .B2(_0695_),
    .X(_0804_));
 sky130_fd_sc_hd__and2_2 _2327_ (.A(net61),
    .B(_0474_),
    .X(_0805_));
 sky130_fd_sc_hd__nor2_1 _2328_ (.A(_0463_),
    .B(_0805_),
    .Y(_0806_));
 sky130_fd_sc_hd__a21o_1 _2329_ (.A1(_0724_),
    .A2(_0762_),
    .B1(_0713_),
    .X(_0807_));
 sky130_fd_sc_hd__o221a_1 _2330_ (.A1(_1837_),
    .A2(_0711_),
    .B1(_0713_),
    .B2(_1787_),
    .C1(_0659_),
    .X(_0808_));
 sky130_fd_sc_hd__a31o_1 _2331_ (.A1(_0658_),
    .A2(_0763_),
    .A3(_0807_),
    .B1(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__o21a_1 _2332_ (.A1(_1832_),
    .A2(_0710_),
    .B1(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__o21ai_1 _2333_ (.A1(_0464_),
    .A2(_0810_),
    .B1(_1820_),
    .Y(_0811_));
 sky130_fd_sc_hd__o211ai_1 _2334_ (.A1(_0464_),
    .A2(_0810_),
    .B1(_0778_),
    .C1(_1820_),
    .Y(_0812_));
 sky130_fd_sc_hd__a211o_1 _2335_ (.A1(_0463_),
    .A2(_0804_),
    .B1(_0806_),
    .C1(_0778_),
    .X(_0813_));
 sky130_fd_sc_hd__a21oi_1 _2336_ (.A1(_0812_),
    .A2(_0813_),
    .B1(_0783_),
    .Y(_0814_));
 sky130_fd_sc_hd__nor2_1 _2337_ (.A(_0799_),
    .B(_0814_),
    .Y(_0815_));
 sky130_fd_sc_hd__or2_1 _2338_ (.A(_0758_),
    .B(_0759_),
    .X(_0816_));
 sky130_fd_sc_hd__a21oi_1 _2339_ (.A1(_0758_),
    .A2(_0759_),
    .B1(_0659_),
    .Y(_0817_));
 sky130_fd_sc_hd__o221a_1 _2340_ (.A1(_1837_),
    .A2(_0750_),
    .B1(_0759_),
    .B2(_1787_),
    .C1(_0659_),
    .X(_0818_));
 sky130_fd_sc_hd__a21oi_1 _2341_ (.A1(_0816_),
    .A2(_0817_),
    .B1(_0818_),
    .Y(_0819_));
 sky130_fd_sc_hd__a21oi_2 _2342_ (.A1(_1831_),
    .A2(_0749_),
    .B1(_0819_),
    .Y(_0820_));
 sky130_fd_sc_hd__mux2_1 _2343_ (.A0(_1804_),
    .A1(_0820_),
    .S(_0463_),
    .X(_0821_));
 sky130_fd_sc_hd__a22o_1 _2344_ (.A1(net789),
    .A2(_1788_),
    .B1(_1837_),
    .B2(_0757_),
    .X(_0822_));
 sky130_fd_sc_hd__mux2_1 _2345_ (.A0(_0822_),
    .A1(_1787_),
    .S(_0758_),
    .X(_0823_));
 sky130_fd_sc_hd__mux2_1 _2346_ (.A0(_1807_),
    .A1(_0823_),
    .S(_0463_),
    .X(_0824_));
 sky130_fd_sc_hd__mux2_1 _2347_ (.A0(_0821_),
    .A1(_0824_),
    .S(_0778_),
    .X(_0825_));
 sky130_fd_sc_hd__inv_2 _2348_ (.A(_0825_),
    .Y(_0826_));
 sky130_fd_sc_hd__and2_1 _2349_ (.A(_1826_),
    .B(_0464_),
    .X(_0827_));
 sky130_fd_sc_hd__or2_1 _2350_ (.A(_0737_),
    .B(_0739_),
    .X(_0828_));
 sky130_fd_sc_hd__a2bb2o_1 _2351_ (.A1_N(_1837_),
    .A2_N(_0739_),
    .B1(_0828_),
    .B2(_1788_),
    .X(_0829_));
 sky130_fd_sc_hd__and2_1 _2352_ (.A(_0760_),
    .B(_0828_),
    .X(_0830_));
 sky130_fd_sc_hd__o21ai_1 _2353_ (.A1(_0760_),
    .A2(_0828_),
    .B1(_0658_),
    .Y(_0831_));
 sky130_fd_sc_hd__o22a_1 _2354_ (.A1(_0658_),
    .A2(_0829_),
    .B1(_0830_),
    .B2(_0831_),
    .X(_0832_));
 sky130_fd_sc_hd__a21oi_2 _2355_ (.A1(_1831_),
    .A2(_0736_),
    .B1(_0832_),
    .Y(_0833_));
 sky130_fd_sc_hd__xnor2_1 _2356_ (.A(\S8x305.ALU_in1[3] ),
    .B(_0722_),
    .Y(_0834_));
 sky130_fd_sc_hd__o221a_1 _2357_ (.A1(_1837_),
    .A2(_0725_),
    .B1(_0834_),
    .B2(_1787_),
    .C1(_0659_),
    .X(_0835_));
 sky130_fd_sc_hd__a21oi_1 _2358_ (.A1(_0738_),
    .A2(_0761_),
    .B1(_0834_),
    .Y(_0836_));
 sky130_fd_sc_hd__a31o_1 _2359_ (.A1(_0738_),
    .A2(_0761_),
    .A3(_0834_),
    .B1(_0659_),
    .X(_0837_));
 sky130_fd_sc_hd__nor2_1 _2360_ (.A(_0836_),
    .B(_0837_),
    .Y(_0838_));
 sky130_fd_sc_hd__o2bb2a_1 _2361_ (.A1_N(_1831_),
    .A2_N(_0722_),
    .B1(_0835_),
    .B2(_0838_),
    .X(_0839_));
 sky130_fd_sc_hd__mux2_1 _2362_ (.A0(_0436_),
    .A1(_0839_),
    .S(_0463_),
    .X(_0840_));
 sky130_fd_sc_hd__a211o_1 _2363_ (.A1(_0463_),
    .A2(_0833_),
    .B1(_0827_),
    .C1(_0777_),
    .X(_0841_));
 sky130_fd_sc_hd__o21ai_1 _2364_ (.A1(_0778_),
    .A2(_0840_),
    .B1(_0841_),
    .Y(_0842_));
 sky130_fd_sc_hd__mux2_1 _2365_ (.A0(_0826_),
    .A1(_0842_),
    .S(_0783_),
    .X(_0843_));
 sky130_fd_sc_hd__and2_1 _2366_ (.A(_0799_),
    .B(_0843_),
    .X(_0844_));
 sky130_fd_sc_hd__a21o_1 _2367_ (.A1(_0796_),
    .A2(_0815_),
    .B1(_0844_),
    .X(_0845_));
 sky130_fd_sc_hd__o21ai_4 _2368_ (.A1(_1799_),
    .A2(net60),
    .B1(_0797_),
    .Y(_0846_));
 sky130_fd_sc_hd__nand2_2 _2369_ (.A(_1803_),
    .B(_0780_),
    .Y(_0847_));
 sky130_fd_sc_hd__and2_1 _2370_ (.A(_1813_),
    .B(_0776_),
    .X(_0848_));
 sky130_fd_sc_hd__nand2_1 _2371_ (.A(_1813_),
    .B(_0776_),
    .Y(_0849_));
 sky130_fd_sc_hd__a21oi_1 _2372_ (.A1(_0692_),
    .A2(_0848_),
    .B1(_0707_),
    .Y(_0850_));
 sky130_fd_sc_hd__nor2_1 _2373_ (.A(_0676_),
    .B(_0848_),
    .Y(_0851_));
 sky130_fd_sc_hd__o21bai_1 _2374_ (.A1(_0458_),
    .A2(_0851_),
    .B1_N(_0847_),
    .Y(_0852_));
 sky130_fd_sc_hd__a2bb2o_1 _2375_ (.A1_N(_0677_),
    .A2_N(_0852_),
    .B1(_0847_),
    .B2(_0850_),
    .X(_0853_));
 sky130_fd_sc_hd__and3_1 _2376_ (.A(_1813_),
    .B(_0746_),
    .C(_0776_),
    .X(_0854_));
 sky130_fd_sc_hd__inv_2 _2377_ (.A(_0854_),
    .Y(_0855_));
 sky130_fd_sc_hd__or3_1 _2378_ (.A(_0459_),
    .B(_0649_),
    .C(_0851_),
    .X(_0856_));
 sky130_fd_sc_hd__mux2_1 _2379_ (.A0(_0856_),
    .A1(_0855_),
    .S(_0847_),
    .X(_0857_));
 sky130_fd_sc_hd__mux2_2 _2380_ (.A0(_0853_),
    .A1(_0857_),
    .S(_0846_),
    .X(_0858_));
 sky130_fd_sc_hd__o21ai_1 _2381_ (.A1(net793),
    .A2(_0858_),
    .B1(net65),
    .Y(_0859_));
 sky130_fd_sc_hd__a21oi_1 _2382_ (.A1(_0845_),
    .A2(_0858_),
    .B1(_0859_),
    .Y(_0860_));
 sky130_fd_sc_hd__a31oi_4 _2383_ (.A1(net65),
    .A2(_1825_),
    .A3(_1833_),
    .B1(_0484_),
    .Y(_0861_));
 sky130_fd_sc_hd__a31o_2 _2384_ (.A1(net65),
    .A2(_1825_),
    .A3(_1833_),
    .B1(_0484_),
    .X(_0862_));
 sky130_fd_sc_hd__nand2_1 _2385_ (.A(_0858_),
    .B(_0861_),
    .Y(_0863_));
 sky130_fd_sc_hd__a211o_1 _2386_ (.A1(_0796_),
    .A2(_0815_),
    .B1(_0844_),
    .C1(_0863_),
    .X(_0864_));
 sky130_fd_sc_hd__nand2_1 _2387_ (.A(_0772_),
    .B(_0862_),
    .Y(_0865_));
 sky130_fd_sc_hd__a31oi_1 _2388_ (.A1(_0456_),
    .A2(_0864_),
    .A3(_0865_),
    .B1(_0462_),
    .Y(_0866_));
 sky130_fd_sc_hd__o31a_1 _2389_ (.A1(_0456_),
    .A2(_0460_),
    .A3(_0860_),
    .B1(_0866_),
    .X(_0867_));
 sky130_fd_sc_hd__a211oi_2 _2390_ (.A1(net488),
    .A2(_0453_),
    .B1(net82),
    .C1(_1740_),
    .Y(_0868_));
 sky130_fd_sc_hd__a211o_1 _2391_ (.A1(net488),
    .A2(_0453_),
    .B1(net83),
    .C1(_1740_),
    .X(_0869_));
 sky130_fd_sc_hd__and3_1 _2392_ (.A(_0456_),
    .B(_0461_),
    .C(_0861_),
    .X(_0870_));
 sky130_fd_sc_hd__or3_2 _2393_ (.A(_0455_),
    .B(_0462_),
    .C(_0862_),
    .X(_0871_));
 sky130_fd_sc_hd__o21a_1 _2394_ (.A1(_0858_),
    .A2(_0871_),
    .B1(_0868_),
    .X(_0872_));
 sky130_fd_sc_hd__or4_2 _2395_ (.A(\cmdr[7] ),
    .B(\cmdr[6] ),
    .C(\cmdr[5] ),
    .D(\cmdr[4] ),
    .X(_0873_));
 sky130_fd_sc_hd__nor3b_4 _2396_ (.A(net31),
    .B(_0873_),
    .C_N(net2),
    .Y(_0874_));
 sky130_fd_sc_hd__mux4_1 _2397_ (.A0(\memory[0][0] ),
    .A1(\memory[1][0] ),
    .A2(\memory[2][0] ),
    .A3(\memory[3][0] ),
    .S0(net90),
    .S1(net88),
    .X(_0875_));
 sky130_fd_sc_hd__nand2b_1 _2398_ (.A_N(net86),
    .B(_0875_),
    .Y(_0876_));
 sky130_fd_sc_hd__mux4_1 _2399_ (.A0(\memory[4][0] ),
    .A1(\memory[6][0] ),
    .A2(\memory[5][0] ),
    .A3(\memory[7][0] ),
    .S0(net87),
    .S1(net89),
    .X(_0877_));
 sky130_fd_sc_hd__a21oi_1 _2400_ (.A1(net86),
    .A2(_0877_),
    .B1(_0003_),
    .Y(_0878_));
 sky130_fd_sc_hd__mux4_1 _2401_ (.A0(\memory[8][0] ),
    .A1(\memory[9][0] ),
    .A2(\memory[10][0] ),
    .A3(\memory[11][0] ),
    .S0(net89),
    .S1(net87),
    .X(_0879_));
 sky130_fd_sc_hd__nand2b_1 _2402_ (.A_N(net86),
    .B(_0879_),
    .Y(_0880_));
 sky130_fd_sc_hd__mux4_1 _2403_ (.A0(\memory[12][0] ),
    .A1(\memory[13][0] ),
    .A2(\memory[14][0] ),
    .A3(\memory[15][0] ),
    .S0(net90),
    .S1(net88),
    .X(_0881_));
 sky130_fd_sc_hd__nand2_1 _2404_ (.A(net86),
    .B(_0881_),
    .Y(_0882_));
 sky130_fd_sc_hd__a32o_1 _2405_ (.A1(_0003_),
    .A2(_0880_),
    .A3(_0882_),
    .B1(_0876_),
    .B2(_0878_),
    .X(_0883_));
 sky130_fd_sc_hd__mux2_1 _2406_ (.A0(_1781_),
    .A1(_0883_),
    .S(_0874_),
    .X(_0884_));
 sky130_fd_sc_hd__or4_1 _2407_ (.A(net496),
    .B(net461),
    .C(net486),
    .D(net516),
    .X(_0885_));
 sky130_fd_sc_hd__or4_1 _2408_ (.A(net466),
    .B(net435),
    .C(net457),
    .D(net481),
    .X(_0886_));
 sky130_fd_sc_hd__nor2_1 _2409_ (.A(_0885_),
    .B(_0886_),
    .Y(_0887_));
 sky130_fd_sc_hd__and3_4 _2410_ (.A(net1),
    .B(_0448_),
    .C(_0887_),
    .X(_0888_));
 sky130_fd_sc_hd__mux2_1 _2411_ (.A0(_0884_),
    .A1(net15),
    .S(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__a21bo_1 _2412_ (.A1(_0462_),
    .A2(_0889_),
    .B1_N(_0872_),
    .X(_0890_));
 sky130_fd_sc_hd__o221a_1 _2413_ (.A1(net793),
    .A2(_0872_),
    .B1(_0890_),
    .B2(_0867_),
    .C1(net100),
    .X(_0004_));
 sky130_fd_sc_hd__a211oi_1 _2414_ (.A1(_0463_),
    .A2(_0804_),
    .B1(_0806_),
    .C1(_0777_),
    .Y(_0891_));
 sky130_fd_sc_hd__a31o_1 _2415_ (.A1(_0777_),
    .A2(_0792_),
    .A3(_0794_),
    .B1(_0891_),
    .X(_0892_));
 sky130_fd_sc_hd__nor2_1 _2416_ (.A(_0777_),
    .B(_0840_),
    .Y(_0893_));
 sky130_fd_sc_hd__a211oi_1 _2417_ (.A1(_0777_),
    .A2(_0811_),
    .B1(_0893_),
    .C1(_0783_),
    .Y(_0894_));
 sky130_fd_sc_hd__a211o_1 _2418_ (.A1(_0783_),
    .A2(_0892_),
    .B1(_0894_),
    .C1(_0799_),
    .X(_0895_));
 sky130_fd_sc_hd__a21oi_1 _2419_ (.A1(_0706_),
    .A2(_0848_),
    .B1(_0677_),
    .Y(_0896_));
 sky130_fd_sc_hd__inv_2 _2420_ (.A(_0896_),
    .Y(_0897_));
 sky130_fd_sc_hd__nand2_1 _2421_ (.A(_0469_),
    .B(_0849_),
    .Y(_0898_));
 sky130_fd_sc_hd__a31o_1 _2422_ (.A1(_0459_),
    .A2(_0676_),
    .A3(_0898_),
    .B1(_0677_),
    .X(_0899_));
 sky130_fd_sc_hd__mux2_1 _2423_ (.A0(_0899_),
    .A1(_0897_),
    .S(_0847_),
    .X(_0900_));
 sky130_fd_sc_hd__and3_1 _2424_ (.A(_0676_),
    .B(_0677_),
    .C(_0898_),
    .X(_0901_));
 sky130_fd_sc_hd__mux2_1 _2425_ (.A0(_0901_),
    .A1(_0849_),
    .S(_0847_),
    .X(_0902_));
 sky130_fd_sc_hd__mux2_1 _2426_ (.A0(_0900_),
    .A1(_0902_),
    .S(_0846_),
    .X(_0903_));
 sky130_fd_sc_hd__or2_1 _2427_ (.A(_0777_),
    .B(_0821_),
    .X(_0904_));
 sky130_fd_sc_hd__a211o_1 _2428_ (.A1(_0463_),
    .A2(_0833_),
    .B1(_0827_),
    .C1(_0778_),
    .X(_0905_));
 sky130_fd_sc_hd__nand2_1 _2429_ (.A(_0777_),
    .B(_0824_),
    .Y(_0906_));
 sky130_fd_sc_hd__nor2_1 _2430_ (.A(_0783_),
    .B(_0906_),
    .Y(_0907_));
 sky130_fd_sc_hd__a31oi_2 _2431_ (.A1(_0783_),
    .A2(_0904_),
    .A3(_0905_),
    .B1(_0907_),
    .Y(_0908_));
 sky130_fd_sc_hd__a21oi_1 _2432_ (.A1(_0799_),
    .A2(_0908_),
    .B1(_0903_),
    .Y(_0909_));
 sky130_fd_sc_hd__a22o_1 _2433_ (.A1(net400),
    .A2(_0903_),
    .B1(_0909_),
    .B2(_0895_),
    .X(_0910_));
 sky130_fd_sc_hd__a21o_1 _2434_ (.A1(net65),
    .A2(_0910_),
    .B1(_0793_),
    .X(_0911_));
 sky130_fd_sc_hd__or2_1 _2435_ (.A(_0791_),
    .B(_0861_),
    .X(_0912_));
 sky130_fd_sc_hd__a21o_1 _2436_ (.A1(_0895_),
    .A2(_0909_),
    .B1(_0862_),
    .X(_0913_));
 sky130_fd_sc_hd__a21o_1 _2437_ (.A1(_0912_),
    .A2(_0913_),
    .B1(_0455_),
    .X(_0914_));
 sky130_fd_sc_hd__o211a_1 _2438_ (.A1(_0456_),
    .A2(_0911_),
    .B1(_0914_),
    .C1(_0461_),
    .X(_0915_));
 sky130_fd_sc_hd__a21oi_1 _2439_ (.A1(_0870_),
    .A2(_0903_),
    .B1(_0869_),
    .Y(_0916_));
 sky130_fd_sc_hd__mux4_1 _2440_ (.A0(\memory[0][1] ),
    .A1(\memory[1][1] ),
    .A2(\memory[2][1] ),
    .A3(\memory[3][1] ),
    .S0(net90),
    .S1(net88),
    .X(_0917_));
 sky130_fd_sc_hd__nand2b_1 _2441_ (.A_N(net85),
    .B(_0917_),
    .Y(_0918_));
 sky130_fd_sc_hd__mux4_1 _2442_ (.A0(\memory[4][1] ),
    .A1(\memory[6][1] ),
    .A2(\memory[5][1] ),
    .A3(\memory[7][1] ),
    .S0(net87),
    .S1(net89),
    .X(_0919_));
 sky130_fd_sc_hd__a21oi_1 _2443_ (.A1(net85),
    .A2(_0919_),
    .B1(_0003_),
    .Y(_0920_));
 sky130_fd_sc_hd__mux4_1 _2444_ (.A0(\memory[8][1] ),
    .A1(\memory[9][1] ),
    .A2(\memory[10][1] ),
    .A3(\memory[11][1] ),
    .S0(net89),
    .S1(net87),
    .X(_0921_));
 sky130_fd_sc_hd__nand2b_1 _2445_ (.A_N(net85),
    .B(_0921_),
    .Y(_0922_));
 sky130_fd_sc_hd__mux4_1 _2446_ (.A0(\memory[12][1] ),
    .A1(\memory[13][1] ),
    .A2(\memory[14][1] ),
    .A3(\memory[15][1] ),
    .S0(net90),
    .S1(net88),
    .X(_0923_));
 sky130_fd_sc_hd__nand2_1 _2447_ (.A(net85),
    .B(_0923_),
    .Y(_0924_));
 sky130_fd_sc_hd__a32o_1 _2448_ (.A1(_0003_),
    .A2(_0922_),
    .A3(_0924_),
    .B1(_0918_),
    .B2(_0920_),
    .X(_0925_));
 sky130_fd_sc_hd__mux2_1 _2449_ (.A0(_1780_),
    .A1(_0925_),
    .S(_0874_),
    .X(_0926_));
 sky130_fd_sc_hd__mux2_1 _2450_ (.A0(_0926_),
    .A1(net14),
    .S(_0888_),
    .X(_0927_));
 sky130_fd_sc_hd__a21bo_1 _2451_ (.A1(_0462_),
    .A2(_0927_),
    .B1_N(_0916_),
    .X(_0928_));
 sky130_fd_sc_hd__o221a_1 _2452_ (.A1(net400),
    .A2(_0916_),
    .B1(_0928_),
    .B2(_0915_),
    .C1(net113),
    .X(_0005_));
 sky130_fd_sc_hd__a21oi_1 _2453_ (.A1(_0812_),
    .A2(_0813_),
    .B1(_0782_),
    .Y(_0929_));
 sky130_fd_sc_hd__nor2_1 _2454_ (.A(_0783_),
    .B(_0842_),
    .Y(_0930_));
 sky130_fd_sc_hd__mux2_1 _2455_ (.A0(_0850_),
    .A1(_0856_),
    .S(_0847_),
    .X(_0931_));
 sky130_fd_sc_hd__or2_1 _2456_ (.A(_0847_),
    .B(_0854_),
    .X(_0932_));
 sky130_fd_sc_hd__inv_2 _2457_ (.A(_0932_),
    .Y(_0933_));
 sky130_fd_sc_hd__mux2_1 _2458_ (.A0(_0931_),
    .A1(_0933_),
    .S(_0846_),
    .X(_0934_));
 sky130_fd_sc_hd__a21o_1 _2459_ (.A1(_0783_),
    .A2(_0825_),
    .B1(_0798_),
    .X(_0935_));
 sky130_fd_sc_hd__o311a_1 _2460_ (.A1(_0799_),
    .A2(_0929_),
    .A3(_0930_),
    .B1(_0934_),
    .C1(_0935_),
    .X(_0936_));
 sky130_fd_sc_hd__o21bai_1 _2461_ (.A1(net79),
    .A2(_0934_),
    .B1_N(_0936_),
    .Y(_0937_));
 sky130_fd_sc_hd__a21o_1 _2462_ (.A1(net65),
    .A2(_0937_),
    .B1(_0805_),
    .X(_0938_));
 sky130_fd_sc_hd__a211o_1 _2463_ (.A1(_1824_),
    .A2(_0937_),
    .B1(_0805_),
    .C1(_0456_),
    .X(_0939_));
 sky130_fd_sc_hd__nor2_1 _2464_ (.A(_0804_),
    .B(_0861_),
    .Y(_0940_));
 sky130_fd_sc_hd__a211o_1 _2465_ (.A1(_0861_),
    .A2(_0936_),
    .B1(_0940_),
    .C1(_0455_),
    .X(_0941_));
 sky130_fd_sc_hd__o21a_1 _2466_ (.A1(_0871_),
    .A2(_0934_),
    .B1(_0868_),
    .X(_0942_));
 sky130_fd_sc_hd__mux4_1 _2467_ (.A0(\memory[0][2] ),
    .A1(\memory[1][2] ),
    .A2(\memory[2][2] ),
    .A3(\memory[3][2] ),
    .S0(net89),
    .S1(net87),
    .X(_0943_));
 sky130_fd_sc_hd__nand2b_1 _2468_ (.A_N(net85),
    .B(_0943_),
    .Y(_0944_));
 sky130_fd_sc_hd__mux4_1 _2469_ (.A0(\memory[4][2] ),
    .A1(\memory[6][2] ),
    .A2(\memory[5][2] ),
    .A3(\memory[7][2] ),
    .S0(net87),
    .S1(net89),
    .X(_0945_));
 sky130_fd_sc_hd__a21oi_1 _2470_ (.A1(net85),
    .A2(_0945_),
    .B1(_0003_),
    .Y(_0946_));
 sky130_fd_sc_hd__mux4_1 _2471_ (.A0(\memory[8][2] ),
    .A1(\memory[9][2] ),
    .A2(\memory[10][2] ),
    .A3(\memory[11][2] ),
    .S0(net90),
    .S1(_0001_),
    .X(_0947_));
 sky130_fd_sc_hd__nand2b_1 _2472_ (.A_N(net85),
    .B(_0947_),
    .Y(_0948_));
 sky130_fd_sc_hd__mux4_2 _2473_ (.A0(\memory[12][2] ),
    .A1(\memory[13][2] ),
    .A2(\memory[14][2] ),
    .A3(\memory[15][2] ),
    .S0(net90),
    .S1(net88),
    .X(_0949_));
 sky130_fd_sc_hd__nand2_1 _2474_ (.A(net85),
    .B(_0949_),
    .Y(_0950_));
 sky130_fd_sc_hd__a32o_1 _2475_ (.A1(_0003_),
    .A2(_0948_),
    .A3(_0950_),
    .B1(_0944_),
    .B2(_0946_),
    .X(_0951_));
 sky130_fd_sc_hd__mux2_1 _2476_ (.A0(_1779_),
    .A1(_0951_),
    .S(_0874_),
    .X(_0952_));
 sky130_fd_sc_hd__mux2_1 _2477_ (.A0(_0952_),
    .A1(net13),
    .S(_0888_),
    .X(_0953_));
 sky130_fd_sc_hd__a21bo_1 _2478_ (.A1(_0462_),
    .A2(_0953_),
    .B1_N(_0942_),
    .X(_0954_));
 sky130_fd_sc_hd__a31o_1 _2479_ (.A1(_0461_),
    .A2(_0939_),
    .A3(_0941_),
    .B1(_0954_),
    .X(_0955_));
 sky130_fd_sc_hd__o211a_1 _2480_ (.A1(net429),
    .A2(_0942_),
    .B1(_0955_),
    .C1(net113),
    .X(_0006_));
 sky130_fd_sc_hd__a211o_1 _2481_ (.A1(_0777_),
    .A2(_0811_),
    .B1(_0893_),
    .C1(_0782_),
    .X(_0956_));
 sky130_fd_sc_hd__a31oi_1 _2482_ (.A1(_0782_),
    .A2(_0904_),
    .A3(_0905_),
    .B1(_0799_),
    .Y(_0957_));
 sky130_fd_sc_hd__a31o_1 _2483_ (.A1(_1803_),
    .A2(_0780_),
    .A3(_0897_),
    .B1(_0901_),
    .X(_0958_));
 sky130_fd_sc_hd__or2_1 _2484_ (.A(_0847_),
    .B(_0849_),
    .X(_0959_));
 sky130_fd_sc_hd__mux2_1 _2485_ (.A0(_0958_),
    .A1(_0959_),
    .S(_0846_),
    .X(_0960_));
 sky130_fd_sc_hd__o21a_1 _2486_ (.A1(_0782_),
    .A2(_0906_),
    .B1(_0799_),
    .X(_0961_));
 sky130_fd_sc_hd__a211oi_1 _2487_ (.A1(_0956_),
    .A2(_0957_),
    .B1(_0960_),
    .C1(_0961_),
    .Y(_0962_));
 sky130_fd_sc_hd__a21o_1 _2488_ (.A1(net759),
    .A2(_0960_),
    .B1(net61),
    .X(_0963_));
 sky130_fd_sc_hd__o22a_1 _2489_ (.A1(_1820_),
    .A2(net65),
    .B1(_0962_),
    .B2(_0963_),
    .X(_0964_));
 sky130_fd_sc_hd__mux2_1 _2490_ (.A0(_0810_),
    .A1(_0962_),
    .S(_0861_),
    .X(_0965_));
 sky130_fd_sc_hd__or2_1 _2491_ (.A(_0455_),
    .B(_0965_),
    .X(_0966_));
 sky130_fd_sc_hd__o211a_1 _2492_ (.A1(_0456_),
    .A2(_0964_),
    .B1(_0966_),
    .C1(_0461_),
    .X(_0967_));
 sky130_fd_sc_hd__a21oi_1 _2493_ (.A1(_0870_),
    .A2(_0960_),
    .B1(_0869_),
    .Y(_0968_));
 sky130_fd_sc_hd__mux4_1 _2494_ (.A0(\memory[0][3] ),
    .A1(\memory[1][3] ),
    .A2(\memory[2][3] ),
    .A3(\memory[3][3] ),
    .S0(net90),
    .S1(net88),
    .X(_0969_));
 sky130_fd_sc_hd__nand2b_1 _2495_ (.A_N(net86),
    .B(_0969_),
    .Y(_0970_));
 sky130_fd_sc_hd__mux4_1 _2496_ (.A0(\memory[4][3] ),
    .A1(\memory[6][3] ),
    .A2(\memory[5][3] ),
    .A3(\memory[7][3] ),
    .S0(net87),
    .S1(net89),
    .X(_0971_));
 sky130_fd_sc_hd__a21oi_1 _2497_ (.A1(net86),
    .A2(_0971_),
    .B1(_0003_),
    .Y(_0972_));
 sky130_fd_sc_hd__mux4_1 _2498_ (.A0(\memory[8][3] ),
    .A1(\memory[9][3] ),
    .A2(\memory[10][3] ),
    .A3(\memory[11][3] ),
    .S0(net89),
    .S1(net87),
    .X(_0973_));
 sky130_fd_sc_hd__nand2b_1 _2499_ (.A_N(net86),
    .B(_0973_),
    .Y(_0974_));
 sky130_fd_sc_hd__mux4_2 _2500_ (.A0(\memory[12][3] ),
    .A1(\memory[13][3] ),
    .A2(\memory[14][3] ),
    .A3(\memory[15][3] ),
    .S0(net90),
    .S1(net88),
    .X(_0975_));
 sky130_fd_sc_hd__nand2_1 _2501_ (.A(net86),
    .B(_0975_),
    .Y(_0976_));
 sky130_fd_sc_hd__a32o_1 _2502_ (.A1(_0003_),
    .A2(_0974_),
    .A3(_0976_),
    .B1(_0970_),
    .B2(_0972_),
    .X(_0977_));
 sky130_fd_sc_hd__mux2_1 _2503_ (.A0(_1778_),
    .A1(_0977_),
    .S(_0874_),
    .X(_0978_));
 sky130_fd_sc_hd__mux2_1 _2504_ (.A0(_0978_),
    .A1(net12),
    .S(_0888_),
    .X(_0979_));
 sky130_fd_sc_hd__a21bo_1 _2505_ (.A1(_0462_),
    .A2(_0979_),
    .B1_N(_0968_),
    .X(_0980_));
 sky130_fd_sc_hd__o221a_1 _2506_ (.A1(net759),
    .A2(_0968_),
    .B1(_0980_),
    .B2(_0967_),
    .C1(net101),
    .X(_0007_));
 sky130_fd_sc_hd__nand2b_1 _2507_ (.A_N(_0846_),
    .B(_0857_),
    .Y(_0981_));
 sky130_fd_sc_hd__nor3_1 _2508_ (.A(_0799_),
    .B(_0843_),
    .C(_0981_),
    .Y(_0982_));
 sky130_fd_sc_hd__a21o_1 _2509_ (.A1(net730),
    .A2(_0981_),
    .B1(_1823_),
    .X(_0983_));
 sky130_fd_sc_hd__o22a_1 _2510_ (.A1(net65),
    .A2(_0436_),
    .B1(_0982_),
    .B2(_0983_),
    .X(_0984_));
 sky130_fd_sc_hd__mux2_1 _2511_ (.A0(_0839_),
    .A1(_0982_),
    .S(_0861_),
    .X(_0985_));
 sky130_fd_sc_hd__or2_1 _2512_ (.A(_0455_),
    .B(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__o211a_1 _2513_ (.A1(_0456_),
    .A2(_0984_),
    .B1(_0986_),
    .C1(_0461_),
    .X(_0987_));
 sky130_fd_sc_hd__a21oi_1 _2514_ (.A1(_0870_),
    .A2(_0981_),
    .B1(_0869_),
    .Y(_0988_));
 sky130_fd_sc_hd__mux4_1 _2515_ (.A0(\memory[0][4] ),
    .A1(\memory[1][4] ),
    .A2(\memory[2][4] ),
    .A3(\memory[3][4] ),
    .S0(net90),
    .S1(net88),
    .X(_0989_));
 sky130_fd_sc_hd__nand2b_1 _2516_ (.A_N(net86),
    .B(_0989_),
    .Y(_0990_));
 sky130_fd_sc_hd__mux4_1 _2517_ (.A0(\memory[4][4] ),
    .A1(\memory[6][4] ),
    .A2(\memory[5][4] ),
    .A3(\memory[7][4] ),
    .S0(net87),
    .S1(net89),
    .X(_0991_));
 sky130_fd_sc_hd__a21oi_1 _2518_ (.A1(net85),
    .A2(_0991_),
    .B1(_0003_),
    .Y(_0992_));
 sky130_fd_sc_hd__mux4_1 _2519_ (.A0(\memory[8][4] ),
    .A1(\memory[9][4] ),
    .A2(\memory[10][4] ),
    .A3(\memory[11][4] ),
    .S0(net89),
    .S1(net87),
    .X(_0993_));
 sky130_fd_sc_hd__nand2b_1 _2520_ (.A_N(net85),
    .B(_0993_),
    .Y(_0994_));
 sky130_fd_sc_hd__mux4_1 _2521_ (.A0(\memory[12][4] ),
    .A1(\memory[13][4] ),
    .A2(\memory[14][4] ),
    .A3(\memory[15][4] ),
    .S0(net90),
    .S1(net88),
    .X(_0995_));
 sky130_fd_sc_hd__nand2_1 _2522_ (.A(net85),
    .B(_0995_),
    .Y(_0996_));
 sky130_fd_sc_hd__a32o_1 _2523_ (.A1(_0003_),
    .A2(_0994_),
    .A3(_0996_),
    .B1(_0990_),
    .B2(_0992_),
    .X(_0997_));
 sky130_fd_sc_hd__mux2_1 _2524_ (.A0(_1777_),
    .A1(_0997_),
    .S(_0874_),
    .X(_0998_));
 sky130_fd_sc_hd__mux2_1 _2525_ (.A0(_0998_),
    .A1(net11),
    .S(_0888_),
    .X(_0999_));
 sky130_fd_sc_hd__a21bo_1 _2526_ (.A1(_0462_),
    .A2(_0999_),
    .B1_N(_0988_),
    .X(_1000_));
 sky130_fd_sc_hd__o221a_1 _2527_ (.A1(net730),
    .A2(_0988_),
    .B1(_1000_),
    .B2(_0987_),
    .C1(net101),
    .X(_0008_));
 sky130_fd_sc_hd__nor2_1 _2528_ (.A(_0846_),
    .B(_0902_),
    .Y(_1001_));
 sky130_fd_sc_hd__and3b_1 _2529_ (.A_N(_0908_),
    .B(_1001_),
    .C(_0798_),
    .X(_1002_));
 sky130_fd_sc_hd__o21ai_1 _2530_ (.A1(net76),
    .A2(_1001_),
    .B1(net65),
    .Y(_1003_));
 sky130_fd_sc_hd__o22a_1 _2531_ (.A1(net65),
    .A2(_1826_),
    .B1(_1002_),
    .B2(_1003_),
    .X(_1004_));
 sky130_fd_sc_hd__a21o_1 _2532_ (.A1(_0833_),
    .A2(_0862_),
    .B1(_0455_),
    .X(_1005_));
 sky130_fd_sc_hd__a21o_1 _2533_ (.A1(_0861_),
    .A2(_1002_),
    .B1(_1005_),
    .X(_1006_));
 sky130_fd_sc_hd__o211a_1 _2534_ (.A1(_0456_),
    .A2(_1004_),
    .B1(_1006_),
    .C1(_0461_),
    .X(_1007_));
 sky130_fd_sc_hd__o21a_1 _2535_ (.A1(_0871_),
    .A2(_1001_),
    .B1(_0868_),
    .X(_1008_));
 sky130_fd_sc_hd__mux4_1 _2536_ (.A0(\memory[0][5] ),
    .A1(\memory[1][5] ),
    .A2(\memory[2][5] ),
    .A3(\memory[3][5] ),
    .S0(net90),
    .S1(net88),
    .X(_1009_));
 sky130_fd_sc_hd__nand2b_1 _2537_ (.A_N(net86),
    .B(_1009_),
    .Y(_1010_));
 sky130_fd_sc_hd__mux4_1 _2538_ (.A0(\memory[4][5] ),
    .A1(\memory[6][5] ),
    .A2(\memory[5][5] ),
    .A3(\memory[7][5] ),
    .S0(net87),
    .S1(_0000_),
    .X(_1011_));
 sky130_fd_sc_hd__a21oi_1 _2539_ (.A1(net86),
    .A2(_1011_),
    .B1(_0003_),
    .Y(_1012_));
 sky130_fd_sc_hd__mux4_1 _2540_ (.A0(\memory[8][5] ),
    .A1(\memory[9][5] ),
    .A2(\memory[10][5] ),
    .A3(\memory[11][5] ),
    .S0(net89),
    .S1(net87),
    .X(_1013_));
 sky130_fd_sc_hd__nand2b_1 _2541_ (.A_N(net86),
    .B(_1013_),
    .Y(_1014_));
 sky130_fd_sc_hd__mux4_1 _2542_ (.A0(\memory[12][5] ),
    .A1(\memory[13][5] ),
    .A2(\memory[14][5] ),
    .A3(\memory[15][5] ),
    .S0(net90),
    .S1(net88),
    .X(_1015_));
 sky130_fd_sc_hd__nand2_1 _2543_ (.A(net86),
    .B(_1015_),
    .Y(_1016_));
 sky130_fd_sc_hd__a32o_1 _2544_ (.A1(_0003_),
    .A2(_1014_),
    .A3(_1016_),
    .B1(_1010_),
    .B2(_1012_),
    .X(_1017_));
 sky130_fd_sc_hd__mux2_1 _2545_ (.A0(_1776_),
    .A1(_1017_),
    .S(_0874_),
    .X(_1018_));
 sky130_fd_sc_hd__mux2_1 _2546_ (.A0(_1018_),
    .A1(net10),
    .S(_0888_),
    .X(_1019_));
 sky130_fd_sc_hd__a21bo_1 _2547_ (.A1(_0462_),
    .A2(_1019_),
    .B1_N(_1008_),
    .X(_1020_));
 sky130_fd_sc_hd__o221a_1 _2548_ (.A1(net809),
    .A2(_1008_),
    .B1(_1020_),
    .B2(_1007_),
    .C1(net100),
    .X(_0009_));
 sky130_fd_sc_hd__or2_1 _2549_ (.A(_0846_),
    .B(_0932_),
    .X(_1021_));
 sky130_fd_sc_hd__and4b_1 _2550_ (.A_N(_1021_),
    .B(_0825_),
    .C(_0798_),
    .D(_0783_),
    .X(_1022_));
 sky130_fd_sc_hd__and2_1 _2551_ (.A(_0820_),
    .B(_0862_),
    .X(_1023_));
 sky130_fd_sc_hd__a21o_1 _2552_ (.A1(net641),
    .A2(_1021_),
    .B1(_1823_),
    .X(_1024_));
 sky130_fd_sc_hd__o22a_1 _2553_ (.A1(_1804_),
    .A2(net65),
    .B1(_1022_),
    .B2(_1024_),
    .X(_1025_));
 sky130_fd_sc_hd__a211o_1 _2554_ (.A1(_0861_),
    .A2(_1022_),
    .B1(_1023_),
    .C1(_0455_),
    .X(_1026_));
 sky130_fd_sc_hd__o211a_1 _2555_ (.A1(_0456_),
    .A2(_1025_),
    .B1(_1026_),
    .C1(_0461_),
    .X(_1027_));
 sky130_fd_sc_hd__a21oi_1 _2556_ (.A1(_0870_),
    .A2(_1021_),
    .B1(_0869_),
    .Y(_1028_));
 sky130_fd_sc_hd__mux4_1 _2557_ (.A0(\memory[0][6] ),
    .A1(\memory[1][6] ),
    .A2(\memory[2][6] ),
    .A3(\memory[3][6] ),
    .S0(net90),
    .S1(net88),
    .X(_1029_));
 sky130_fd_sc_hd__nand2b_1 _2558_ (.A_N(net86),
    .B(_1029_),
    .Y(_1030_));
 sky130_fd_sc_hd__mux4_1 _2559_ (.A0(\memory[4][6] ),
    .A1(\memory[6][6] ),
    .A2(\memory[5][6] ),
    .A3(\memory[7][6] ),
    .S0(net87),
    .S1(net89),
    .X(_1031_));
 sky130_fd_sc_hd__a21oi_1 _2560_ (.A1(net85),
    .A2(_1031_),
    .B1(_0003_),
    .Y(_1032_));
 sky130_fd_sc_hd__mux4_1 _2561_ (.A0(\memory[8][6] ),
    .A1(\memory[9][6] ),
    .A2(\memory[10][6] ),
    .A3(\memory[11][6] ),
    .S0(net89),
    .S1(net87),
    .X(_1033_));
 sky130_fd_sc_hd__nand2b_1 _2562_ (.A_N(_0002_),
    .B(_1033_),
    .Y(_1034_));
 sky130_fd_sc_hd__mux4_1 _2563_ (.A0(\memory[12][6] ),
    .A1(\memory[13][6] ),
    .A2(\memory[14][6] ),
    .A3(\memory[15][6] ),
    .S0(net90),
    .S1(net88),
    .X(_1035_));
 sky130_fd_sc_hd__nand2_1 _2564_ (.A(net86),
    .B(_1035_),
    .Y(_1036_));
 sky130_fd_sc_hd__a32o_1 _2565_ (.A1(_0003_),
    .A2(_1034_),
    .A3(_1036_),
    .B1(_1030_),
    .B2(_1032_),
    .X(_1037_));
 sky130_fd_sc_hd__mux2_1 _2566_ (.A0(_1775_),
    .A1(_1037_),
    .S(_0874_),
    .X(_1038_));
 sky130_fd_sc_hd__mux2_1 _2567_ (.A0(_1038_),
    .A1(net9),
    .S(_0888_),
    .X(_1039_));
 sky130_fd_sc_hd__a21bo_1 _2568_ (.A1(_0462_),
    .A2(_1039_),
    .B1_N(_1028_),
    .X(_1040_));
 sky130_fd_sc_hd__o221a_1 _2569_ (.A1(net641),
    .A2(_1028_),
    .B1(_1040_),
    .B2(_1027_),
    .C1(net101),
    .X(_0010_));
 sky130_fd_sc_hd__nor2_1 _2570_ (.A(_0846_),
    .B(_0959_),
    .Y(_1041_));
 sky130_fd_sc_hd__and4_1 _2571_ (.A(_0777_),
    .B(_0783_),
    .C(_0798_),
    .D(_0824_),
    .X(_1042_));
 sky130_fd_sc_hd__mux2_1 _2572_ (.A0(net680),
    .A1(_1042_),
    .S(_1041_),
    .X(_1043_));
 sky130_fd_sc_hd__mux2_1 _2573_ (.A0(_1807_),
    .A1(_1043_),
    .S(net65),
    .X(_1044_));
 sky130_fd_sc_hd__a21o_1 _2574_ (.A1(_0823_),
    .A2(_0862_),
    .B1(_0455_),
    .X(_1045_));
 sky130_fd_sc_hd__a31o_1 _2575_ (.A1(_0861_),
    .A2(_1041_),
    .A3(_1042_),
    .B1(_1045_),
    .X(_1046_));
 sky130_fd_sc_hd__o211a_1 _2576_ (.A1(_0456_),
    .A2(_1044_),
    .B1(_1046_),
    .C1(_0461_),
    .X(_1047_));
 sky130_fd_sc_hd__o21a_1 _2577_ (.A1(_0871_),
    .A2(_1041_),
    .B1(_0868_),
    .X(_1048_));
 sky130_fd_sc_hd__mux4_1 _2578_ (.A0(\memory[0][7] ),
    .A1(\memory[1][7] ),
    .A2(\memory[2][7] ),
    .A3(\memory[3][7] ),
    .S0(net89),
    .S1(net87),
    .X(_1049_));
 sky130_fd_sc_hd__nand2b_1 _2579_ (.A_N(net85),
    .B(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__mux4_1 _2580_ (.A0(\memory[4][7] ),
    .A1(\memory[6][7] ),
    .A2(\memory[5][7] ),
    .A3(\memory[7][7] ),
    .S0(net88),
    .S1(net89),
    .X(_1051_));
 sky130_fd_sc_hd__a21oi_1 _2581_ (.A1(net85),
    .A2(_1051_),
    .B1(_0003_),
    .Y(_1052_));
 sky130_fd_sc_hd__mux4_1 _2582_ (.A0(\memory[8][7] ),
    .A1(\memory[9][7] ),
    .A2(\memory[10][7] ),
    .A3(\memory[11][7] ),
    .S0(net89),
    .S1(net87),
    .X(_1053_));
 sky130_fd_sc_hd__nand2b_1 _2583_ (.A_N(net85),
    .B(_1053_),
    .Y(_1054_));
 sky130_fd_sc_hd__mux4_2 _2584_ (.A0(\memory[12][7] ),
    .A1(\memory[13][7] ),
    .A2(\memory[14][7] ),
    .A3(\memory[15][7] ),
    .S0(net90),
    .S1(net88),
    .X(_1055_));
 sky130_fd_sc_hd__nand2_1 _2585_ (.A(net85),
    .B(_1055_),
    .Y(_1056_));
 sky130_fd_sc_hd__a32o_1 _2586_ (.A1(_0003_),
    .A2(_1054_),
    .A3(_1056_),
    .B1(_1050_),
    .B2(_1052_),
    .X(_1057_));
 sky130_fd_sc_hd__mux2_1 _2587_ (.A0(_1774_),
    .A1(_1057_),
    .S(_0874_),
    .X(_1058_));
 sky130_fd_sc_hd__mux2_1 _2588_ (.A0(_1058_),
    .A1(net8),
    .S(_0888_),
    .X(_1059_));
 sky130_fd_sc_hd__a21bo_1 _2589_ (.A1(_0462_),
    .A2(_1059_),
    .B1_N(_1048_),
    .X(_1060_));
 sky130_fd_sc_hd__o221a_1 _2590_ (.A1(net680),
    .A2(_1048_),
    .B1(_1060_),
    .B2(_1047_),
    .C1(net101),
    .X(_0011_));
 sky130_fd_sc_hd__nor2_1 _2591_ (.A(_1782_),
    .B(net31),
    .Y(_1061_));
 sky130_fd_sc_hd__or4b_2 _2592_ (.A(_1782_),
    .B(_0873_),
    .C(net31),
    .D_N(net34),
    .X(_1062_));
 sky130_fd_sc_hd__nand2_1 _2593_ (.A(\cmdr[3] ),
    .B(\cmdr[2] ),
    .Y(_1063_));
 sky130_fd_sc_hd__or2_2 _2594_ (.A(_1062_),
    .B(_1063_),
    .X(_1064_));
 sky130_fd_sc_hd__or3b_4 _2595_ (.A(\cmdr[0] ),
    .B(_1064_),
    .C_N(\cmdr[1] ),
    .X(_1065_));
 sky130_fd_sc_hd__mux2_1 _2596_ (.A0(net81),
    .A1(net374),
    .S(_1065_),
    .X(_0012_));
 sky130_fd_sc_hd__mux2_1 _2597_ (.A0(net80),
    .A1(net338),
    .S(_1065_),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_1 _2598_ (.A0(net79),
    .A1(net310),
    .S(_1065_),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _2599_ (.A0(net78),
    .A1(net376),
    .S(_1065_),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _2600_ (.A0(net77),
    .A1(net362),
    .S(_1065_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _2601_ (.A0(net76),
    .A1(net300),
    .S(_1065_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _2602_ (.A0(net75),
    .A1(net302),
    .S(_1065_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _2603_ (.A0(net74),
    .A1(net322),
    .S(_1065_),
    .X(_0019_));
 sky130_fd_sc_hd__or4_1 _2604_ (.A(_0721_),
    .B(_0732_),
    .C(_0748_),
    .D(_0754_),
    .X(_1066_));
 sky130_fd_sc_hd__o41a_1 _2605_ (.A1(_0506_),
    .A2(_0543_),
    .A3(_0561_),
    .A4(_0755_),
    .B1(_1066_),
    .X(_1067_));
 sky130_fd_sc_hd__nand3_1 _2606_ (.A(_0651_),
    .B(_0680_),
    .C(_0694_),
    .Y(_1068_));
 sky130_fd_sc_hd__or4_1 _2607_ (.A(_0588_),
    .B(_0606_),
    .C(_0624_),
    .D(_0642_),
    .X(_1069_));
 sky130_fd_sc_hd__o22a_1 _2608_ (.A1(_0709_),
    .A2(_1068_),
    .B1(_1069_),
    .B2(net65),
    .X(_1070_));
 sky130_fd_sc_hd__or2_1 _2609_ (.A(_1067_),
    .B(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__and3_2 _2610_ (.A(_1792_),
    .B(_0658_),
    .C(_1071_),
    .X(_1072_));
 sky130_fd_sc_hd__nand2_1 _2611_ (.A(net599),
    .B(net84),
    .Y(_1073_));
 sky130_fd_sc_hd__nand2_1 _2612_ (.A(net599),
    .B(_0461_),
    .Y(_1074_));
 sky130_fd_sc_hd__nor2_2 _2613_ (.A(_0465_),
    .B(_1074_),
    .Y(_1075_));
 sky130_fd_sc_hd__or2_2 _2614_ (.A(_0465_),
    .B(_1074_),
    .X(_1076_));
 sky130_fd_sc_hd__nor2_2 _2615_ (.A(_1072_),
    .B(_1076_),
    .Y(_1077_));
 sky130_fd_sc_hd__or3_4 _2616_ (.A(_1787_),
    .B(_1791_),
    .C(_1797_),
    .X(_1078_));
 sky130_fd_sc_hd__nand2b_4 _2617_ (.A_N(_1072_),
    .B(_1078_),
    .Y(_1079_));
 sky130_fd_sc_hd__inv_2 _2618_ (.A(_1079_),
    .Y(_1080_));
 sky130_fd_sc_hd__and3_2 _2619_ (.A(net470),
    .B(net801),
    .C(net740),
    .X(_1081_));
 sky130_fd_sc_hd__nand2_1 _2620_ (.A(net750),
    .B(_1081_),
    .Y(_1082_));
 sky130_fd_sc_hd__nand3_1 _2621_ (.A(net742),
    .B(net750),
    .C(_1081_),
    .Y(_1083_));
 sky130_fd_sc_hd__and4_1 _2622_ (.A(\S8x305.PC[4] ),
    .B(\S8x305.PC[3] ),
    .C(\S8x305.PC[5] ),
    .D(_1081_),
    .X(_1084_));
 sky130_fd_sc_hd__and2_1 _2623_ (.A(\S8x305.PC[6] ),
    .B(_1084_),
    .X(_1085_));
 sky130_fd_sc_hd__and3_1 _2624_ (.A(net463),
    .B(net737),
    .C(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__a21oi_1 _2625_ (.A1(net472),
    .A2(_1085_),
    .B1(net463),
    .Y(_1087_));
 sky130_fd_sc_hd__o32a_1 _2626_ (.A1(_1079_),
    .A2(net464),
    .A3(net473),
    .B1(_1078_),
    .B2(_1811_),
    .X(_1088_));
 sky130_fd_sc_hd__nand2_1 _2627_ (.A(_1077_),
    .B(net474),
    .Y(_1089_));
 sky130_fd_sc_hd__o211a_1 _2628_ (.A1(net463),
    .A2(_1077_),
    .B1(_1089_),
    .C1(net103),
    .X(_0020_));
 sky130_fd_sc_hd__and2_1 _2629_ (.A(net441),
    .B(_1086_),
    .X(_1090_));
 sky130_fd_sc_hd__nor2_1 _2630_ (.A(net441),
    .B(net464),
    .Y(_1091_));
 sky130_fd_sc_hd__o32a_1 _2631_ (.A1(_1079_),
    .A2(_1090_),
    .A3(_1091_),
    .B1(_1078_),
    .B2(net62),
    .X(_1092_));
 sky130_fd_sc_hd__nand2_1 _2632_ (.A(_1077_),
    .B(net465),
    .Y(_1093_));
 sky130_fd_sc_hd__o211a_1 _2633_ (.A1(net441),
    .A2(_1077_),
    .B1(_1093_),
    .C1(net103),
    .X(_0021_));
 sky130_fd_sc_hd__xnor2_1 _2634_ (.A(net556),
    .B(_1090_),
    .Y(_1094_));
 sky130_fd_sc_hd__o221ai_1 _2635_ (.A1(_1828_),
    .A2(_1078_),
    .B1(_1079_),
    .B2(_1094_),
    .C1(_1077_),
    .Y(_1095_));
 sky130_fd_sc_hd__o211a_1 _2636_ (.A1(net556),
    .A2(_1077_),
    .B1(_1095_),
    .C1(net103),
    .X(_0022_));
 sky130_fd_sc_hd__and3_1 _2637_ (.A(net122),
    .B(net556),
    .C(_1090_),
    .X(_1096_));
 sky130_fd_sc_hd__a21oi_1 _2638_ (.A1(net556),
    .A2(_1090_),
    .B1(net122),
    .Y(_1097_));
 sky130_fd_sc_hd__o32ai_1 _2639_ (.A1(_1079_),
    .A2(_1096_),
    .A3(_1097_),
    .B1(_1078_),
    .B2(_0435_),
    .Y(_1098_));
 sky130_fd_sc_hd__or2_1 _2640_ (.A(net122),
    .B(_1077_),
    .X(_1099_));
 sky130_fd_sc_hd__o311a_1 _2641_ (.A1(_1072_),
    .A2(_1076_),
    .A3(_1098_),
    .B1(_1099_),
    .C1(net103),
    .X(_0023_));
 sky130_fd_sc_hd__xnor2_1 _2642_ (.A(net445),
    .B(_1096_),
    .Y(_1100_));
 sky130_fd_sc_hd__o221a_1 _2643_ (.A1(net61),
    .A2(_1078_),
    .B1(_1079_),
    .B2(_1100_),
    .C1(_1077_),
    .X(_1101_));
 sky130_fd_sc_hd__o21ai_1 _2644_ (.A1(net445),
    .A2(_1077_),
    .B1(net103),
    .Y(_1102_));
 sky130_fd_sc_hd__nor2_1 _2645_ (.A(_1101_),
    .B(_1102_),
    .Y(_0024_));
 sky130_fd_sc_hd__or4_4 _2646_ (.A(_1771_),
    .B(_1799_),
    .C(net66),
    .D(_0487_),
    .X(_1103_));
 sky130_fd_sc_hd__nor2_8 _2647_ (.A(_0443_),
    .B(_1103_),
    .Y(_1104_));
 sky130_fd_sc_hd__inv_2 _2648_ (.A(_1104_),
    .Y(_1105_));
 sky130_fd_sc_hd__a21oi_2 _2649_ (.A1(_1825_),
    .A2(_0488_),
    .B1(_1104_),
    .Y(_1106_));
 sky130_fd_sc_hd__a21o_1 _2650_ (.A1(_1825_),
    .A2(_0488_),
    .B1(_1104_),
    .X(_1107_));
 sky130_fd_sc_hd__or3b_4 _2651_ (.A(_0437_),
    .B(_1106_),
    .C_N(_1830_),
    .X(_1108_));
 sky130_fd_sc_hd__nor2_2 _2652_ (.A(_0445_),
    .B(_1108_),
    .Y(_1109_));
 sky130_fd_sc_hd__or2_2 _2653_ (.A(_0445_),
    .B(_1108_),
    .X(_1110_));
 sky130_fd_sc_hd__and3_1 _2654_ (.A(net107),
    .B(net622),
    .C(_1110_),
    .X(_1111_));
 sky130_fd_sc_hd__mux2_8 _2655_ (.A0(_0823_),
    .A1(_1044_),
    .S(_1104_),
    .X(_1112_));
 sky130_fd_sc_hd__a21o_1 _2656_ (.A1(_1109_),
    .A2(_1112_),
    .B1(_1111_),
    .X(_0025_));
 sky130_fd_sc_hd__and3_1 _2657_ (.A(net109),
    .B(net613),
    .C(_1110_),
    .X(_1113_));
 sky130_fd_sc_hd__mux2_8 _2658_ (.A0(_0820_),
    .A1(_1025_),
    .S(_1104_),
    .X(_1114_));
 sky130_fd_sc_hd__a21o_1 _2659_ (.A1(_1109_),
    .A2(_1114_),
    .B1(_1113_),
    .X(_0026_));
 sky130_fd_sc_hd__and3_1 _2660_ (.A(net107),
    .B(net566),
    .C(_1110_),
    .X(_1115_));
 sky130_fd_sc_hd__mux2_8 _2661_ (.A0(_0833_),
    .A1(_1004_),
    .S(_1104_),
    .X(_1116_));
 sky130_fd_sc_hd__a21o_1 _2662_ (.A1(_1109_),
    .A2(_1116_),
    .B1(_1115_),
    .X(_0027_));
 sky130_fd_sc_hd__and3_1 _2663_ (.A(net107),
    .B(net586),
    .C(_1110_),
    .X(_1117_));
 sky130_fd_sc_hd__mux2_8 _2664_ (.A0(_0839_),
    .A1(_0984_),
    .S(_1104_),
    .X(_1118_));
 sky130_fd_sc_hd__a21o_1 _2665_ (.A1(_1109_),
    .A2(_1118_),
    .B1(_1117_),
    .X(_0028_));
 sky130_fd_sc_hd__and3_1 _2666_ (.A(net109),
    .B(net628),
    .C(_1110_),
    .X(_1119_));
 sky130_fd_sc_hd__mux2_8 _2667_ (.A0(_0810_),
    .A1(_0964_),
    .S(_1104_),
    .X(_1120_));
 sky130_fd_sc_hd__a21o_1 _2668_ (.A1(_1109_),
    .A2(_1120_),
    .B1(_1119_),
    .X(_0029_));
 sky130_fd_sc_hd__and3_1 _2669_ (.A(net110),
    .B(net492),
    .C(_1110_),
    .X(_1121_));
 sky130_fd_sc_hd__nor2_1 _2670_ (.A(_0804_),
    .B(_1104_),
    .Y(_1122_));
 sky130_fd_sc_hd__a21o_4 _2671_ (.A1(_0938_),
    .A2(_1104_),
    .B1(_1122_),
    .X(_1123_));
 sky130_fd_sc_hd__a21o_1 _2672_ (.A1(_1109_),
    .A2(_1123_),
    .B1(_1121_),
    .X(_0030_));
 sky130_fd_sc_hd__and3_1 _2673_ (.A(net108),
    .B(net548),
    .C(_1110_),
    .X(_1124_));
 sky130_fd_sc_hd__mux2_8 _2674_ (.A0(_0791_),
    .A1(_0911_),
    .S(_1104_),
    .X(_1125_));
 sky130_fd_sc_hd__a21o_1 _2675_ (.A1(_1109_),
    .A2(_1125_),
    .B1(_1124_),
    .X(_0031_));
 sky130_fd_sc_hd__and3_1 _2676_ (.A(net108),
    .B(net498),
    .C(_1110_),
    .X(_1126_));
 sky130_fd_sc_hd__or2_1 _2677_ (.A(_0772_),
    .B(_1104_),
    .X(_1127_));
 sky130_fd_sc_hd__o31a_4 _2678_ (.A1(_0460_),
    .A2(_0860_),
    .A3(_1105_),
    .B1(_1127_),
    .X(_1128_));
 sky130_fd_sc_hd__a21o_1 _2679_ (.A1(_1109_),
    .A2(_1128_),
    .B1(_1126_),
    .X(_0032_));
 sky130_fd_sc_hd__and2_2 _2680_ (.A(_1836_),
    .B(_1061_),
    .X(_1129_));
 sky130_fd_sc_hd__nand2_4 _2681_ (.A(_1836_),
    .B(_1061_),
    .Y(_1130_));
 sky130_fd_sc_hd__or2_1 _2682_ (.A(net690),
    .B(_1129_),
    .X(_1131_));
 sky130_fd_sc_hd__o211a_1 _2683_ (.A1(net680),
    .A2(_1130_),
    .B1(_1131_),
    .C1(net99),
    .X(_0033_));
 sky130_fd_sc_hd__or2_1 _2684_ (.A(net666),
    .B(_1129_),
    .X(_1132_));
 sky130_fd_sc_hd__o211a_1 _2685_ (.A1(net641),
    .A2(_1130_),
    .B1(_1132_),
    .C1(net99),
    .X(_0034_));
 sky130_fd_sc_hd__or2_1 _2686_ (.A(net811),
    .B(_1129_),
    .X(_1133_));
 sky130_fd_sc_hd__o211a_1 _2687_ (.A1(net809),
    .A2(_1130_),
    .B1(_1133_),
    .C1(net99),
    .X(_0035_));
 sky130_fd_sc_hd__or2_1 _2688_ (.A(net734),
    .B(_1129_),
    .X(_1134_));
 sky130_fd_sc_hd__o211a_1 _2689_ (.A1(net730),
    .A2(_1130_),
    .B1(_1134_),
    .C1(net99),
    .X(_0036_));
 sky130_fd_sc_hd__nor2_2 _2690_ (.A(_1817_),
    .B(_1108_),
    .Y(_1135_));
 sky130_fd_sc_hd__or2_2 _2691_ (.A(_1817_),
    .B(_1108_),
    .X(_1136_));
 sky130_fd_sc_hd__and3_1 _2692_ (.A(net107),
    .B(net577),
    .C(_1136_),
    .X(_1137_));
 sky130_fd_sc_hd__a21o_1 _2693_ (.A1(_1112_),
    .A2(_1135_),
    .B1(_1137_),
    .X(_0037_));
 sky130_fd_sc_hd__and3_1 _2694_ (.A(net109),
    .B(net619),
    .C(_1136_),
    .X(_1138_));
 sky130_fd_sc_hd__a21o_1 _2695_ (.A1(_1114_),
    .A2(_1135_),
    .B1(_1138_),
    .X(_0038_));
 sky130_fd_sc_hd__and3_1 _2696_ (.A(net113),
    .B(net537),
    .C(_1136_),
    .X(_1139_));
 sky130_fd_sc_hd__a21o_1 _2697_ (.A1(_1116_),
    .A2(_1135_),
    .B1(_1139_),
    .X(_0039_));
 sky130_fd_sc_hd__and3_1 _2698_ (.A(net113),
    .B(net590),
    .C(_1136_),
    .X(_1140_));
 sky130_fd_sc_hd__a21o_1 _2699_ (.A1(_1118_),
    .A2(_1135_),
    .B1(_1140_),
    .X(_0040_));
 sky130_fd_sc_hd__and3_1 _2700_ (.A(net109),
    .B(net598),
    .C(_1136_),
    .X(_1141_));
 sky130_fd_sc_hd__a21o_1 _2701_ (.A1(_1120_),
    .A2(_1135_),
    .B1(_1141_),
    .X(_0041_));
 sky130_fd_sc_hd__and3_1 _2702_ (.A(net110),
    .B(net652),
    .C(_1136_),
    .X(_1142_));
 sky130_fd_sc_hd__a21o_1 _2703_ (.A1(_1123_),
    .A2(_1135_),
    .B1(_1142_),
    .X(_0042_));
 sky130_fd_sc_hd__and3_1 _2704_ (.A(net108),
    .B(net539),
    .C(_1136_),
    .X(_1143_));
 sky130_fd_sc_hd__a21o_1 _2705_ (.A1(_1125_),
    .A2(_1135_),
    .B1(_1143_),
    .X(_0043_));
 sky130_fd_sc_hd__and3_1 _2706_ (.A(net108),
    .B(net615),
    .C(_1136_),
    .X(_1144_));
 sky130_fd_sc_hd__a21o_1 _2707_ (.A1(_1128_),
    .A2(_1135_),
    .B1(_1144_),
    .X(_0044_));
 sky130_fd_sc_hd__nor2_2 _2708_ (.A(net40),
    .B(net92),
    .Y(_1145_));
 sky130_fd_sc_hd__nor2_2 _2709_ (.A(_1806_),
    .B(_1814_),
    .Y(_1146_));
 sky130_fd_sc_hd__or2_1 _2710_ (.A(_1806_),
    .B(_1814_),
    .X(_1147_));
 sky130_fd_sc_hd__and3b_2 _2711_ (.A_N(_1830_),
    .B(_0437_),
    .C(_1107_),
    .X(_1148_));
 sky130_fd_sc_hd__and2_2 _2712_ (.A(_1146_),
    .B(_1148_),
    .X(_1149_));
 sky130_fd_sc_hd__a22o_1 _2713_ (.A1(net168),
    .A2(_1145_),
    .B1(_1149_),
    .B2(_1114_),
    .X(_0045_));
 sky130_fd_sc_hd__a22o_1 _2714_ (.A1(net146),
    .A2(_1145_),
    .B1(_1149_),
    .B2(_1116_),
    .X(_0046_));
 sky130_fd_sc_hd__a22o_1 _2715_ (.A1(net152),
    .A2(_1145_),
    .B1(_1149_),
    .B2(_1118_),
    .X(_0047_));
 sky130_fd_sc_hd__a22o_1 _2716_ (.A1(net140),
    .A2(_1145_),
    .B1(_1149_),
    .B2(_1120_),
    .X(_0048_));
 sky130_fd_sc_hd__a22o_1 _2717_ (.A1(net208),
    .A2(_1145_),
    .B1(_1149_),
    .B2(_1123_),
    .X(_0049_));
 sky130_fd_sc_hd__a22o_1 _2718_ (.A1(net128),
    .A2(_1145_),
    .B1(_1149_),
    .B2(_1125_),
    .X(_0050_));
 sky130_fd_sc_hd__a22o_1 _2719_ (.A1(net156),
    .A2(_1145_),
    .B1(_1149_),
    .B2(_1128_),
    .X(_0051_));
 sky130_fd_sc_hd__xnor2_1 _2720_ (.A(net729),
    .B(_1083_),
    .Y(_1150_));
 sky130_fd_sc_hd__mux2_1 _2721_ (.A0(_1150_),
    .A1(_0805_),
    .S(_1072_),
    .X(_1151_));
 sky130_fd_sc_hd__a21oi_2 _2722_ (.A1(net66),
    .A2(_1072_),
    .B1(_1076_),
    .Y(_1152_));
 sky130_fd_sc_hd__mux2_1 _2723_ (.A0(_0474_),
    .A1(_1151_),
    .S(_1078_),
    .X(_1153_));
 sky130_fd_sc_hd__mux2_1 _2724_ (.A0(net729),
    .A1(_1153_),
    .S(_1152_),
    .X(_1154_));
 sky130_fd_sc_hd__and2_1 _2725_ (.A(net104),
    .B(_1154_),
    .X(_0052_));
 sky130_fd_sc_hd__nor2_1 _2726_ (.A(\S8x305.PC[6] ),
    .B(_1084_),
    .Y(_1155_));
 sky130_fd_sc_hd__or3_1 _2727_ (.A(_1072_),
    .B(_1085_),
    .C(_1155_),
    .X(_1156_));
 sky130_fd_sc_hd__a21bo_1 _2728_ (.A1(_0793_),
    .A2(_1072_),
    .B1_N(_1156_),
    .X(_1157_));
 sky130_fd_sc_hd__mux2_1 _2729_ (.A0(_0469_),
    .A1(_1157_),
    .S(_1078_),
    .X(_1158_));
 sky130_fd_sc_hd__mux2_1 _2730_ (.A0(net800),
    .A1(_1158_),
    .S(_1152_),
    .X(_1159_));
 sky130_fd_sc_hd__and2_1 _2731_ (.A(net104),
    .B(_1159_),
    .X(_0053_));
 sky130_fd_sc_hd__xor2_1 _2732_ (.A(net472),
    .B(_1085_),
    .X(_1160_));
 sky130_fd_sc_hd__mux2_1 _2733_ (.A0(_1160_),
    .A1(_0460_),
    .S(_1072_),
    .X(_1161_));
 sky130_fd_sc_hd__mux2_1 _2734_ (.A0(_0459_),
    .A1(_1161_),
    .S(_1078_),
    .X(_1162_));
 sky130_fd_sc_hd__mux2_1 _2735_ (.A0(net472),
    .A1(_1162_),
    .S(_1152_),
    .X(_1163_));
 sky130_fd_sc_hd__and2_1 _2736_ (.A(net104),
    .B(_1163_),
    .X(_0054_));
 sky130_fd_sc_hd__and3_1 _2737_ (.A(net459),
    .B(_0488_),
    .C(_0658_),
    .X(_1164_));
 sky130_fd_sc_hd__and2_1 _2738_ (.A(net104),
    .B(net825),
    .X(_1165_));
 sky130_fd_sc_hd__o21a_1 _2739_ (.A1(_0655_),
    .A2(_0768_),
    .B1(_0656_),
    .X(_1166_));
 sky130_fd_sc_hd__mux2_1 _2740_ (.A0(_1165_),
    .A1(_1166_),
    .S(_1164_),
    .X(_1167_));
 sky130_fd_sc_hd__mux2_1 _2741_ (.A0(_1167_),
    .A1(_1112_),
    .S(_1149_),
    .X(_0055_));
 sky130_fd_sc_hd__and2_2 _2742_ (.A(_0444_),
    .B(_1148_),
    .X(_1168_));
 sky130_fd_sc_hd__nand2_2 _2743_ (.A(_0444_),
    .B(_1148_),
    .Y(_1169_));
 sky130_fd_sc_hd__and3_1 _2744_ (.A(net108),
    .B(net573),
    .C(_1169_),
    .X(_1170_));
 sky130_fd_sc_hd__a21o_1 _2745_ (.A1(_1112_),
    .A2(_1168_),
    .B1(_1170_),
    .X(_0056_));
 sky130_fd_sc_hd__and3_1 _2746_ (.A(net105),
    .B(net528),
    .C(_1169_),
    .X(_1171_));
 sky130_fd_sc_hd__a21o_1 _2747_ (.A1(_1114_),
    .A2(_1168_),
    .B1(_1171_),
    .X(_0057_));
 sky130_fd_sc_hd__and3_1 _2748_ (.A(net105),
    .B(net493),
    .C(_1169_),
    .X(_1172_));
 sky130_fd_sc_hd__a21o_1 _2749_ (.A1(_1116_),
    .A2(_1168_),
    .B1(_1172_),
    .X(_0058_));
 sky130_fd_sc_hd__and3_1 _2750_ (.A(net105),
    .B(net636),
    .C(_1169_),
    .X(_1173_));
 sky130_fd_sc_hd__a21o_1 _2751_ (.A1(_1118_),
    .A2(_1168_),
    .B1(_1173_),
    .X(_0059_));
 sky130_fd_sc_hd__and3_1 _2752_ (.A(net105),
    .B(net630),
    .C(_1169_),
    .X(_1174_));
 sky130_fd_sc_hd__a21o_1 _2753_ (.A1(_1120_),
    .A2(_1168_),
    .B1(_1174_),
    .X(_0060_));
 sky130_fd_sc_hd__and3_1 _2754_ (.A(net108),
    .B(net563),
    .C(_1169_),
    .X(_1175_));
 sky130_fd_sc_hd__a21o_1 _2755_ (.A1(_1123_),
    .A2(_1168_),
    .B1(_1175_),
    .X(_0061_));
 sky130_fd_sc_hd__and3_1 _2756_ (.A(net108),
    .B(net596),
    .C(_1169_),
    .X(_1176_));
 sky130_fd_sc_hd__a21o_1 _2757_ (.A1(_1125_),
    .A2(_1168_),
    .B1(_1176_),
    .X(_0062_));
 sky130_fd_sc_hd__and3_1 _2758_ (.A(net108),
    .B(net507),
    .C(_1169_),
    .X(_1177_));
 sky130_fd_sc_hd__a21o_1 _2759_ (.A1(_1128_),
    .A2(_1168_),
    .B1(_1177_),
    .X(_0063_));
 sky130_fd_sc_hd__and3_2 _2760_ (.A(_1830_),
    .B(_0437_),
    .C(_1107_),
    .X(_1178_));
 sky130_fd_sc_hd__and2_2 _2761_ (.A(_1816_),
    .B(_1178_),
    .X(_1179_));
 sky130_fd_sc_hd__nand2_2 _2762_ (.A(_1816_),
    .B(_1178_),
    .Y(_1180_));
 sky130_fd_sc_hd__and3_1 _2763_ (.A(net108),
    .B(net646),
    .C(_1180_),
    .X(_1181_));
 sky130_fd_sc_hd__a21o_1 _2764_ (.A1(_1112_),
    .A2(_1179_),
    .B1(_1181_),
    .X(_0064_));
 sky130_fd_sc_hd__and3_1 _2765_ (.A(net105),
    .B(net568),
    .C(_1180_),
    .X(_1182_));
 sky130_fd_sc_hd__a21o_1 _2766_ (.A1(_1114_),
    .A2(_1179_),
    .B1(_1182_),
    .X(_0065_));
 sky130_fd_sc_hd__and3_1 _2767_ (.A(net105),
    .B(net534),
    .C(_1180_),
    .X(_1183_));
 sky130_fd_sc_hd__a21o_1 _2768_ (.A1(_1116_),
    .A2(_1179_),
    .B1(_1183_),
    .X(_0066_));
 sky130_fd_sc_hd__and3_1 _2769_ (.A(net105),
    .B(net571),
    .C(_1180_),
    .X(_1184_));
 sky130_fd_sc_hd__a21o_1 _2770_ (.A1(_1118_),
    .A2(_1179_),
    .B1(_1184_),
    .X(_0067_));
 sky130_fd_sc_hd__and3_1 _2771_ (.A(net105),
    .B(net651),
    .C(_1180_),
    .X(_1185_));
 sky130_fd_sc_hd__a21o_1 _2772_ (.A1(_1120_),
    .A2(_1179_),
    .B1(_1185_),
    .X(_0068_));
 sky130_fd_sc_hd__and3_1 _2773_ (.A(net107),
    .B(net635),
    .C(_1180_),
    .X(_1186_));
 sky130_fd_sc_hd__a21o_1 _2774_ (.A1(_1123_),
    .A2(_1179_),
    .B1(_1186_),
    .X(_0069_));
 sky130_fd_sc_hd__and3_1 _2775_ (.A(net107),
    .B(net591),
    .C(_1180_),
    .X(_1187_));
 sky130_fd_sc_hd__a21o_1 _2776_ (.A1(_1125_),
    .A2(_1179_),
    .B1(_1187_),
    .X(_0070_));
 sky130_fd_sc_hd__and3_1 _2777_ (.A(net108),
    .B(net602),
    .C(_1180_),
    .X(_1188_));
 sky130_fd_sc_hd__a21o_1 _2778_ (.A1(_1128_),
    .A2(_1179_),
    .B1(_1188_),
    .X(_0071_));
 sky130_fd_sc_hd__and2_2 _2779_ (.A(_1816_),
    .B(_1148_),
    .X(_1189_));
 sky130_fd_sc_hd__nand2_2 _2780_ (.A(_1816_),
    .B(_1148_),
    .Y(_1190_));
 sky130_fd_sc_hd__and3_1 _2781_ (.A(net108),
    .B(net513),
    .C(_1190_),
    .X(_1191_));
 sky130_fd_sc_hd__a21o_1 _2782_ (.A1(_1112_),
    .A2(_1189_),
    .B1(_1191_),
    .X(_0072_));
 sky130_fd_sc_hd__and3_1 _2783_ (.A(net105),
    .B(net575),
    .C(_1190_),
    .X(_1192_));
 sky130_fd_sc_hd__a21o_1 _2784_ (.A1(_1114_),
    .A2(_1189_),
    .B1(_1192_),
    .X(_0073_));
 sky130_fd_sc_hd__and3_1 _2785_ (.A(net105),
    .B(net521),
    .C(_1190_),
    .X(_1193_));
 sky130_fd_sc_hd__a21o_1 _2786_ (.A1(_1116_),
    .A2(_1189_),
    .B1(_1193_),
    .X(_0074_));
 sky130_fd_sc_hd__and3_1 _2787_ (.A(net105),
    .B(net510),
    .C(_1190_),
    .X(_1194_));
 sky130_fd_sc_hd__a21o_1 _2788_ (.A1(_1118_),
    .A2(_1189_),
    .B1(_1194_),
    .X(_0075_));
 sky130_fd_sc_hd__and3_1 _2789_ (.A(net105),
    .B(net555),
    .C(_1190_),
    .X(_1195_));
 sky130_fd_sc_hd__a21o_1 _2790_ (.A1(_1120_),
    .A2(_1189_),
    .B1(_1195_),
    .X(_0076_));
 sky130_fd_sc_hd__and3_1 _2791_ (.A(net108),
    .B(net515),
    .C(_1190_),
    .X(_1196_));
 sky130_fd_sc_hd__a21o_1 _2792_ (.A1(_1123_),
    .A2(_1189_),
    .B1(_1196_),
    .X(_0077_));
 sky130_fd_sc_hd__and3_1 _2793_ (.A(net105),
    .B(net608),
    .C(_1190_),
    .X(_1197_));
 sky130_fd_sc_hd__a21o_1 _2794_ (.A1(_1125_),
    .A2(_1189_),
    .B1(_1197_),
    .X(_0078_));
 sky130_fd_sc_hd__and3_1 _2795_ (.A(net108),
    .B(net545),
    .C(_1190_),
    .X(_1198_));
 sky130_fd_sc_hd__a21o_1 _2796_ (.A1(_1128_),
    .A2(_1189_),
    .B1(_1198_),
    .X(_0079_));
 sky130_fd_sc_hd__and2_2 _2797_ (.A(_0444_),
    .B(_1178_),
    .X(_1199_));
 sky130_fd_sc_hd__nand2_2 _2798_ (.A(_0444_),
    .B(_1178_),
    .Y(_1200_));
 sky130_fd_sc_hd__and3_1 _2799_ (.A(net108),
    .B(net653),
    .C(_1200_),
    .X(_1201_));
 sky130_fd_sc_hd__a21o_1 _2800_ (.A1(_1112_),
    .A2(_1199_),
    .B1(_1201_),
    .X(_0080_));
 sky130_fd_sc_hd__and3_1 _2801_ (.A(net105),
    .B(net559),
    .C(_1200_),
    .X(_1202_));
 sky130_fd_sc_hd__a21o_1 _2802_ (.A1(_1114_),
    .A2(_1199_),
    .B1(_1202_),
    .X(_0081_));
 sky130_fd_sc_hd__and3_1 _2803_ (.A(net105),
    .B(net567),
    .C(_1200_),
    .X(_1203_));
 sky130_fd_sc_hd__a21o_1 _2804_ (.A1(_1116_),
    .A2(_1199_),
    .B1(_1203_),
    .X(_0082_));
 sky130_fd_sc_hd__and3_1 _2805_ (.A(net105),
    .B(net589),
    .C(_1200_),
    .X(_1204_));
 sky130_fd_sc_hd__a21o_1 _2806_ (.A1(_1118_),
    .A2(_1199_),
    .B1(_1204_),
    .X(_0083_));
 sky130_fd_sc_hd__and3_1 _2807_ (.A(net106),
    .B(net606),
    .C(_1200_),
    .X(_1205_));
 sky130_fd_sc_hd__a21o_1 _2808_ (.A1(_1120_),
    .A2(_1199_),
    .B1(_1205_),
    .X(_0084_));
 sky130_fd_sc_hd__and3_1 _2809_ (.A(net107),
    .B(net616),
    .C(_1200_),
    .X(_1206_));
 sky130_fd_sc_hd__a21o_1 _2810_ (.A1(_1123_),
    .A2(_1199_),
    .B1(_1206_),
    .X(_0085_));
 sky130_fd_sc_hd__and3_1 _2811_ (.A(net107),
    .B(net538),
    .C(_1200_),
    .X(_1207_));
 sky130_fd_sc_hd__a21o_1 _2812_ (.A1(_1125_),
    .A2(_1199_),
    .B1(_1207_),
    .X(_0086_));
 sky130_fd_sc_hd__and3_1 _2813_ (.A(net108),
    .B(net648),
    .C(_1200_),
    .X(_1208_));
 sky130_fd_sc_hd__a21o_1 _2814_ (.A1(_1128_),
    .A2(_1199_),
    .B1(_1208_),
    .X(_0087_));
 sky130_fd_sc_hd__and2_2 _2815_ (.A(_1146_),
    .B(_1178_),
    .X(_1209_));
 sky130_fd_sc_hd__nand2_2 _2816_ (.A(_1146_),
    .B(_1178_),
    .Y(_1210_));
 sky130_fd_sc_hd__and3_1 _2817_ (.A(net107),
    .B(net553),
    .C(_1210_),
    .X(_1211_));
 sky130_fd_sc_hd__a21o_1 _2818_ (.A1(_1112_),
    .A2(_1209_),
    .B1(_1211_),
    .X(_0088_));
 sky130_fd_sc_hd__and3_1 _2819_ (.A(net106),
    .B(net511),
    .C(_1210_),
    .X(_1212_));
 sky130_fd_sc_hd__a21o_1 _2820_ (.A1(_1114_),
    .A2(_1209_),
    .B1(_1212_),
    .X(_0089_));
 sky130_fd_sc_hd__and3_1 _2821_ (.A(net106),
    .B(net581),
    .C(_1210_),
    .X(_1213_));
 sky130_fd_sc_hd__a21o_1 _2822_ (.A1(_1116_),
    .A2(_1209_),
    .B1(_1213_),
    .X(_0090_));
 sky130_fd_sc_hd__and3_1 _2823_ (.A(net106),
    .B(net535),
    .C(_1210_),
    .X(_1214_));
 sky130_fd_sc_hd__a21o_1 _2824_ (.A1(_1118_),
    .A2(_1209_),
    .B1(_1214_),
    .X(_0091_));
 sky130_fd_sc_hd__and3_1 _2825_ (.A(net106),
    .B(net531),
    .C(_1210_),
    .X(_1215_));
 sky130_fd_sc_hd__a21o_1 _2826_ (.A1(_1120_),
    .A2(_1209_),
    .B1(_1215_),
    .X(_0092_));
 sky130_fd_sc_hd__and3_1 _2827_ (.A(net107),
    .B(net618),
    .C(_1210_),
    .X(_1216_));
 sky130_fd_sc_hd__a21o_1 _2828_ (.A1(_1123_),
    .A2(_1209_),
    .B1(_1216_),
    .X(_0093_));
 sky130_fd_sc_hd__and3_1 _2829_ (.A(net107),
    .B(net491),
    .C(_1210_),
    .X(_1217_));
 sky130_fd_sc_hd__a21o_1 _2830_ (.A1(_1125_),
    .A2(_1209_),
    .B1(_1217_),
    .X(_0094_));
 sky130_fd_sc_hd__and3_1 _2831_ (.A(net107),
    .B(net611),
    .C(_1210_),
    .X(_1218_));
 sky130_fd_sc_hd__a21o_1 _2832_ (.A1(_1128_),
    .A2(_1209_),
    .B1(_1218_),
    .X(_0095_));
 sky130_fd_sc_hd__nor2_2 _2833_ (.A(_1806_),
    .B(_1815_),
    .Y(_1219_));
 sky130_fd_sc_hd__or2_1 _2834_ (.A(_1806_),
    .B(_1815_),
    .X(_1220_));
 sky130_fd_sc_hd__nor2_2 _2835_ (.A(_1108_),
    .B(_1220_),
    .Y(_1221_));
 sky130_fd_sc_hd__or2_2 _2836_ (.A(_1108_),
    .B(_1220_),
    .X(_1222_));
 sky130_fd_sc_hd__and3_1 _2837_ (.A(net109),
    .B(net706),
    .C(_1222_),
    .X(_1223_));
 sky130_fd_sc_hd__a21o_1 _2838_ (.A1(_1112_),
    .A2(_1221_),
    .B1(_1223_),
    .X(_0096_));
 sky130_fd_sc_hd__and3_1 _2839_ (.A(net109),
    .B(net609),
    .C(_1222_),
    .X(_1224_));
 sky130_fd_sc_hd__a21o_1 _2840_ (.A1(_1114_),
    .A2(_1221_),
    .B1(_1224_),
    .X(_0097_));
 sky130_fd_sc_hd__and3_1 _2841_ (.A(net109),
    .B(net583),
    .C(_1222_),
    .X(_1225_));
 sky130_fd_sc_hd__a21o_1 _2842_ (.A1(_1116_),
    .A2(_1221_),
    .B1(_1225_),
    .X(_0098_));
 sky130_fd_sc_hd__and3_1 _2843_ (.A(net109),
    .B(net588),
    .C(_1222_),
    .X(_1226_));
 sky130_fd_sc_hd__a21o_1 _2844_ (.A1(_1118_),
    .A2(_1221_),
    .B1(_1226_),
    .X(_0099_));
 sky130_fd_sc_hd__and3_1 _2845_ (.A(net109),
    .B(net625),
    .C(_1222_),
    .X(_1227_));
 sky130_fd_sc_hd__a21o_1 _2846_ (.A1(_1120_),
    .A2(_1221_),
    .B1(_1227_),
    .X(_0100_));
 sky130_fd_sc_hd__and3_1 _2847_ (.A(net109),
    .B(net624),
    .C(_1222_),
    .X(_1228_));
 sky130_fd_sc_hd__a21o_1 _2848_ (.A1(_1123_),
    .A2(_1221_),
    .B1(_1228_),
    .X(_0101_));
 sky130_fd_sc_hd__and3_1 _2849_ (.A(net110),
    .B(net585),
    .C(_1222_),
    .X(_1229_));
 sky130_fd_sc_hd__a21o_1 _2850_ (.A1(_1125_),
    .A2(_1221_),
    .B1(_1229_),
    .X(_0102_));
 sky130_fd_sc_hd__and3_1 _2851_ (.A(net110),
    .B(net558),
    .C(_1222_),
    .X(_1230_));
 sky130_fd_sc_hd__a21o_1 _2852_ (.A1(_1128_),
    .A2(_1221_),
    .B1(_1230_),
    .X(_0103_));
 sky130_fd_sc_hd__and2_2 _2853_ (.A(_1178_),
    .B(_1219_),
    .X(_1231_));
 sky130_fd_sc_hd__nand2_2 _2854_ (.A(_1178_),
    .B(_1219_),
    .Y(_1232_));
 sky130_fd_sc_hd__and3_1 _2855_ (.A(net107),
    .B(net655),
    .C(_1232_),
    .X(_1233_));
 sky130_fd_sc_hd__a21o_1 _2856_ (.A1(_1112_),
    .A2(_1231_),
    .B1(_1233_),
    .X(_0104_));
 sky130_fd_sc_hd__and3_1 _2857_ (.A(net106),
    .B(net650),
    .C(_1232_),
    .X(_1234_));
 sky130_fd_sc_hd__a21o_1 _2858_ (.A1(_1114_),
    .A2(_1231_),
    .B1(_1234_),
    .X(_0105_));
 sky130_fd_sc_hd__and3_1 _2859_ (.A(net106),
    .B(net518),
    .C(_1232_),
    .X(_1235_));
 sky130_fd_sc_hd__a21o_1 _2860_ (.A1(_1116_),
    .A2(_1231_),
    .B1(_1235_),
    .X(_0106_));
 sky130_fd_sc_hd__and3_1 _2861_ (.A(net106),
    .B(net550),
    .C(_1232_),
    .X(_1236_));
 sky130_fd_sc_hd__a21o_1 _2862_ (.A1(_1118_),
    .A2(_1231_),
    .B1(_1236_),
    .X(_0107_));
 sky130_fd_sc_hd__and3_1 _2863_ (.A(net106),
    .B(net604),
    .C(_1232_),
    .X(_1237_));
 sky130_fd_sc_hd__a21o_1 _2864_ (.A1(_1120_),
    .A2(_1231_),
    .B1(_1237_),
    .X(_0108_));
 sky130_fd_sc_hd__and3_1 _2865_ (.A(net107),
    .B(net638),
    .C(_1232_),
    .X(_1238_));
 sky130_fd_sc_hd__a21o_1 _2866_ (.A1(_1123_),
    .A2(_1231_),
    .B1(_1238_),
    .X(_0109_));
 sky130_fd_sc_hd__and3_1 _2867_ (.A(net107),
    .B(net597),
    .C(_1232_),
    .X(_1239_));
 sky130_fd_sc_hd__a21o_1 _2868_ (.A1(_1125_),
    .A2(_1231_),
    .B1(_1239_),
    .X(_0110_));
 sky130_fd_sc_hd__and3_1 _2869_ (.A(net107),
    .B(net593),
    .C(_1232_),
    .X(_1240_));
 sky130_fd_sc_hd__a21o_1 _2870_ (.A1(_1128_),
    .A2(_1231_),
    .B1(_1240_),
    .X(_0111_));
 sky130_fd_sc_hd__and2_2 _2871_ (.A(_1148_),
    .B(_1219_),
    .X(_1241_));
 sky130_fd_sc_hd__nand2_2 _2872_ (.A(_1148_),
    .B(_1219_),
    .Y(_1242_));
 sky130_fd_sc_hd__and3_1 _2873_ (.A(net104),
    .B(net551),
    .C(_1242_),
    .X(_1243_));
 sky130_fd_sc_hd__a21o_1 _2874_ (.A1(_1112_),
    .A2(_1241_),
    .B1(_1243_),
    .X(_0112_));
 sky130_fd_sc_hd__and3_1 _2875_ (.A(net104),
    .B(net533),
    .C(_1242_),
    .X(_1244_));
 sky130_fd_sc_hd__a21o_1 _2876_ (.A1(_1114_),
    .A2(_1241_),
    .B1(_1244_),
    .X(_0113_));
 sky130_fd_sc_hd__and3_1 _2877_ (.A(net104),
    .B(net715),
    .C(_1242_),
    .X(_1245_));
 sky130_fd_sc_hd__a21o_1 _2878_ (.A1(_1116_),
    .A2(_1241_),
    .B1(_1245_),
    .X(_0114_));
 sky130_fd_sc_hd__and3_1 _2879_ (.A(net104),
    .B(net584),
    .C(_1242_),
    .X(_1246_));
 sky130_fd_sc_hd__a21o_1 _2880_ (.A1(_1118_),
    .A2(_1241_),
    .B1(_1246_),
    .X(_0115_));
 sky130_fd_sc_hd__and3_1 _2881_ (.A(net104),
    .B(net579),
    .C(_1242_),
    .X(_1247_));
 sky130_fd_sc_hd__a21o_1 _2882_ (.A1(_1120_),
    .A2(_1241_),
    .B1(_1247_),
    .X(_0116_));
 sky130_fd_sc_hd__and3_1 _2883_ (.A(net104),
    .B(net527),
    .C(_1242_),
    .X(_1248_));
 sky130_fd_sc_hd__a21o_1 _2884_ (.A1(_1123_),
    .A2(_1241_),
    .B1(_1248_),
    .X(_0117_));
 sky130_fd_sc_hd__and3_1 _2885_ (.A(net104),
    .B(net509),
    .C(_1242_),
    .X(_1249_));
 sky130_fd_sc_hd__a21o_1 _2886_ (.A1(_1125_),
    .A2(_1241_),
    .B1(_1249_),
    .X(_0118_));
 sky130_fd_sc_hd__and3_1 _2887_ (.A(net104),
    .B(net524),
    .C(_1242_),
    .X(_1250_));
 sky130_fd_sc_hd__a21o_1 _2888_ (.A1(_1128_),
    .A2(_1241_),
    .B1(_1250_),
    .X(_0119_));
 sky130_fd_sc_hd__or2_1 _2889_ (.A(net693),
    .B(net431),
    .X(_1251_));
 sky130_fd_sc_hd__nor4_1 _2890_ (.A(net688),
    .B(net817),
    .C(\ROM_spi_cycle[0] ),
    .D(_1251_),
    .Y(_1252_));
 sky130_fd_sc_hd__or4_4 _2891_ (.A(net688),
    .B(net817),
    .C(\ROM_spi_cycle[0] ),
    .D(_1251_),
    .X(_1253_));
 sky130_fd_sc_hd__nor2_1 _2892_ (.A(net477),
    .B(net768),
    .Y(_1254_));
 sky130_fd_sc_hd__or2_2 _2893_ (.A(net477),
    .B(net768),
    .X(_1255_));
 sky130_fd_sc_hd__nor3_2 _2894_ (.A(net720),
    .B(net722),
    .C(net698),
    .Y(_1256_));
 sky130_fd_sc_hd__or3_1 _2895_ (.A(net720),
    .B(net722),
    .C(net698),
    .X(_1257_));
 sky130_fd_sc_hd__nor2_1 _2896_ (.A(net661),
    .B(\startup_cycle[2] ),
    .Y(_1258_));
 sky130_fd_sc_hd__or2_1 _2897_ (.A(net661),
    .B(\startup_cycle[2] ),
    .X(_1259_));
 sky130_fd_sc_hd__and3_4 _2898_ (.A(_1254_),
    .B(_1256_),
    .C(_1258_),
    .X(_1260_));
 sky130_fd_sc_hd__or3_1 _2899_ (.A(_1255_),
    .B(_1257_),
    .C(_1259_),
    .X(_1261_));
 sky130_fd_sc_hd__nand2_2 _2900_ (.A(net64),
    .B(_1260_),
    .Y(_1262_));
 sky130_fd_sc_hd__or2_2 _2901_ (.A(\mem_cycle[3] ),
    .B(\mem_cycle[2] ),
    .X(_1263_));
 sky130_fd_sc_hd__or4_2 _2902_ (.A(\mem_cycle[5] ),
    .B(\mem_cycle[4] ),
    .C(\mem_cycle[1] ),
    .D(\mem_cycle[0] ),
    .X(_1264_));
 sky130_fd_sc_hd__nor2_1 _2903_ (.A(_1263_),
    .B(_1264_),
    .Y(_1265_));
 sky130_fd_sc_hd__or2_1 _2904_ (.A(_1263_),
    .B(_1264_),
    .X(_1266_));
 sky130_fd_sc_hd__a22o_1 _2905_ (.A1(\S8x305.A[12] ),
    .A2(_1754_),
    .B1(_1760_),
    .B2(\S8x305.A[3] ),
    .X(_1267_));
 sky130_fd_sc_hd__a22o_1 _2906_ (.A1(_1746_),
    .A2(\last_A[4] ),
    .B1(_1761_),
    .B2(\S8x305.A[2] ),
    .X(_1268_));
 sky130_fd_sc_hd__a22o_1 _2907_ (.A1(\S8x305.A[9] ),
    .A2(_1757_),
    .B1(_1759_),
    .B2(\S8x305.A[4] ),
    .X(_1269_));
 sky130_fd_sc_hd__a221o_1 _2908_ (.A1(\S8x305.A[0] ),
    .A2(_1752_),
    .B1(\last_A[9] ),
    .B2(_1742_),
    .C1(_1267_),
    .X(_1270_));
 sky130_fd_sc_hd__o22a_1 _2909_ (.A1(_1743_),
    .A2(\last_A[7] ),
    .B1(_1762_),
    .B2(net786),
    .X(_1271_));
 sky130_fd_sc_hd__o221a_1 _2910_ (.A1(net815),
    .A2(_1755_),
    .B1(_1756_),
    .B2(net453),
    .C1(_1271_),
    .X(_1272_));
 sky130_fd_sc_hd__o22a_1 _2911_ (.A1(net370),
    .A2(_1751_),
    .B1(_1754_),
    .B2(net773),
    .X(_1273_));
 sky130_fd_sc_hd__o221a_1 _2912_ (.A1(_1741_),
    .A2(net836),
    .B1(\last_A[6] ),
    .B2(_1744_),
    .C1(_1273_),
    .X(_1274_));
 sky130_fd_sc_hd__a221o_1 _2913_ (.A1(_1750_),
    .A2(\ROM_addr_buff[1] ),
    .B1(\last_A[2] ),
    .B2(_1748_),
    .C1(_1268_),
    .X(_1275_));
 sky130_fd_sc_hd__a221o_1 _2914_ (.A1(\S8x305.A[11] ),
    .A2(_1755_),
    .B1(\last_A[6] ),
    .B2(_1744_),
    .C1(_1275_),
    .X(_1276_));
 sky130_fd_sc_hd__a22o_1 _2915_ (.A1(_1743_),
    .A2(\last_A[7] ),
    .B1(\last_A[5] ),
    .B2(_1745_),
    .X(_1277_));
 sky130_fd_sc_hd__a221o_1 _2916_ (.A1(\S8x305.A[5] ),
    .A2(_1758_),
    .B1(_1762_),
    .B2(\S8x305.A[1] ),
    .C1(_1277_),
    .X(_1278_));
 sky130_fd_sc_hd__a221o_1 _2917_ (.A1(net370),
    .A2(_1751_),
    .B1(\last_A[3] ),
    .B2(_1747_),
    .C1(_1269_),
    .X(_1279_));
 sky130_fd_sc_hd__or4_1 _2918_ (.A(_1266_),
    .B(_1270_),
    .C(_1278_),
    .D(_1279_),
    .X(_1280_));
 sky130_fd_sc_hd__nor2_1 _2919_ (.A(_1276_),
    .B(_1280_),
    .Y(_1281_));
 sky130_fd_sc_hd__a31o_2 _2920_ (.A1(_1272_),
    .A2(net837),
    .A3(_1281_),
    .B1(_1262_),
    .X(_1282_));
 sky130_fd_sc_hd__nand2_1 _2921_ (.A(net796),
    .B(net835),
    .Y(_1283_));
 sky130_fd_sc_hd__nor2_1 _2922_ (.A(_1282_),
    .B(_1283_),
    .Y(_1284_));
 sky130_fd_sc_hd__nand2_1 _2923_ (.A(net830),
    .B(net443),
    .Y(_1285_));
 sky130_fd_sc_hd__or4_4 _2924_ (.A(_1764_),
    .B(_1282_),
    .C(_1283_),
    .D(_1285_),
    .X(_1286_));
 sky130_fd_sc_hd__nor2_2 _2925_ (.A(net826),
    .B(_1286_),
    .Y(_1287_));
 sky130_fd_sc_hd__or3_1 _2926_ (.A(net4),
    .B(\mem_cycle[5] ),
    .C(_1286_),
    .X(_1288_));
 sky130_fd_sc_hd__o211a_1 _2927_ (.A1(net425),
    .A2(_1287_),
    .B1(_1288_),
    .C1(net97),
    .X(_0120_));
 sky130_fd_sc_hd__or3_1 _2928_ (.A(net5),
    .B(\mem_cycle[5] ),
    .C(_1286_),
    .X(_1289_));
 sky130_fd_sc_hd__o211a_1 _2929_ (.A1(net421),
    .A2(_1287_),
    .B1(_1289_),
    .C1(net97),
    .X(_0121_));
 sky130_fd_sc_hd__or3_1 _2930_ (.A(net6),
    .B(\mem_cycle[5] ),
    .C(_1286_),
    .X(_1290_));
 sky130_fd_sc_hd__o211a_1 _2931_ (.A1(net405),
    .A2(_1287_),
    .B1(_1290_),
    .C1(net97),
    .X(_0122_));
 sky130_fd_sc_hd__or3_1 _2932_ (.A(net7),
    .B(\mem_cycle[5] ),
    .C(_1286_),
    .X(_1291_));
 sky130_fd_sc_hd__o211a_1 _2933_ (.A1(net427),
    .A2(_1287_),
    .B1(_1291_),
    .C1(net97),
    .X(_0123_));
 sky130_fd_sc_hd__or3b_1 _2934_ (.A(\mem_cycle[0] ),
    .B(_1263_),
    .C_N(net796),
    .X(_1292_));
 sky130_fd_sc_hd__nor3_1 _2935_ (.A(_1763_),
    .B(net822),
    .C(_1292_),
    .Y(_1293_));
 sky130_fd_sc_hd__and2b_1 _2936_ (.A_N(_1282_),
    .B(net827),
    .X(_1294_));
 sky130_fd_sc_hd__or2_1 _2937_ (.A(_1266_),
    .B(_1282_),
    .X(_1295_));
 sky130_fd_sc_hd__o211a_1 _2938_ (.A1(net599),
    .A2(_1294_),
    .B1(net58),
    .C1(net97),
    .X(_0124_));
 sky130_fd_sc_hd__nor2_1 _2939_ (.A(_1782_),
    .B(net32),
    .Y(_1296_));
 sky130_fd_sc_hd__and3_4 _2940_ (.A(net34),
    .B(_0887_),
    .C(_1296_),
    .X(_1297_));
 sky130_fd_sc_hd__o21ai_1 _2941_ (.A1(net633),
    .A2(_1297_),
    .B1(net102),
    .Y(_1298_));
 sky130_fd_sc_hd__a21oi_1 _2942_ (.A1(net74),
    .A2(_1297_),
    .B1(_1298_),
    .Y(_0125_));
 sky130_fd_sc_hd__o21ai_1 _2943_ (.A1(net620),
    .A2(_1297_),
    .B1(net102),
    .Y(_1299_));
 sky130_fd_sc_hd__a21oi_1 _2944_ (.A1(net75),
    .A2(_1297_),
    .B1(_1299_),
    .Y(_0126_));
 sky130_fd_sc_hd__o21ai_1 _2945_ (.A1(net704),
    .A2(_1297_),
    .B1(net102),
    .Y(_1300_));
 sky130_fd_sc_hd__a21oi_1 _2946_ (.A1(net76),
    .A2(_1297_),
    .B1(_1300_),
    .Y(_0127_));
 sky130_fd_sc_hd__o21ai_1 _2947_ (.A1(net657),
    .A2(_1297_),
    .B1(net102),
    .Y(_1301_));
 sky130_fd_sc_hd__a21oi_1 _2948_ (.A1(net77),
    .A2(_1297_),
    .B1(_1301_),
    .Y(_0128_));
 sky130_fd_sc_hd__o21ai_1 _2949_ (.A1(net668),
    .A2(_1297_),
    .B1(net102),
    .Y(_1302_));
 sky130_fd_sc_hd__a21oi_1 _2950_ (.A1(net78),
    .A2(_1297_),
    .B1(_1302_),
    .Y(_0129_));
 sky130_fd_sc_hd__o21ai_1 _2951_ (.A1(net665),
    .A2(_1297_),
    .B1(net102),
    .Y(_1303_));
 sky130_fd_sc_hd__a21oi_1 _2952_ (.A1(net79),
    .A2(_1297_),
    .B1(_1303_),
    .Y(_0130_));
 sky130_fd_sc_hd__o21ai_1 _2953_ (.A1(net719),
    .A2(_1297_),
    .B1(net102),
    .Y(_1304_));
 sky130_fd_sc_hd__a21oi_1 _2954_ (.A1(net80),
    .A2(_1297_),
    .B1(_1304_),
    .Y(_0131_));
 sky130_fd_sc_hd__o21ai_1 _2955_ (.A1(net764),
    .A2(_1297_),
    .B1(net94),
    .Y(_1305_));
 sky130_fd_sc_hd__a21oi_1 _2956_ (.A1(net81),
    .A2(_1297_),
    .B1(_1305_),
    .Y(_0132_));
 sky130_fd_sc_hd__nor2_1 _2957_ (.A(net726),
    .B(net64),
    .Y(_1306_));
 sky130_fd_sc_hd__nand2_1 _2958_ (.A(net661),
    .B(\startup_cycle[2] ),
    .Y(_1307_));
 sky130_fd_sc_hd__and2_1 _2959_ (.A(net477),
    .B(net768),
    .X(_1308_));
 sky130_fd_sc_hd__and3_2 _2960_ (.A(net661),
    .B(\startup_cycle[2] ),
    .C(_1308_),
    .X(_1309_));
 sky130_fd_sc_hd__a31o_1 _2961_ (.A1(_1768_),
    .A2(\startup_cycle[2] ),
    .A3(_1254_),
    .B1(_1309_),
    .X(_1310_));
 sky130_fd_sc_hd__nand2_1 _2962_ (.A(net477),
    .B(_1769_),
    .Y(_1311_));
 sky130_fd_sc_hd__nor2_1 _2963_ (.A(_1768_),
    .B(\startup_cycle[2] ),
    .Y(_1312_));
 sky130_fd_sc_hd__a31o_1 _2964_ (.A1(\startup_cycle[1] ),
    .A2(_1769_),
    .A3(_1312_),
    .B1(_1310_),
    .X(_1313_));
 sky130_fd_sc_hd__a2bb2o_1 _2965_ (.A1_N(_1255_),
    .A2_N(_1307_),
    .B1(_1308_),
    .B2(_1312_),
    .X(_1314_));
 sky130_fd_sc_hd__o21a_1 _2966_ (.A1(_1313_),
    .A2(_1314_),
    .B1(_1256_),
    .X(_1315_));
 sky130_fd_sc_hd__and4_1 _2967_ (.A(_1768_),
    .B(\startup_cycle[2] ),
    .C(_1256_),
    .D(_1308_),
    .X(_1316_));
 sky130_fd_sc_hd__nor2_1 _2968_ (.A(_1315_),
    .B(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__nor2_1 _2969_ (.A(\startup_cycle[1] ),
    .B(_1769_),
    .Y(_1318_));
 sky130_fd_sc_hd__a311o_1 _2970_ (.A1(_1256_),
    .A2(_1258_),
    .A3(_1318_),
    .B1(_1316_),
    .C1(_1315_),
    .X(_1319_));
 sky130_fd_sc_hd__o21ba_1 _2971_ (.A1(_1253_),
    .A2(_1319_),
    .B1_N(_1306_),
    .X(_1320_));
 sky130_fd_sc_hd__nand2_1 _2972_ (.A(net726),
    .B(\ROM_spi_cycle[0] ),
    .Y(_1321_));
 sky130_fd_sc_hd__o211a_1 _2973_ (.A1(\ROM_spi_cycle[0] ),
    .A2(_1320_),
    .B1(net727),
    .C1(net93),
    .X(_0133_));
 sky130_fd_sc_hd__or2_1 _2974_ (.A(_1770_),
    .B(_1251_),
    .X(_1322_));
 sky130_fd_sc_hd__a31o_1 _2975_ (.A1(net726),
    .A2(\ROM_spi_cycle[0] ),
    .A3(_1322_),
    .B1(net817),
    .X(_1323_));
 sky130_fd_sc_hd__and3_1 _2976_ (.A(net726),
    .B(net817),
    .C(\ROM_spi_cycle[0] ),
    .X(_1324_));
 sky130_fd_sc_hd__and3b_1 _2977_ (.A_N(_1324_),
    .B(net93),
    .C(net818),
    .X(_0134_));
 sky130_fd_sc_hd__and2_1 _2978_ (.A(net431),
    .B(_1324_),
    .X(_1325_));
 sky130_fd_sc_hd__nor2_1 _2979_ (.A(net91),
    .B(_1325_),
    .Y(_1326_));
 sky130_fd_sc_hd__o21a_1 _2980_ (.A1(net431),
    .A2(_1324_),
    .B1(_1326_),
    .X(_0135_));
 sky130_fd_sc_hd__or2_1 _2981_ (.A(net693),
    .B(_1325_),
    .X(_1327_));
 sky130_fd_sc_hd__nand2_1 _2982_ (.A(net693),
    .B(_1325_),
    .Y(_1328_));
 sky130_fd_sc_hd__and3_1 _2983_ (.A(net93),
    .B(_1327_),
    .C(net694),
    .X(_0136_));
 sky130_fd_sc_hd__nand2_1 _2984_ (.A(\ROM_spi_cycle[3] ),
    .B(net431),
    .Y(_1329_));
 sky130_fd_sc_hd__mux2_1 _2985_ (.A0(_1251_),
    .A1(_1329_),
    .S(\ROM_spi_cycle[1] ),
    .X(_1330_));
 sky130_fd_sc_hd__nand2_1 _2986_ (.A(_1770_),
    .B(_1328_),
    .Y(_1331_));
 sky130_fd_sc_hd__o311a_1 _2987_ (.A1(_1770_),
    .A2(_1321_),
    .A3(_1330_),
    .B1(_1331_),
    .C1(net93),
    .X(_0137_));
 sky130_fd_sc_hd__nor2_2 _2988_ (.A(_1253_),
    .B(_1260_),
    .Y(_1332_));
 sky130_fd_sc_hd__nor2_1 _2989_ (.A(_1259_),
    .B(_1311_),
    .Y(_1333_));
 sky130_fd_sc_hd__and4b_1 _2990_ (.A_N(net722),
    .B(net698),
    .C(_1333_),
    .D(net720),
    .X(_1334_));
 sky130_fd_sc_hd__o21a_1 _2991_ (.A1(net768),
    .A2(_1334_),
    .B1(_1332_),
    .X(_1335_));
 sky130_fd_sc_hd__nor2_1 _2992_ (.A(net768),
    .B(_1332_),
    .Y(_1336_));
 sky130_fd_sc_hd__o21ai_1 _2993_ (.A1(_1335_),
    .A2(net769),
    .B1(net94),
    .Y(_0138_));
 sky130_fd_sc_hd__o21ai_1 _2994_ (.A1(net477),
    .A2(_1335_),
    .B1(net94),
    .Y(_1337_));
 sky130_fd_sc_hd__a21oi_1 _2995_ (.A1(net477),
    .A2(_1335_),
    .B1(_1337_),
    .Y(_0139_));
 sky130_fd_sc_hd__a21o_1 _2996_ (.A1(net64),
    .A2(_1308_),
    .B1(net806),
    .X(_1338_));
 sky130_fd_sc_hd__nand3_1 _2997_ (.A(net806),
    .B(net64),
    .C(_1308_),
    .Y(_1339_));
 sky130_fd_sc_hd__and3_1 _2998_ (.A(net93),
    .B(_1338_),
    .C(net807),
    .X(_0140_));
 sky130_fd_sc_hd__a221oi_1 _2999_ (.A1(net64),
    .A2(_1309_),
    .B1(_1339_),
    .B2(_1768_),
    .C1(net91),
    .Y(_0141_));
 sky130_fd_sc_hd__a21oi_1 _3000_ (.A1(_1309_),
    .A2(_1332_),
    .B1(net698),
    .Y(_1340_));
 sky130_fd_sc_hd__and3_1 _3001_ (.A(net698),
    .B(_1309_),
    .C(_1332_),
    .X(_1341_));
 sky130_fd_sc_hd__a2111oi_1 _3002_ (.A1(_1332_),
    .A2(_1334_),
    .B1(net699),
    .C1(_1341_),
    .D1(net91),
    .Y(_0142_));
 sky130_fd_sc_hd__and3_1 _3003_ (.A(net722),
    .B(net698),
    .C(_1309_),
    .X(_1342_));
 sky130_fd_sc_hd__nand2_1 _3004_ (.A(_1332_),
    .B(_1342_),
    .Y(_1343_));
 sky130_fd_sc_hd__o211a_1 _3005_ (.A1(net722),
    .A2(_1341_),
    .B1(_1343_),
    .C1(net94),
    .X(_0143_));
 sky130_fd_sc_hd__o311a_1 _3006_ (.A1(_1260_),
    .A2(_1334_),
    .A3(_1342_),
    .B1(net64),
    .C1(net720),
    .X(_1344_));
 sky130_fd_sc_hd__a211oi_1 _3007_ (.A1(_1767_),
    .A2(_1343_),
    .B1(_1344_),
    .C1(net91),
    .Y(_0144_));
 sky130_fd_sc_hd__or2_1 _3008_ (.A(_1282_),
    .B(_1293_),
    .X(_1345_));
 sky130_fd_sc_hd__nand2_1 _3009_ (.A(net835),
    .B(net838),
    .Y(_1346_));
 sky130_fd_sc_hd__o21ai_1 _3010_ (.A1(net835),
    .A2(_1345_),
    .B1(_1346_),
    .Y(_1347_));
 sky130_fd_sc_hd__and3_1 _3011_ (.A(\last_addr[3] ),
    .B(\last_addr[2] ),
    .C(\last_addr[1] ),
    .X(_1348_));
 sky130_fd_sc_hd__and2_1 _3012_ (.A(\last_addr[4] ),
    .B(_1348_),
    .X(_1349_));
 sky130_fd_sc_hd__and3_1 _3013_ (.A(\last_addr[5] ),
    .B(\last_addr[4] ),
    .C(_1348_),
    .X(_1350_));
 sky130_fd_sc_hd__and3_1 _3014_ (.A(\last_addr[7] ),
    .B(\last_addr[6] ),
    .C(_1350_),
    .X(_1351_));
 sky130_fd_sc_hd__and3_1 _3015_ (.A(\last_addr[9] ),
    .B(\last_addr[8] ),
    .C(_1351_),
    .X(_1352_));
 sky130_fd_sc_hd__and2_1 _3016_ (.A(\last_addr[10] ),
    .B(_1352_),
    .X(_1353_));
 sky130_fd_sc_hd__and3_1 _3017_ (.A(net716),
    .B(net774),
    .C(_1353_),
    .X(_1354_));
 sky130_fd_sc_hd__a21oi_1 _3018_ (.A1(net774),
    .A2(_1353_),
    .B1(net716),
    .Y(_1355_));
 sky130_fd_sc_hd__nor2_1 _3019_ (.A(_1354_),
    .B(_1355_),
    .Y(_1356_));
 sky130_fd_sc_hd__xnor2_1 _3020_ (.A(net774),
    .B(_1353_),
    .Y(_1357_));
 sky130_fd_sc_hd__a22o_1 _3021_ (.A1(\last_addr[13] ),
    .A2(_1354_),
    .B1(_1357_),
    .B2(net718),
    .X(_1358_));
 sky130_fd_sc_hd__o21ba_1 _3022_ (.A1(net718),
    .A2(_1357_),
    .B1_N(_1358_),
    .X(_1359_));
 sky130_fd_sc_hd__nor2_1 _3023_ (.A(net682),
    .B(_1352_),
    .Y(_1360_));
 sky130_fd_sc_hd__or3_1 _3024_ (.A(net767),
    .B(_1353_),
    .C(_1360_),
    .X(_1361_));
 sky130_fd_sc_hd__o21ai_1 _3025_ (.A1(_1353_),
    .A2(_1360_),
    .B1(net767),
    .Y(_1362_));
 sky130_fd_sc_hd__a21oi_1 _3026_ (.A1(\last_addr[8] ),
    .A2(_1351_),
    .B1(\last_addr[9] ),
    .Y(_1363_));
 sky130_fd_sc_hd__nor2_1 _3027_ (.A(_1352_),
    .B(_1363_),
    .Y(_1364_));
 sky130_fd_sc_hd__xnor2_1 _3028_ (.A(\ROM_addr_buff[9] ),
    .B(_1364_),
    .Y(_1365_));
 sky130_fd_sc_hd__xnor2_1 _3029_ (.A(\last_addr[8] ),
    .B(_1351_),
    .Y(_1366_));
 sky130_fd_sc_hd__xnor2_1 _3030_ (.A(\ROM_addr_buff[8] ),
    .B(_1366_),
    .Y(_1367_));
 sky130_fd_sc_hd__a21oi_1 _3031_ (.A1(\last_addr[6] ),
    .A2(_1350_),
    .B1(\last_addr[7] ),
    .Y(_1368_));
 sky130_fd_sc_hd__or2_1 _3032_ (.A(_1351_),
    .B(_1368_),
    .X(_1369_));
 sky130_fd_sc_hd__xnor2_1 _3033_ (.A(\ROM_addr_buff[7] ),
    .B(_1369_),
    .Y(_1370_));
 sky130_fd_sc_hd__xnor2_1 _3034_ (.A(\ROM_addr_buff[6] ),
    .B(\last_addr[6] ),
    .Y(_1371_));
 sky130_fd_sc_hd__nor2_1 _3035_ (.A(\last_addr[5] ),
    .B(_1349_),
    .Y(_1372_));
 sky130_fd_sc_hd__or3_1 _3036_ (.A(\mem_cycle[4] ),
    .B(net848),
    .C(_1263_),
    .X(_1373_));
 sky130_fd_sc_hd__and3b_4 _3037_ (.A_N(_1373_),
    .B(_1763_),
    .C(net835),
    .X(_1374_));
 sky130_fd_sc_hd__xnor2_1 _3038_ (.A(\ROM_addr_buff[1] ),
    .B(\last_addr[1] ),
    .Y(_1375_));
 sky130_fd_sc_hd__nor2_1 _3039_ (.A(\last_addr[4] ),
    .B(_1348_),
    .Y(_1376_));
 sky130_fd_sc_hd__or2_1 _3040_ (.A(_1349_),
    .B(_1376_),
    .X(_1377_));
 sky130_fd_sc_hd__or2_1 _3041_ (.A(_1350_),
    .B(_1372_),
    .X(_1378_));
 sky130_fd_sc_hd__a21oi_1 _3042_ (.A1(\last_addr[2] ),
    .A2(\last_addr[1] ),
    .B1(\last_addr[3] ),
    .Y(_1379_));
 sky130_fd_sc_hd__or2_1 _3043_ (.A(_1348_),
    .B(_1379_),
    .X(_1380_));
 sky130_fd_sc_hd__xnor2_1 _3044_ (.A(\ROM_addr_buff[3] ),
    .B(_1380_),
    .Y(_1381_));
 sky130_fd_sc_hd__xnor2_1 _3045_ (.A(\last_addr[2] ),
    .B(\last_addr[1] ),
    .Y(_1382_));
 sky130_fd_sc_hd__xnor2_1 _3046_ (.A(\ROM_addr_buff[2] ),
    .B(_1382_),
    .Y(_1383_));
 sky130_fd_sc_hd__xnor2_1 _3047_ (.A(\ROM_addr_buff[4] ),
    .B(_1377_),
    .Y(_1384_));
 sky130_fd_sc_hd__xnor2_1 _3048_ (.A(net841),
    .B(_1356_),
    .Y(_1385_));
 sky130_fd_sc_hd__o21a_1 _3049_ (.A1(\last_addr[13] ),
    .A2(_1354_),
    .B1(net738),
    .X(_1386_));
 sky130_fd_sc_hd__nor3_1 _3050_ (.A(net738),
    .B(\last_addr[13] ),
    .C(_1354_),
    .Y(_1387_));
 sky130_fd_sc_hd__xnor2_1 _3051_ (.A(\ROM_addr_buff[5] ),
    .B(_1378_),
    .Y(_1388_));
 sky130_fd_sc_hd__or4b_1 _3052_ (.A(\last_addr[0] ),
    .B(_1375_),
    .C(_1383_),
    .D_N(_1374_),
    .X(_1389_));
 sky130_fd_sc_hd__or4_1 _3053_ (.A(_1381_),
    .B(_1384_),
    .C(_1388_),
    .D(_1389_),
    .X(_1390_));
 sky130_fd_sc_hd__xnor2_1 _3054_ (.A(_1350_),
    .B(_1371_),
    .Y(_1391_));
 sky130_fd_sc_hd__or4_1 _3055_ (.A(_1367_),
    .B(_1370_),
    .C(_1390_),
    .D(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__and4b_1 _3056_ (.A_N(_1392_),
    .B(_1362_),
    .C(_1361_),
    .D(_1365_),
    .X(_1393_));
 sky130_fd_sc_hd__o2111a_1 _3057_ (.A1(_1386_),
    .A2(_1387_),
    .B1(_1393_),
    .C1(_1385_),
    .D1(_1359_),
    .X(_1394_));
 sky130_fd_sc_hd__and2b_1 _3058_ (.A_N(_1282_),
    .B(net842),
    .X(_1395_));
 sky130_fd_sc_hd__o21a_1 _3059_ (.A1(_1347_),
    .A2(_1395_),
    .B1(net94),
    .X(_0145_));
 sky130_fd_sc_hd__xnor2_1 _3060_ (.A(net796),
    .B(net835),
    .Y(_1396_));
 sky130_fd_sc_hd__o2bb2a_1 _3061_ (.A1_N(net796),
    .A2_N(_1282_),
    .B1(_1345_),
    .B2(_1396_),
    .X(_1397_));
 sky130_fd_sc_hd__nor2_1 _3062_ (.A(net91),
    .B(_1397_),
    .Y(_0146_));
 sky130_fd_sc_hd__o21ai_1 _3063_ (.A1(net443),
    .A2(_1284_),
    .B1(net97),
    .Y(_1398_));
 sky130_fd_sc_hd__a21oi_1 _3064_ (.A1(net443),
    .A2(_1284_),
    .B1(_1398_),
    .Y(_0147_));
 sky130_fd_sc_hd__nand2b_1 _3065_ (.A_N(net830),
    .B(_1282_),
    .Y(_1399_));
 sky130_fd_sc_hd__nor2_1 _3066_ (.A(_1765_),
    .B(_1283_),
    .Y(_1400_));
 sky130_fd_sc_hd__xor2_1 _3067_ (.A(net830),
    .B(_1400_),
    .X(_1401_));
 sky130_fd_sc_hd__o311a_1 _3068_ (.A1(_1282_),
    .A2(_1394_),
    .A3(_1401_),
    .B1(net831),
    .C1(net95),
    .X(_0148_));
 sky130_fd_sc_hd__a31o_1 _3069_ (.A1(\mem_cycle[3] ),
    .A2(net443),
    .A3(_1284_),
    .B1(net822),
    .X(_1402_));
 sky130_fd_sc_hd__a21oi_1 _3070_ (.A1(_1286_),
    .A2(net823),
    .B1(_1395_),
    .Y(_1403_));
 sky130_fd_sc_hd__nor2_1 _3071_ (.A(net91),
    .B(net824),
    .Y(_0149_));
 sky130_fd_sc_hd__and2_1 _3072_ (.A(net826),
    .B(_1286_),
    .X(_1404_));
 sky130_fd_sc_hd__nor2_1 _3073_ (.A(net827),
    .B(_1374_),
    .Y(_1405_));
 sky130_fd_sc_hd__o221a_1 _3074_ (.A1(_1287_),
    .A2(_1404_),
    .B1(_1405_),
    .B2(net838),
    .C1(net97),
    .X(_0150_));
 sky130_fd_sc_hd__nand2_1 _3075_ (.A(\startup_cycle[2] ),
    .B(_1318_),
    .Y(_1406_));
 sky130_fd_sc_hd__nand2_1 _3076_ (.A(_1254_),
    .B(_1312_),
    .Y(_1407_));
 sky130_fd_sc_hd__and3b_1 _3077_ (.A_N(_1333_),
    .B(_1406_),
    .C(_1407_),
    .X(_1408_));
 sky130_fd_sc_hd__or3_1 _3078_ (.A(_1767_),
    .B(net722),
    .C(net698),
    .X(_1409_));
 sky130_fd_sc_hd__o32a_1 _3079_ (.A1(_1307_),
    .A2(_1311_),
    .A3(_1409_),
    .B1(_1408_),
    .B2(_1257_),
    .X(_1410_));
 sky130_fd_sc_hd__nand2_1 _3080_ (.A(_1261_),
    .B(_1410_),
    .Y(_1411_));
 sky130_fd_sc_hd__nor2_1 _3081_ (.A(_1319_),
    .B(_1411_),
    .Y(_1412_));
 sky130_fd_sc_hd__a21o_1 _3082_ (.A1(_1260_),
    .A2(_1265_),
    .B1(_1253_),
    .X(_1413_));
 sky130_fd_sc_hd__or4b_2 _3083_ (.A(\mem_cycle[5] ),
    .B(\mem_cycle[4] ),
    .C(\mem_cycle[0] ),
    .D_N(\mem_cycle[1] ),
    .X(_1414_));
 sky130_fd_sc_hd__inv_2 _3084_ (.A(_1414_),
    .Y(_1415_));
 sky130_fd_sc_hd__or2_1 _3085_ (.A(_1263_),
    .B(_1414_),
    .X(_1416_));
 sky130_fd_sc_hd__or3b_1 _3086_ (.A(_1261_),
    .B(_1265_),
    .C_N(_1416_),
    .X(_1417_));
 sky130_fd_sc_hd__nor2_1 _3087_ (.A(_1374_),
    .B(_1417_),
    .Y(_1418_));
 sky130_fd_sc_hd__or2_1 _3088_ (.A(_1261_),
    .B(_1416_),
    .X(_1419_));
 sky130_fd_sc_hd__a2111o_1 _3089_ (.A1(_1260_),
    .A2(_1394_),
    .B1(_1412_),
    .C1(_1413_),
    .D1(_1418_),
    .X(_1420_));
 sky130_fd_sc_hd__and3b_1 _3090_ (.A_N(_1420_),
    .B(_1419_),
    .C(_1411_),
    .X(_1421_));
 sky130_fd_sc_hd__a211o_1 _3091_ (.A1(net744),
    .A2(_1420_),
    .B1(_1421_),
    .C1(net91),
    .X(_0151_));
 sky130_fd_sc_hd__nand2_1 _3092_ (.A(_1763_),
    .B(\mem_cycle[4] ),
    .Y(_1422_));
 sky130_fd_sc_hd__or3_1 _3093_ (.A(\mem_cycle[3] ),
    .B(_1765_),
    .C(_1264_),
    .X(_1423_));
 sky130_fd_sc_hd__o211a_1 _3094_ (.A1(\mem_cycle[0] ),
    .A2(_1373_),
    .B1(_1422_),
    .C1(_1423_),
    .X(_1424_));
 sky130_fd_sc_hd__or4b_1 _3095_ (.A(\mem_cycle[5] ),
    .B(\mem_cycle[4] ),
    .C(\mem_cycle[0] ),
    .D_N(\mem_cycle[3] ),
    .X(_1425_));
 sky130_fd_sc_hd__or4_1 _3096_ (.A(\mem_cycle[1] ),
    .B(\mem_cycle[0] ),
    .C(_1263_),
    .D(_1422_),
    .X(_1426_));
 sky130_fd_sc_hd__inv_2 _3097_ (.A(_1426_),
    .Y(_1427_));
 sky130_fd_sc_hd__o211a_1 _3098_ (.A1(_1765_),
    .A2(_1414_),
    .B1(_1425_),
    .C1(_1426_),
    .X(_1428_));
 sky130_fd_sc_hd__or3_1 _3099_ (.A(_1763_),
    .B(\mem_cycle[4] ),
    .C(_1263_),
    .X(_1429_));
 sky130_fd_sc_hd__nor3_1 _3100_ (.A(net796),
    .B(_1766_),
    .C(_1429_),
    .Y(_1430_));
 sky130_fd_sc_hd__a31oi_1 _3101_ (.A1(_1763_),
    .A2(net835),
    .A3(_1373_),
    .B1(_1430_),
    .Y(_1431_));
 sky130_fd_sc_hd__and4_1 _3102_ (.A(_1405_),
    .B(_1424_),
    .C(_1428_),
    .D(_1431_),
    .X(_1432_));
 sky130_fd_sc_hd__o311a_1 _3103_ (.A1(_1265_),
    .A2(_1394_),
    .A3(_1432_),
    .B1(_1260_),
    .C1(net64),
    .X(_1433_));
 sky130_fd_sc_hd__or3b_1 _3104_ (.A(\startup_cycle[6] ),
    .B(net722),
    .C_N(net698),
    .X(_1434_));
 sky130_fd_sc_hd__or2_1 _3105_ (.A(_1258_),
    .B(_1434_),
    .X(_1435_));
 sky130_fd_sc_hd__nand2_2 _3106_ (.A(_1767_),
    .B(net722),
    .Y(_1436_));
 sky130_fd_sc_hd__a31o_1 _3107_ (.A1(_1409_),
    .A2(_1435_),
    .A3(_1436_),
    .B1(_1255_),
    .X(_1437_));
 sky130_fd_sc_hd__nand2b_1 _3108_ (.A_N(_1409_),
    .B(_1307_),
    .Y(_1438_));
 sky130_fd_sc_hd__a31o_1 _3109_ (.A1(_1434_),
    .A2(_1436_),
    .A3(_1438_),
    .B1(_1311_),
    .X(_1439_));
 sky130_fd_sc_hd__a311o_1 _3110_ (.A1(_1332_),
    .A2(_1437_),
    .A3(_1439_),
    .B1(_1433_),
    .C1(_1306_),
    .X(_1440_));
 sky130_fd_sc_hd__a21oi_1 _3111_ (.A1(_1260_),
    .A2(_1431_),
    .B1(_1253_),
    .Y(_1441_));
 sky130_fd_sc_hd__a2bb2o_1 _3112_ (.A1_N(net820),
    .A2_N(net64),
    .B1(_1437_),
    .B2(_1441_),
    .X(_1442_));
 sky130_fd_sc_hd__mux2_1 _3113_ (.A0(_1442_),
    .A1(net846),
    .S(_1440_),
    .X(_1443_));
 sky130_fd_sc_hd__and2_1 _3114_ (.A(net94),
    .B(net847),
    .X(_0152_));
 sky130_fd_sc_hd__nand2b_1 _3115_ (.A_N(_1417_),
    .B(_1428_),
    .Y(_1444_));
 sky130_fd_sc_hd__a21o_1 _3116_ (.A1(_1266_),
    .A2(_1444_),
    .B1(_1262_),
    .X(_1445_));
 sky130_fd_sc_hd__a21o_1 _3117_ (.A1(net726),
    .A2(net820),
    .B1(net64),
    .X(_1446_));
 sky130_fd_sc_hd__or4_1 _3118_ (.A(\startup_cycle[6] ),
    .B(net722),
    .C(_1255_),
    .D(_1259_),
    .X(_1447_));
 sky130_fd_sc_hd__or3_1 _3119_ (.A(net698),
    .B(_1407_),
    .C(_1436_),
    .X(_1448_));
 sky130_fd_sc_hd__nor4_1 _3120_ (.A(net698),
    .B(_1255_),
    .C(_1307_),
    .D(_1436_),
    .Y(_1449_));
 sky130_fd_sc_hd__nand3b_1 _3121_ (.A_N(_1449_),
    .B(_1447_),
    .C(_1448_),
    .Y(_1450_));
 sky130_fd_sc_hd__o311a_1 _3122_ (.A1(_1253_),
    .A2(_1260_),
    .A3(_1450_),
    .B1(_1446_),
    .C1(_1445_),
    .X(_1451_));
 sky130_fd_sc_hd__nand2_1 _3123_ (.A(net830),
    .B(_1765_),
    .Y(_1452_));
 sky130_fd_sc_hd__nor2_1 _3124_ (.A(_1264_),
    .B(_1452_),
    .Y(_1453_));
 sky130_fd_sc_hd__nor2_1 _3125_ (.A(_1414_),
    .B(_1452_),
    .Y(_1454_));
 sky130_fd_sc_hd__a221o_1 _3126_ (.A1(\ROM_addr_buff[8] ),
    .A2(_1453_),
    .B1(_1454_),
    .B2(\ROM_addr_buff[4] ),
    .C1(_1427_),
    .X(_1455_));
 sky130_fd_sc_hd__a31o_1 _3127_ (.A1(\ROM_addr_buff[12] ),
    .A2(_1416_),
    .A3(_1425_),
    .B1(_1455_),
    .X(_1456_));
 sky130_fd_sc_hd__a211o_1 _3128_ (.A1(_1260_),
    .A2(_1456_),
    .B1(_1449_),
    .C1(_1253_),
    .X(_1457_));
 sky130_fd_sc_hd__o21a_1 _3129_ (.A1(net423),
    .A2(net821),
    .B1(_1457_),
    .X(_1458_));
 sky130_fd_sc_hd__mux2_1 _3130_ (.A0(net833),
    .A1(_1458_),
    .S(_1451_),
    .X(_1459_));
 sky130_fd_sc_hd__and2_1 _3131_ (.A(net93),
    .B(net834),
    .X(_0153_));
 sky130_fd_sc_hd__nor2_1 _3132_ (.A(_1292_),
    .B(_1422_),
    .Y(_1460_));
 sky130_fd_sc_hd__nor2_1 _3133_ (.A(_1417_),
    .B(_1460_),
    .Y(_1461_));
 sky130_fd_sc_hd__nand3_1 _3134_ (.A(\startup_cycle[4] ),
    .B(_1254_),
    .C(_1258_),
    .Y(_1462_));
 sky130_fd_sc_hd__o21a_1 _3135_ (.A1(_1436_),
    .A2(_1462_),
    .B1(_1447_),
    .X(_1463_));
 sky130_fd_sc_hd__or3_1 _3136_ (.A(_1413_),
    .B(_1461_),
    .C(_1463_),
    .X(_1464_));
 sky130_fd_sc_hd__o2bb2a_1 _3137_ (.A1_N(_1260_),
    .A2_N(_1460_),
    .B1(_1462_),
    .B2(_1436_),
    .X(_1465_));
 sky130_fd_sc_hd__nor2_1 _3138_ (.A(_1464_),
    .B(_1465_),
    .Y(_1466_));
 sky130_fd_sc_hd__a211o_1 _3139_ (.A1(net447),
    .A2(_1464_),
    .B1(_1466_),
    .C1(net91),
    .X(_0154_));
 sky130_fd_sc_hd__or4_1 _3140_ (.A(_1253_),
    .B(_1255_),
    .C(_1259_),
    .D(_1434_),
    .X(_1467_));
 sky130_fd_sc_hd__a21o_1 _3141_ (.A1(net214),
    .A2(_1467_),
    .B1(net91),
    .X(_0155_));
 sky130_fd_sc_hd__o21a_2 _3142_ (.A1(\ROM_spi_cycle[0] ),
    .A2(net64),
    .B1(_1320_),
    .X(_1468_));
 sky130_fd_sc_hd__o21ai_4 _3143_ (.A1(\ROM_spi_cycle[0] ),
    .A2(net64),
    .B1(_1320_),
    .Y(_1469_));
 sky130_fd_sc_hd__a21o_1 _3144_ (.A1(_1256_),
    .A2(_1313_),
    .B1(_1317_),
    .X(_1470_));
 sky130_fd_sc_hd__a21o_1 _3145_ (.A1(net64),
    .A2(_1470_),
    .B1(_1469_),
    .X(_1471_));
 sky130_fd_sc_hd__o211a_1 _3146_ (.A1(net392),
    .A2(_1468_),
    .B1(_1471_),
    .C1(net93),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _3147_ (.A0(net392),
    .A1(_1311_),
    .S(net64),
    .X(_1472_));
 sky130_fd_sc_hd__or2_1 _3148_ (.A(_1469_),
    .B(_1472_),
    .X(_1473_));
 sky130_fd_sc_hd__o211a_1 _3149_ (.A1(net409),
    .A2(_1468_),
    .B1(_1473_),
    .C1(net93),
    .X(_0157_));
 sky130_fd_sc_hd__nor2_1 _3150_ (.A(_1253_),
    .B(_1315_),
    .Y(_1474_));
 sky130_fd_sc_hd__a211o_1 _3151_ (.A1(net409),
    .A2(_1253_),
    .B1(_1469_),
    .C1(_1474_),
    .X(_1475_));
 sky130_fd_sc_hd__o211a_1 _3152_ (.A1(net417),
    .A2(_1468_),
    .B1(_1475_),
    .C1(net93),
    .X(_0158_));
 sky130_fd_sc_hd__a21oi_1 _3153_ (.A1(_1256_),
    .A2(_1310_),
    .B1(_1317_),
    .Y(_1476_));
 sky130_fd_sc_hd__nor2_1 _3154_ (.A(_1253_),
    .B(_1476_),
    .Y(_1477_));
 sky130_fd_sc_hd__a211o_1 _3155_ (.A1(\ROM_spi_dat_out[2] ),
    .A2(_1253_),
    .B1(_1469_),
    .C1(_1477_),
    .X(_1478_));
 sky130_fd_sc_hd__o211a_1 _3156_ (.A1(net413),
    .A2(_1468_),
    .B1(_1478_),
    .C1(net93),
    .X(_0159_));
 sky130_fd_sc_hd__or2_1 _3157_ (.A(_1253_),
    .B(_1317_),
    .X(_1479_));
 sky130_fd_sc_hd__o21ai_1 _3158_ (.A1(net413),
    .A2(net64),
    .B1(_1479_),
    .Y(_1480_));
 sky130_fd_sc_hd__nand2_1 _3159_ (.A(_1468_),
    .B(_1480_),
    .Y(_1481_));
 sky130_fd_sc_hd__o211a_1 _3160_ (.A1(net419),
    .A2(_1468_),
    .B1(_1481_),
    .C1(net93),
    .X(_0160_));
 sky130_fd_sc_hd__a211o_1 _3161_ (.A1(\ROM_spi_dat_out[4] ),
    .A2(_1253_),
    .B1(_1469_),
    .C1(_1477_),
    .X(_1482_));
 sky130_fd_sc_hd__o211a_1 _3162_ (.A1(net415),
    .A2(_1468_),
    .B1(_1482_),
    .C1(net93),
    .X(_0161_));
 sky130_fd_sc_hd__and2_1 _3163_ (.A(_1256_),
    .B(_1309_),
    .X(_1483_));
 sky130_fd_sc_hd__o22a_1 _3164_ (.A1(net415),
    .A2(net64),
    .B1(_1479_),
    .B2(_1483_),
    .X(_1484_));
 sky130_fd_sc_hd__or2_1 _3165_ (.A(net500),
    .B(_1468_),
    .X(_1485_));
 sky130_fd_sc_hd__o211a_1 _3166_ (.A1(_1469_),
    .A2(_1484_),
    .B1(net501),
    .C1(net93),
    .X(_0162_));
 sky130_fd_sc_hd__a211o_1 _3167_ (.A1(\ROM_spi_dat_out[6] ),
    .A2(_1253_),
    .B1(_1469_),
    .C1(_1477_),
    .X(_1486_));
 sky130_fd_sc_hd__o211a_1 _3168_ (.A1(net423),
    .A2(_1468_),
    .B1(_1486_),
    .C1(net93),
    .X(_0163_));
 sky130_fd_sc_hd__nor2_2 _3169_ (.A(_1262_),
    .B(_1265_),
    .Y(_1487_));
 sky130_fd_sc_hd__and2_1 _3170_ (.A(_1374_),
    .B(_1487_),
    .X(_1488_));
 sky130_fd_sc_hd__nand2_8 _3171_ (.A(_1374_),
    .B(_1487_),
    .Y(_1489_));
 sky130_fd_sc_hd__a21o_1 _3172_ (.A1(net124),
    .A2(_1489_),
    .B1(net91),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _3173_ (.A0(net780),
    .A1(\last_addr[1] ),
    .S(_1489_),
    .X(_1490_));
 sky130_fd_sc_hd__or2_1 _3174_ (.A(net92),
    .B(net781),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _3175_ (.A0(\ROM_addr_buff[2] ),
    .A1(net802),
    .S(_1489_),
    .X(_1491_));
 sky130_fd_sc_hd__or2_1 _3176_ (.A(net92),
    .B(net803),
    .X(_0166_));
 sky130_fd_sc_hd__or2_1 _3177_ (.A(net696),
    .B(_1488_),
    .X(_1492_));
 sky130_fd_sc_hd__o211a_1 _3178_ (.A1(net692),
    .A2(_1489_),
    .B1(_1492_),
    .C1(net95),
    .X(_0167_));
 sky130_fd_sc_hd__or2_1 _3179_ (.A(net762),
    .B(_1488_),
    .X(_1493_));
 sky130_fd_sc_hd__o211a_1 _3180_ (.A1(net758),
    .A2(_1489_),
    .B1(_1493_),
    .C1(net95),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _3181_ (.A0(\ROM_addr_buff[5] ),
    .A1(net674),
    .S(_1489_),
    .X(_1494_));
 sky130_fd_sc_hd__or2_1 _3182_ (.A(net92),
    .B(net675),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _3183_ (.A0(net766),
    .A1(net798),
    .S(_1489_),
    .X(_1495_));
 sky130_fd_sc_hd__or2_1 _3184_ (.A(net91),
    .B(net799),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _3185_ (.A0(\ROM_addr_buff[7] ),
    .A1(net711),
    .S(_1489_),
    .X(_1496_));
 sky130_fd_sc_hd__or2_1 _3186_ (.A(net91),
    .B(net712),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _3187_ (.A0(net736),
    .A1(net791),
    .S(_1489_),
    .X(_1497_));
 sky130_fd_sc_hd__or2_1 _3188_ (.A(net91),
    .B(net792),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _3189_ (.A0(\ROM_addr_buff[9] ),
    .A1(net670),
    .S(_1489_),
    .X(_1498_));
 sky130_fd_sc_hd__or2_1 _3190_ (.A(net91),
    .B(net671),
    .X(_0173_));
 sky130_fd_sc_hd__or2_1 _3191_ (.A(net682),
    .B(_1488_),
    .X(_1499_));
 sky130_fd_sc_hd__o211a_1 _3192_ (.A1(net850),
    .A2(_1489_),
    .B1(_1499_),
    .C1(net93),
    .X(_0174_));
 sky130_fd_sc_hd__or2_1 _3193_ (.A(net774),
    .B(_1488_),
    .X(_1500_));
 sky130_fd_sc_hd__o211a_1 _3194_ (.A1(net718),
    .A2(_1489_),
    .B1(_1500_),
    .C1(net93),
    .X(_0175_));
 sky130_fd_sc_hd__or2_1 _3195_ (.A(net716),
    .B(_1488_),
    .X(_1501_));
 sky130_fd_sc_hd__o211a_1 _3196_ (.A1(\ROM_addr_buff[12] ),
    .A2(_1489_),
    .B1(_1501_),
    .C1(net94),
    .X(_0176_));
 sky130_fd_sc_hd__or2_1 _3197_ (.A(\last_addr[13] ),
    .B(_1488_),
    .X(_1502_));
 sky130_fd_sc_hd__o211a_1 _3198_ (.A1(net738),
    .A2(_1489_),
    .B1(_1502_),
    .C1(net95),
    .X(_0177_));
 sky130_fd_sc_hd__and2_1 _3199_ (.A(net726),
    .B(net64),
    .X(_1503_));
 sky130_fd_sc_hd__o21a_1 _3200_ (.A1(_1306_),
    .A2(_1503_),
    .B1(net94),
    .X(_0178_));
 sky130_fd_sc_hd__nand2_2 _3201_ (.A(_1836_),
    .B(_1296_),
    .Y(_1504_));
 sky130_fd_sc_hd__a31o_1 _3202_ (.A1(net35),
    .A2(_1836_),
    .A3(_0448_),
    .B1(net516),
    .X(_1505_));
 sky130_fd_sc_hd__o211a_1 _3203_ (.A1(\S8x305.iv_latch[0] ),
    .A2(_1504_),
    .B1(_1505_),
    .C1(net99),
    .X(_0179_));
 sky130_fd_sc_hd__a31o_1 _3204_ (.A1(net35),
    .A2(_1836_),
    .A3(_0448_),
    .B1(net486),
    .X(_1506_));
 sky130_fd_sc_hd__o211a_1 _3205_ (.A1(net851),
    .A2(_1504_),
    .B1(_1506_),
    .C1(net99),
    .X(_0180_));
 sky130_fd_sc_hd__a31o_1 _3206_ (.A1(net35),
    .A2(_1836_),
    .A3(_0448_),
    .B1(net461),
    .X(_1507_));
 sky130_fd_sc_hd__o211a_1 _3207_ (.A1(\S8x305.iv_latch[2] ),
    .A2(_1504_),
    .B1(_1507_),
    .C1(net99),
    .X(_0181_));
 sky130_fd_sc_hd__a31o_1 _3208_ (.A1(net35),
    .A2(_1836_),
    .A3(_0448_),
    .B1(net496),
    .X(_1508_));
 sky130_fd_sc_hd__o211a_1 _3209_ (.A1(\S8x305.iv_latch[3] ),
    .A2(_1504_),
    .B1(_1508_),
    .C1(net99),
    .X(_0182_));
 sky130_fd_sc_hd__a31o_1 _3210_ (.A1(net35),
    .A2(_1836_),
    .A3(_0448_),
    .B1(net481),
    .X(_1509_));
 sky130_fd_sc_hd__o211a_1 _3211_ (.A1(\S8x305.iv_latch[4] ),
    .A2(_1504_),
    .B1(_1509_),
    .C1(net99),
    .X(_0183_));
 sky130_fd_sc_hd__a31o_1 _3212_ (.A1(net35),
    .A2(_1836_),
    .A3(_0448_),
    .B1(net457),
    .X(_1510_));
 sky130_fd_sc_hd__o211a_1 _3213_ (.A1(net429),
    .A2(_1504_),
    .B1(_1510_),
    .C1(net100),
    .X(_0184_));
 sky130_fd_sc_hd__a31o_1 _3214_ (.A1(net35),
    .A2(_1836_),
    .A3(_0448_),
    .B1(net435),
    .X(_1511_));
 sky130_fd_sc_hd__o211a_1 _3215_ (.A1(net400),
    .A2(_1504_),
    .B1(_1511_),
    .C1(net100),
    .X(_0185_));
 sky130_fd_sc_hd__a31o_1 _3216_ (.A1(net35),
    .A2(_1836_),
    .A3(_0448_),
    .B1(net466),
    .X(_1512_));
 sky130_fd_sc_hd__o211a_1 _3217_ (.A1(\S8x305.iv_latch[7] ),
    .A2(_1504_),
    .B1(_1512_),
    .C1(net100),
    .X(_0186_));
 sky130_fd_sc_hd__or2_1 _3218_ (.A(net505),
    .B(_1129_),
    .X(_1513_));
 sky130_fd_sc_hd__o211a_1 _3219_ (.A1(\S8x305.iv_latch[4] ),
    .A2(_1130_),
    .B1(_1513_),
    .C1(net99),
    .X(_0191_));
 sky130_fd_sc_hd__or2_1 _3220_ (.A(\cmdr[5] ),
    .B(_1129_),
    .X(_1514_));
 sky130_fd_sc_hd__o211a_1 _3221_ (.A1(net429),
    .A2(_1130_),
    .B1(_1514_),
    .C1(net99),
    .X(_0192_));
 sky130_fd_sc_hd__or2_1 _3222_ (.A(net439),
    .B(_1129_),
    .X(_1515_));
 sky130_fd_sc_hd__o211a_1 _3223_ (.A1(net400),
    .A2(_1130_),
    .B1(_1515_),
    .C1(net99),
    .X(_0193_));
 sky130_fd_sc_hd__or2_1 _3224_ (.A(net475),
    .B(_1129_),
    .X(_1516_));
 sky130_fd_sc_hd__o211a_1 _3225_ (.A1(\S8x305.iv_latch[7] ),
    .A2(_1130_),
    .B1(_1516_),
    .C1(net99),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _3226_ (.A0(_1749_),
    .A1(_1762_),
    .S(net57),
    .X(_1517_));
 sky130_fd_sc_hd__nand2_1 _3227_ (.A(net103),
    .B(net752),
    .Y(_0195_));
 sky130_fd_sc_hd__mux2_1 _3228_ (.A0(_1748_),
    .A1(_1761_),
    .S(net58),
    .X(_1518_));
 sky130_fd_sc_hd__nand2_1 _3229_ (.A(net95),
    .B(net456),
    .Y(_0196_));
 sky130_fd_sc_hd__mux2_1 _3230_ (.A0(_1747_),
    .A1(_1760_),
    .S(net57),
    .X(_1519_));
 sky130_fd_sc_hd__nand2_1 _3231_ (.A(net95),
    .B(net544),
    .Y(_0197_));
 sky130_fd_sc_hd__mux2_1 _3232_ (.A0(_1746_),
    .A1(_1759_),
    .S(net58),
    .X(_1520_));
 sky130_fd_sc_hd__nand2_1 _3233_ (.A(net95),
    .B(net484),
    .Y(_0198_));
 sky130_fd_sc_hd__mux2_1 _3234_ (.A0(_1745_),
    .A1(_1758_),
    .S(net57),
    .X(_1521_));
 sky130_fd_sc_hd__nand2_1 _3235_ (.A(net95),
    .B(net640),
    .Y(_0199_));
 sky130_fd_sc_hd__mux2_1 _3236_ (.A0(net753),
    .A1(\last_A[6] ),
    .S(net58),
    .X(_1522_));
 sky130_fd_sc_hd__or2_1 _3237_ (.A(net92),
    .B(net754),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _3238_ (.A0(net672),
    .A1(\last_A[7] ),
    .S(net57),
    .X(_1523_));
 sky130_fd_sc_hd__or2_1 _3239_ (.A(net92),
    .B(net673),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _3240_ (.A0(_1742_),
    .A1(_1757_),
    .S(net57),
    .X(_1524_));
 sky130_fd_sc_hd__nand2_1 _3241_ (.A(net96),
    .B(net495),
    .Y(_0202_));
 sky130_fd_sc_hd__mux2_1 _3242_ (.A0(_1741_),
    .A1(_1756_),
    .S(net58),
    .X(_1525_));
 sky130_fd_sc_hd__nand2_1 _3243_ (.A(net96),
    .B(net454),
    .Y(_0203_));
 sky130_fd_sc_hd__mux2_1 _3244_ (.A0(\S8x305.A[11] ),
    .A1(net724),
    .S(net58),
    .X(_1526_));
 sky130_fd_sc_hd__or2_1 _3245_ (.A(net92),
    .B(net725),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _3246_ (.A0(\S8x305.A[12] ),
    .A1(net708),
    .S(net57),
    .X(_1527_));
 sky130_fd_sc_hd__or2_1 _3247_ (.A(net92),
    .B(net709),
    .X(_0205_));
 sky130_fd_sc_hd__or3b_4 _3248_ (.A(_1064_),
    .B(\cmdr[1] ),
    .C_N(\cmdr[0] ),
    .X(_1528_));
 sky130_fd_sc_hd__mux2_1 _3249_ (.A0(net81),
    .A1(net194),
    .S(_1528_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _3250_ (.A0(net80),
    .A1(net368),
    .S(_1528_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _3251_ (.A0(net79),
    .A1(net298),
    .S(_1528_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _3252_ (.A0(net78),
    .A1(net134),
    .S(_1528_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _3253_ (.A0(net77),
    .A1(net138),
    .S(_1528_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _3254_ (.A0(net76),
    .A1(net150),
    .S(_1528_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_1 _3255_ (.A0(net75),
    .A1(net240),
    .S(_1528_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _3256_ (.A0(net74),
    .A1(net254),
    .S(_1528_),
    .X(_0213_));
 sky130_fd_sc_hd__nor2_2 _3257_ (.A(_1108_),
    .B(_1147_),
    .Y(_1529_));
 sky130_fd_sc_hd__or2_2 _3258_ (.A(_1108_),
    .B(_1147_),
    .X(_1530_));
 sky130_fd_sc_hd__and3_1 _3259_ (.A(net109),
    .B(net561),
    .C(_1530_),
    .X(_1531_));
 sky130_fd_sc_hd__a21o_1 _3260_ (.A1(_1112_),
    .A2(_1529_),
    .B1(_1531_),
    .X(_0214_));
 sky130_fd_sc_hd__and3_1 _3261_ (.A(net109),
    .B(net522),
    .C(_1530_),
    .X(_1532_));
 sky130_fd_sc_hd__a21o_1 _3262_ (.A1(_1114_),
    .A2(_1529_),
    .B1(_1532_),
    .X(_0215_));
 sky130_fd_sc_hd__and3_1 _3263_ (.A(net109),
    .B(net645),
    .C(_1530_),
    .X(_1533_));
 sky130_fd_sc_hd__a21o_1 _3264_ (.A1(_1116_),
    .A2(_1529_),
    .B1(_1533_),
    .X(_0216_));
 sky130_fd_sc_hd__and3_1 _3265_ (.A(net109),
    .B(net637),
    .C(_1530_),
    .X(_1534_));
 sky130_fd_sc_hd__a21o_1 _3266_ (.A1(_1118_),
    .A2(_1529_),
    .B1(_1534_),
    .X(_0217_));
 sky130_fd_sc_hd__and3_1 _3267_ (.A(net109),
    .B(net595),
    .C(_1530_),
    .X(_1535_));
 sky130_fd_sc_hd__a21o_1 _3268_ (.A1(_1120_),
    .A2(_1529_),
    .B1(_1535_),
    .X(_0218_));
 sky130_fd_sc_hd__and3_1 _3269_ (.A(net109),
    .B(net564),
    .C(_1530_),
    .X(_1536_));
 sky130_fd_sc_hd__a21o_1 _3270_ (.A1(_1123_),
    .A2(_1529_),
    .B1(_1536_),
    .X(_0219_));
 sky130_fd_sc_hd__and3_1 _3271_ (.A(net110),
    .B(net614),
    .C(_1530_),
    .X(_1537_));
 sky130_fd_sc_hd__a21o_1 _3272_ (.A1(_1125_),
    .A2(_1529_),
    .B1(_1537_),
    .X(_0220_));
 sky130_fd_sc_hd__and3_1 _3273_ (.A(net110),
    .B(net557),
    .C(_1530_),
    .X(_1538_));
 sky130_fd_sc_hd__a21o_1 _3274_ (.A1(_1128_),
    .A2(_1529_),
    .B1(_1538_),
    .X(_0221_));
 sky130_fd_sc_hd__or3_1 _3275_ (.A(net826),
    .B(_1764_),
    .C(_1262_),
    .X(_1539_));
 sky130_fd_sc_hd__or3_2 _3276_ (.A(_1283_),
    .B(_1452_),
    .C(_1539_),
    .X(_1540_));
 sky130_fd_sc_hd__mux2_1 _3277_ (.A0(net4),
    .A1(net804),
    .S(_1540_),
    .X(_1541_));
 sky130_fd_sc_hd__and2_1 _3278_ (.A(net97),
    .B(_1541_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _3279_ (.A0(net5),
    .A1(net755),
    .S(_1540_),
    .X(_1542_));
 sky130_fd_sc_hd__and2_1 _3280_ (.A(net99),
    .B(net756),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _3281_ (.A0(net6),
    .A1(net663),
    .S(_1540_),
    .X(_1543_));
 sky130_fd_sc_hd__and2_1 _3282_ (.A(net97),
    .B(net664),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _3283_ (.A0(net7),
    .A1(net782),
    .S(_1540_),
    .X(_1544_));
 sky130_fd_sc_hd__and2_1 _3284_ (.A(net99),
    .B(net783),
    .X(_0225_));
 sky130_fd_sc_hd__or4_4 _3285_ (.A(\mem_cycle[1] ),
    .B(_1766_),
    .C(_1285_),
    .D(_1539_),
    .X(_1545_));
 sky130_fd_sc_hd__mux2_1 _3286_ (.A0(net4),
    .A1(net678),
    .S(_1545_),
    .X(_1546_));
 sky130_fd_sc_hd__and2_1 _3287_ (.A(net97),
    .B(net679),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _3288_ (.A0(net5),
    .A1(net748),
    .S(_1545_),
    .X(_1547_));
 sky130_fd_sc_hd__and2_1 _3289_ (.A(net97),
    .B(net749),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _3290_ (.A0(net6),
    .A1(net676),
    .S(_1545_),
    .X(_1548_));
 sky130_fd_sc_hd__and2_1 _3291_ (.A(net98),
    .B(net677),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _3292_ (.A0(net7),
    .A1(net776),
    .S(_1545_),
    .X(_1549_));
 sky130_fd_sc_hd__and2_1 _3293_ (.A(net98),
    .B(net777),
    .X(_0229_));
 sky130_fd_sc_hd__nand2_2 _3294_ (.A(net797),
    .B(_1487_),
    .Y(_1550_));
 sky130_fd_sc_hd__mux2_1 _3295_ (.A0(net4),
    .A1(net772),
    .S(_1550_),
    .X(_1551_));
 sky130_fd_sc_hd__and2_1 _3296_ (.A(net97),
    .B(_1551_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _3297_ (.A0(net5),
    .A1(net746),
    .S(_1550_),
    .X(_1552_));
 sky130_fd_sc_hd__and2_1 _3298_ (.A(net97),
    .B(net747),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _3299_ (.A0(net6),
    .A1(net732),
    .S(_1550_),
    .X(_1553_));
 sky130_fd_sc_hd__and2_1 _3300_ (.A(net97),
    .B(net733),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _3301_ (.A0(net7),
    .A1(net794),
    .S(_1550_),
    .X(_1554_));
 sky130_fd_sc_hd__and2_1 _3302_ (.A(net97),
    .B(net795),
    .X(_0233_));
 sky130_fd_sc_hd__o211a_1 _3303_ (.A1(net738),
    .A2(\mem_cycle[3] ),
    .B1(net443),
    .C1(_1415_),
    .X(_1555_));
 sky130_fd_sc_hd__nor2_1 _3304_ (.A(_1264_),
    .B(_1285_),
    .Y(_1556_));
 sky130_fd_sc_hd__a22o_1 _3305_ (.A1(\ROM_addr_buff[9] ),
    .A2(_1453_),
    .B1(_1556_),
    .B2(\ROM_addr_buff[1] ),
    .X(_1557_));
 sky130_fd_sc_hd__a211o_1 _3306_ (.A1(net761),
    .A2(_1454_),
    .B1(_1555_),
    .C1(_1557_),
    .X(_1558_));
 sky130_fd_sc_hd__and3b_1 _3307_ (.A_N(_1413_),
    .B(_1444_),
    .C(_1450_),
    .X(_1559_));
 sky130_fd_sc_hd__nand2_1 _3308_ (.A(_1448_),
    .B(_1559_),
    .Y(_1560_));
 sky130_fd_sc_hd__a21o_1 _3309_ (.A1(_1260_),
    .A2(_1558_),
    .B1(_1560_),
    .X(_1561_));
 sky130_fd_sc_hd__o211a_1 _3310_ (.A1(net778),
    .A2(_1559_),
    .B1(_1561_),
    .C1(net94),
    .X(_0234_));
 sky130_fd_sc_hd__a22o_1 _3311_ (.A1(net767),
    .A2(_1453_),
    .B1(_1556_),
    .B2(\ROM_addr_buff[2] ),
    .X(_1562_));
 sky130_fd_sc_hd__a211o_1 _3312_ (.A1(net766),
    .A2(_1454_),
    .B1(_1562_),
    .C1(_1427_),
    .X(_1563_));
 sky130_fd_sc_hd__a21o_1 _3313_ (.A1(_1260_),
    .A2(_1563_),
    .B1(_1449_),
    .X(_1564_));
 sky130_fd_sc_hd__mux2_1 _3314_ (.A0(net828),
    .A1(_1564_),
    .S(_1559_),
    .X(_1565_));
 sky130_fd_sc_hd__or2_1 _3315_ (.A(net91),
    .B(net829),
    .X(_0235_));
 sky130_fd_sc_hd__o211a_1 _3316_ (.A1(net790),
    .A2(net443),
    .B1(_1415_),
    .C1(net830),
    .X(_1566_));
 sky130_fd_sc_hd__a22o_1 _3317_ (.A1(net718),
    .A2(_1453_),
    .B1(_1556_),
    .B2(net692),
    .X(_1567_));
 sky130_fd_sc_hd__o21a_1 _3318_ (.A1(_1566_),
    .A2(_1567_),
    .B1(_1260_),
    .X(_1568_));
 sky130_fd_sc_hd__o22a_1 _3319_ (.A1(net839),
    .A2(_1559_),
    .B1(_1560_),
    .B2(_1568_),
    .X(_1569_));
 sky130_fd_sc_hd__or2_1 _3320_ (.A(net91),
    .B(net840),
    .X(_0236_));
 sky130_fd_sc_hd__nor2_1 _3321_ (.A(_1830_),
    .B(_0437_),
    .Y(_1570_));
 sky130_fd_sc_hd__and3_2 _3322_ (.A(_1816_),
    .B(_1107_),
    .C(_1570_),
    .X(_1571_));
 sky130_fd_sc_hd__or3b_4 _3323_ (.A(_1817_),
    .B(_1106_),
    .C_N(_1570_),
    .X(_1572_));
 sky130_fd_sc_hd__and3_1 _3324_ (.A(net111),
    .B(net643),
    .C(_1572_),
    .X(_1573_));
 sky130_fd_sc_hd__a21o_1 _3325_ (.A1(_1112_),
    .A2(_1571_),
    .B1(_1573_),
    .X(_0237_));
 sky130_fd_sc_hd__and3_1 _3326_ (.A(net112),
    .B(net627),
    .C(_1572_),
    .X(_1574_));
 sky130_fd_sc_hd__a21o_1 _3327_ (.A1(_1114_),
    .A2(_1571_),
    .B1(_1574_),
    .X(_0238_));
 sky130_fd_sc_hd__and3_1 _3328_ (.A(net112),
    .B(net632),
    .C(_1572_),
    .X(_1575_));
 sky130_fd_sc_hd__a21o_1 _3329_ (.A1(_1116_),
    .A2(_1571_),
    .B1(_1575_),
    .X(_0239_));
 sky130_fd_sc_hd__and3_1 _3330_ (.A(net111),
    .B(net587),
    .C(_1572_),
    .X(_1576_));
 sky130_fd_sc_hd__a21o_1 _3331_ (.A1(_1118_),
    .A2(_1571_),
    .B1(_1576_),
    .X(_0240_));
 sky130_fd_sc_hd__and3_1 _3332_ (.A(net111),
    .B(net536),
    .C(_1572_),
    .X(_1577_));
 sky130_fd_sc_hd__a21o_1 _3333_ (.A1(_1120_),
    .A2(_1571_),
    .B1(_1577_),
    .X(_0241_));
 sky130_fd_sc_hd__and3_1 _3334_ (.A(net111),
    .B(net582),
    .C(_1572_),
    .X(_1578_));
 sky130_fd_sc_hd__a21o_1 _3335_ (.A1(_1123_),
    .A2(_1571_),
    .B1(_1578_),
    .X(_0242_));
 sky130_fd_sc_hd__and3_1 _3336_ (.A(net111),
    .B(net570),
    .C(_1572_),
    .X(_1579_));
 sky130_fd_sc_hd__a21o_1 _3337_ (.A1(_1125_),
    .A2(_1571_),
    .B1(_1579_),
    .X(_0243_));
 sky130_fd_sc_hd__and3_1 _3338_ (.A(net110),
    .B(net659),
    .C(_1572_),
    .X(_1580_));
 sky130_fd_sc_hd__a21o_1 _3339_ (.A1(_1128_),
    .A2(_1571_),
    .B1(_1580_),
    .X(_0244_));
 sky130_fd_sc_hd__and3_2 _3340_ (.A(_0444_),
    .B(_1107_),
    .C(_1570_),
    .X(_1581_));
 sky130_fd_sc_hd__or3b_4 _3341_ (.A(_0445_),
    .B(_1106_),
    .C_N(_1570_),
    .X(_1582_));
 sky130_fd_sc_hd__and3_1 _3342_ (.A(net112),
    .B(net519),
    .C(_1582_),
    .X(_1583_));
 sky130_fd_sc_hd__a21o_1 _3343_ (.A1(_1112_),
    .A2(_1581_),
    .B1(_1583_),
    .X(_0245_));
 sky130_fd_sc_hd__and3_1 _3344_ (.A(net112),
    .B(net523),
    .C(_1582_),
    .X(_1584_));
 sky130_fd_sc_hd__a21o_1 _3345_ (.A1(_1114_),
    .A2(_1581_),
    .B1(_1584_),
    .X(_0246_));
 sky130_fd_sc_hd__and3_1 _3346_ (.A(net110),
    .B(net610),
    .C(_1582_),
    .X(_1585_));
 sky130_fd_sc_hd__a21o_1 _3347_ (.A1(_1116_),
    .A2(_1581_),
    .B1(_1585_),
    .X(_0247_));
 sky130_fd_sc_hd__and3_1 _3348_ (.A(net112),
    .B(net485),
    .C(_1582_),
    .X(_1586_));
 sky130_fd_sc_hd__a21o_1 _3349_ (.A1(_1118_),
    .A2(_1581_),
    .B1(_1586_),
    .X(_0248_));
 sky130_fd_sc_hd__and3_1 _3350_ (.A(net112),
    .B(net617),
    .C(_1582_),
    .X(_1587_));
 sky130_fd_sc_hd__a21o_1 _3351_ (.A1(_1120_),
    .A2(_1581_),
    .B1(_1587_),
    .X(_0249_));
 sky130_fd_sc_hd__and3_1 _3352_ (.A(net112),
    .B(net547),
    .C(_1582_),
    .X(_1588_));
 sky130_fd_sc_hd__a21o_1 _3353_ (.A1(_1123_),
    .A2(_1581_),
    .B1(_1588_),
    .X(_0250_));
 sky130_fd_sc_hd__and3_1 _3354_ (.A(net111),
    .B(net549),
    .C(_1582_),
    .X(_1589_));
 sky130_fd_sc_hd__a21o_1 _3355_ (.A1(_1125_),
    .A2(_1581_),
    .B1(_1589_),
    .X(_0251_));
 sky130_fd_sc_hd__and3_1 _3356_ (.A(net110),
    .B(net503),
    .C(_1582_),
    .X(_1590_));
 sky130_fd_sc_hd__a21o_1 _3357_ (.A1(_1128_),
    .A2(_1581_),
    .B1(_1590_),
    .X(_0252_));
 sky130_fd_sc_hd__and3_2 _3358_ (.A(_1107_),
    .B(_1219_),
    .C(_1570_),
    .X(_1591_));
 sky130_fd_sc_hd__or3b_4 _3359_ (.A(_1106_),
    .B(_1220_),
    .C_N(_1570_),
    .X(_1592_));
 sky130_fd_sc_hd__and3_1 _3360_ (.A(net110),
    .B(net541),
    .C(_1592_),
    .X(_1593_));
 sky130_fd_sc_hd__a21o_1 _3361_ (.A1(_1112_),
    .A2(_1591_),
    .B1(_1593_),
    .X(_0253_));
 sky130_fd_sc_hd__and3_1 _3362_ (.A(net111),
    .B(net540),
    .C(_1592_),
    .X(_1594_));
 sky130_fd_sc_hd__a21o_1 _3363_ (.A1(_1114_),
    .A2(_1591_),
    .B1(_1594_),
    .X(_0254_));
 sky130_fd_sc_hd__and3_1 _3364_ (.A(net110),
    .B(net530),
    .C(_1592_),
    .X(_1595_));
 sky130_fd_sc_hd__a21o_1 _3365_ (.A1(_1116_),
    .A2(_1591_),
    .B1(_1595_),
    .X(_0255_));
 sky130_fd_sc_hd__and3_1 _3366_ (.A(net111),
    .B(net572),
    .C(_1592_),
    .X(_1596_));
 sky130_fd_sc_hd__a21o_1 _3367_ (.A1(_1118_),
    .A2(_1591_),
    .B1(_1596_),
    .X(_0256_));
 sky130_fd_sc_hd__and3_1 _3368_ (.A(net111),
    .B(net592),
    .C(_1592_),
    .X(_1597_));
 sky130_fd_sc_hd__a21o_1 _3369_ (.A1(_1120_),
    .A2(_1591_),
    .B1(_1597_),
    .X(_0257_));
 sky130_fd_sc_hd__and3_1 _3370_ (.A(net111),
    .B(net565),
    .C(_1592_),
    .X(_1598_));
 sky130_fd_sc_hd__a21o_1 _3371_ (.A1(_1123_),
    .A2(_1591_),
    .B1(_1598_),
    .X(_0258_));
 sky130_fd_sc_hd__and3_1 _3372_ (.A(net111),
    .B(net526),
    .C(_1592_),
    .X(_1599_));
 sky130_fd_sc_hd__a21o_1 _3373_ (.A1(_1125_),
    .A2(_1591_),
    .B1(_1599_),
    .X(_0259_));
 sky130_fd_sc_hd__and3_1 _3374_ (.A(net110),
    .B(net499),
    .C(_1592_),
    .X(_1600_));
 sky130_fd_sc_hd__a21o_1 _3375_ (.A1(_1128_),
    .A2(_1591_),
    .B1(_1600_),
    .X(_0260_));
 sky130_fd_sc_hd__or3_4 _3376_ (.A(\cmdr[1] ),
    .B(\cmdr[0] ),
    .C(_1064_),
    .X(_1601_));
 sky130_fd_sc_hd__mux2_1 _3377_ (.A0(net81),
    .A1(net360),
    .S(_1601_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _3378_ (.A0(net80),
    .A1(net342),
    .S(_1601_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _3379_ (.A0(net79),
    .A1(net284),
    .S(_1601_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _3380_ (.A0(net78),
    .A1(net348),
    .S(_1601_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _3381_ (.A0(net77),
    .A1(net364),
    .S(_1601_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _3382_ (.A0(net76),
    .A1(net278),
    .S(_1601_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _3383_ (.A0(net75),
    .A1(net204),
    .S(_1601_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _3384_ (.A0(net74),
    .A1(net220),
    .S(_1601_),
    .X(_0268_));
 sky130_fd_sc_hd__nand2_1 _3385_ (.A(\cmdr[1] ),
    .B(\cmdr[0] ),
    .Y(_1602_));
 sky130_fd_sc_hd__or2_1 _3386_ (.A(_1062_),
    .B(_1602_),
    .X(_1603_));
 sky130_fd_sc_hd__nand2b_2 _3387_ (.A_N(\cmdr[2] ),
    .B(\cmdr[3] ),
    .Y(_1604_));
 sky130_fd_sc_hd__or2_4 _3388_ (.A(_1603_),
    .B(_1604_),
    .X(_1605_));
 sky130_fd_sc_hd__mux2_1 _3389_ (.A0(net81),
    .A1(net196),
    .S(_1605_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _3390_ (.A0(net80),
    .A1(net290),
    .S(_1605_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _3391_ (.A0(net79),
    .A1(net132),
    .S(_1605_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _3392_ (.A0(net78),
    .A1(net218),
    .S(_1605_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _3393_ (.A0(net77),
    .A1(net222),
    .S(_1605_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _3394_ (.A0(net76),
    .A1(net232),
    .S(_1605_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _3395_ (.A0(net75),
    .A1(net136),
    .S(_1605_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _3396_ (.A0(net74),
    .A1(net252),
    .S(_1605_),
    .X(_0276_));
 sky130_fd_sc_hd__or3b_2 _3397_ (.A(\cmdr[0] ),
    .B(_1062_),
    .C_N(\cmdr[1] ),
    .X(_1606_));
 sky130_fd_sc_hd__or2_4 _3398_ (.A(_1604_),
    .B(_1606_),
    .X(_1607_));
 sky130_fd_sc_hd__mux2_1 _3399_ (.A0(net81),
    .A1(net306),
    .S(_1607_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _3400_ (.A0(net80),
    .A1(net268),
    .S(_1607_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _3401_ (.A0(net79),
    .A1(net172),
    .S(_1607_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _3402_ (.A0(net78),
    .A1(net312),
    .S(_1607_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _3403_ (.A0(net77),
    .A1(net350),
    .S(_1607_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _3404_ (.A0(net76),
    .A1(net318),
    .S(_1607_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _3405_ (.A0(net75),
    .A1(net264),
    .S(_1607_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _3406_ (.A0(net74),
    .A1(net294),
    .S(_1607_),
    .X(_0284_));
 sky130_fd_sc_hd__or3_2 _3407_ (.A(\cmdr[1] ),
    .B(\cmdr[0] ),
    .C(_1062_),
    .X(_1608_));
 sky130_fd_sc_hd__or3_4 _3408_ (.A(\cmdr[3] ),
    .B(\cmdr[2] ),
    .C(_1608_),
    .X(_1609_));
 sky130_fd_sc_hd__mux2_1 _3409_ (.A0(net81),
    .A1(net286),
    .S(_1609_),
    .X(_0285_));
 sky130_fd_sc_hd__mux2_1 _3410_ (.A0(net80),
    .A1(net224),
    .S(_1609_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _3411_ (.A0(net79),
    .A1(net388),
    .S(_1609_),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _3412_ (.A0(net78),
    .A1(net186),
    .S(_1609_),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _3413_ (.A0(net77),
    .A1(net358),
    .S(_1609_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _3414_ (.A0(net76),
    .A1(net274),
    .S(_1609_),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _3415_ (.A0(net75),
    .A1(net344),
    .S(_1609_),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _3416_ (.A0(net74),
    .A1(net332),
    .S(_1609_),
    .X(_0292_));
 sky130_fd_sc_hd__or2_4 _3417_ (.A(_1604_),
    .B(_1608_),
    .X(_1610_));
 sky130_fd_sc_hd__mux2_1 _3418_ (.A0(net81),
    .A1(net226),
    .S(_1610_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _3419_ (.A0(net80),
    .A1(net280),
    .S(_1610_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _3420_ (.A0(net79),
    .A1(net212),
    .S(_1610_),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _3421_ (.A0(net78),
    .A1(net162),
    .S(_1610_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _3422_ (.A0(net77),
    .A1(net262),
    .S(_1610_),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _3423_ (.A0(net76),
    .A1(net206),
    .S(_1610_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _3424_ (.A0(net75),
    .A1(net244),
    .S(_1610_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _3425_ (.A0(net74),
    .A1(net216),
    .S(_1610_),
    .X(_0300_));
 sky130_fd_sc_hd__nand2b_2 _3426_ (.A_N(\cmdr[3] ),
    .B(\cmdr[2] ),
    .Y(_1611_));
 sky130_fd_sc_hd__or2_4 _3427_ (.A(_1603_),
    .B(_1611_),
    .X(_1612_));
 sky130_fd_sc_hd__mux2_1 _3428_ (.A0(net50),
    .A1(net170),
    .S(_1612_),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _3429_ (.A0(net80),
    .A1(net228),
    .S(_1612_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _3430_ (.A0(net79),
    .A1(net200),
    .S(_1612_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _3431_ (.A0(net78),
    .A1(net182),
    .S(_1612_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _3432_ (.A0(net77),
    .A1(net174),
    .S(_1612_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _3433_ (.A0(net76),
    .A1(net336),
    .S(_1612_),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _3434_ (.A0(net75),
    .A1(net188),
    .S(_1612_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _3435_ (.A0(net74),
    .A1(net202),
    .S(_1612_),
    .X(_0308_));
 sky130_fd_sc_hd__or2_4 _3436_ (.A(_1606_),
    .B(_1611_),
    .X(_1613_));
 sky130_fd_sc_hd__mux2_1 _3437_ (.A0(net50),
    .A1(net352),
    .S(_1613_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _3438_ (.A0(net80),
    .A1(net242),
    .S(_1613_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _3439_ (.A0(net79),
    .A1(net166),
    .S(_1613_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _3440_ (.A0(net78),
    .A1(net234),
    .S(_1613_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _3441_ (.A0(net77),
    .A1(net326),
    .S(_1613_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _3442_ (.A0(net76),
    .A1(net236),
    .S(_1613_),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _3443_ (.A0(net56),
    .A1(net246),
    .S(_1613_),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_1 _3444_ (.A0(net74),
    .A1(net198),
    .S(_1613_),
    .X(_0316_));
 sky130_fd_sc_hd__or2_4 _3445_ (.A(_1608_),
    .B(_1611_),
    .X(_1614_));
 sky130_fd_sc_hd__mux2_1 _3446_ (.A0(net50),
    .A1(net316),
    .S(_1614_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _3447_ (.A0(net80),
    .A1(net154),
    .S(_1614_),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _3448_ (.A0(net79),
    .A1(net130),
    .S(_1614_),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _3449_ (.A0(net78),
    .A1(net164),
    .S(_1614_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _3450_ (.A0(net77),
    .A1(net230),
    .S(_1614_),
    .X(_0321_));
 sky130_fd_sc_hd__mux2_1 _3451_ (.A0(net76),
    .A1(net324),
    .S(_1614_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _3452_ (.A0(net56),
    .A1(net126),
    .S(_1614_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _3453_ (.A0(net74),
    .A1(net190),
    .S(_1614_),
    .X(_0324_));
 sky130_fd_sc_hd__or3b_4 _3454_ (.A(_1062_),
    .B(\cmdr[1] ),
    .C_N(\cmdr[0] ),
    .X(_1615_));
 sky130_fd_sc_hd__nor2_4 _3455_ (.A(_1611_),
    .B(_1615_),
    .Y(_1616_));
 sky130_fd_sc_hd__mux2_1 _3456_ (.A0(net479),
    .A1(net81),
    .S(_1616_),
    .X(_1617_));
 sky130_fd_sc_hd__or2_1 _3457_ (.A(_1771_),
    .B(net480),
    .X(_0325_));
 sky130_fd_sc_hd__nand2_1 _3458_ (.A(net400),
    .B(_1616_),
    .Y(_1618_));
 sky130_fd_sc_hd__o211a_1 _3459_ (.A1(net849),
    .A2(_1616_),
    .B1(net401),
    .C1(net101),
    .X(_0326_));
 sky130_fd_sc_hd__nand2_1 _3460_ (.A(net429),
    .B(_1616_),
    .Y(_1619_));
 sky130_fd_sc_hd__o211a_1 _3461_ (.A1(net394),
    .A2(_1616_),
    .B1(_1619_),
    .C1(net101),
    .X(_0327_));
 sky130_fd_sc_hd__nand2_1 _3462_ (.A(\S8x305.iv_latch[4] ),
    .B(_1616_),
    .Y(_1620_));
 sky130_fd_sc_hd__o211a_1 _3463_ (.A1(net411),
    .A2(_1616_),
    .B1(_1620_),
    .C1(net101),
    .X(_0328_));
 sky130_fd_sc_hd__nand2_1 _3464_ (.A(\S8x305.iv_latch[3] ),
    .B(_1616_),
    .Y(_1621_));
 sky130_fd_sc_hd__o211a_1 _3465_ (.A1(net396),
    .A2(_1616_),
    .B1(_1621_),
    .C1(net101),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _3466_ (.A0(net468),
    .A1(net76),
    .S(_1616_),
    .X(_1622_));
 sky130_fd_sc_hd__or2_1 _3467_ (.A(_1771_),
    .B(net469),
    .X(_0330_));
 sky130_fd_sc_hd__nand2_1 _3468_ (.A(net852),
    .B(_1616_),
    .Y(_1623_));
 sky130_fd_sc_hd__o211a_1 _3469_ (.A1(net398),
    .A2(_1616_),
    .B1(_1623_),
    .C1(net101),
    .X(_0331_));
 sky130_fd_sc_hd__nand2_1 _3470_ (.A(\S8x305.iv_latch[0] ),
    .B(_1616_),
    .Y(_1624_));
 sky130_fd_sc_hd__o211a_1 _3471_ (.A1(net403),
    .A2(_1616_),
    .B1(_1624_),
    .C1(net101),
    .X(_0332_));
 sky130_fd_sc_hd__nand2_1 _3472_ (.A(_1752_),
    .B(net57),
    .Y(_1625_));
 sky130_fd_sc_hd__o211a_1 _3473_ (.A1(net702),
    .A2(net57),
    .B1(_1625_),
    .C1(net96),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _3474_ (.A0(net786),
    .A1(net844),
    .S(net57),
    .X(_1626_));
 sky130_fd_sc_hd__and2_1 _3475_ (.A(net96),
    .B(_1626_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _3476_ (.A0(net455),
    .A1(net692),
    .S(net58),
    .X(_1627_));
 sky130_fd_sc_hd__and2_1 _3477_ (.A(net95),
    .B(_1627_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _3478_ (.A0(net543),
    .A1(net758),
    .S(net57),
    .X(_1628_));
 sky130_fd_sc_hd__and2_1 _3479_ (.A(net95),
    .B(_1628_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _3480_ (.A0(net483),
    .A1(net761),
    .S(net57),
    .X(_1629_));
 sky130_fd_sc_hd__and2_1 _3481_ (.A(net95),
    .B(_1629_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _3482_ (.A0(net639),
    .A1(net766),
    .S(net57),
    .X(_1630_));
 sky130_fd_sc_hd__and2_1 _3483_ (.A(net96),
    .B(_1630_),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _3484_ (.A0(net753),
    .A1(net790),
    .S(net58),
    .X(_1631_));
 sky130_fd_sc_hd__and2_1 _3485_ (.A(net95),
    .B(_1631_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _3486_ (.A0(net672),
    .A1(net736),
    .S(net57),
    .X(_1632_));
 sky130_fd_sc_hd__and2_1 _3487_ (.A(net96),
    .B(_1632_),
    .X(_0340_));
 sky130_fd_sc_hd__nand2_1 _3488_ (.A(_1751_),
    .B(net57),
    .Y(_1633_));
 sky130_fd_sc_hd__o211a_1 _3489_ (.A1(net370),
    .A2(net58),
    .B1(_1633_),
    .C1(net96),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _3490_ (.A0(net494),
    .A1(net767),
    .S(net57),
    .X(_1634_));
 sky130_fd_sc_hd__and2_1 _3491_ (.A(net95),
    .B(_1634_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _3492_ (.A0(net453),
    .A1(net718),
    .S(net58),
    .X(_1635_));
 sky130_fd_sc_hd__and2_1 _3493_ (.A(net95),
    .B(_1635_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _3494_ (.A0(net815),
    .A1(\ROM_addr_buff[12] ),
    .S(net58),
    .X(_1636_));
 sky130_fd_sc_hd__and2_1 _3495_ (.A(net95),
    .B(net816),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _3496_ (.A0(net773),
    .A1(net738),
    .S(net57),
    .X(_1637_));
 sky130_fd_sc_hd__and2_1 _3497_ (.A(net95),
    .B(_1637_),
    .X(_0345_));
 sky130_fd_sc_hd__xnor2_1 _3498_ (.A(_1807_),
    .B(_0756_),
    .Y(_1638_));
 sky130_fd_sc_hd__nor2_1 _3499_ (.A(net59),
    .B(_1638_),
    .Y(_1639_));
 sky130_fd_sc_hd__a21o_1 _3500_ (.A1(net740),
    .A2(net59),
    .B1(net489),
    .X(_1640_));
 sky130_fd_sc_hd__o221a_1 _3501_ (.A1(net702),
    .A2(net600),
    .B1(_1639_),
    .B2(_1640_),
    .C1(net96),
    .X(_0346_));
 sky130_fd_sc_hd__xor2_2 _3502_ (.A(_1804_),
    .B(_0506_),
    .X(_1641_));
 sky130_fd_sc_hd__a21oi_1 _3503_ (.A1(_1807_),
    .A2(_0525_),
    .B1(_1641_),
    .Y(_1642_));
 sky130_fd_sc_hd__a31o_1 _3504_ (.A1(_1807_),
    .A2(_0525_),
    .A3(_1641_),
    .B1(net66),
    .X(_1643_));
 sky130_fd_sc_hd__or2_1 _3505_ (.A(_1642_),
    .B(_1643_),
    .X(_1644_));
 sky130_fd_sc_hd__xor2_2 _3506_ (.A(_1804_),
    .B(_0748_),
    .X(_1645_));
 sky130_fd_sc_hd__and2_1 _3507_ (.A(_1807_),
    .B(_0754_),
    .X(_1646_));
 sky130_fd_sc_hd__o21ai_1 _3508_ (.A1(_1645_),
    .A2(_1646_),
    .B1(net66),
    .Y(_1647_));
 sky130_fd_sc_hd__a21o_1 _3509_ (.A1(_1645_),
    .A2(_1646_),
    .B1(_1647_),
    .X(_1648_));
 sky130_fd_sc_hd__a21oi_1 _3510_ (.A1(_1644_),
    .A2(_1648_),
    .B1(net59),
    .Y(_1649_));
 sky130_fd_sc_hd__a21o_1 _3511_ (.A1(\S8x305.PC[1] ),
    .A2(net59),
    .B1(net489),
    .X(_1650_));
 sky130_fd_sc_hd__o221a_1 _3512_ (.A1(net786),
    .A2(net600),
    .B1(_1649_),
    .B2(_1650_),
    .C1(net96),
    .X(_0347_));
 sky130_fd_sc_hd__nor2_1 _3513_ (.A(_1826_),
    .B(_0731_),
    .Y(_1651_));
 sky130_fd_sc_hd__nand2_1 _3514_ (.A(_1826_),
    .B(_0731_),
    .Y(_1652_));
 sky130_fd_sc_hd__nand2b_1 _3515_ (.A_N(_1651_),
    .B(_1652_),
    .Y(_1653_));
 sky130_fd_sc_hd__a22oi_2 _3516_ (.A1(_1804_),
    .A2(_0748_),
    .B1(_1645_),
    .B2(_1646_),
    .Y(_1654_));
 sky130_fd_sc_hd__xnor2_1 _3517_ (.A(_1653_),
    .B(_1654_),
    .Y(_1655_));
 sky130_fd_sc_hd__xnor2_1 _3518_ (.A(_1826_),
    .B(_0561_),
    .Y(_1656_));
 sky130_fd_sc_hd__a32oi_2 _3519_ (.A1(_1807_),
    .A2(_0525_),
    .A3(_1641_),
    .B1(_0506_),
    .B2(_1804_),
    .Y(_1657_));
 sky130_fd_sc_hd__xnor2_1 _3520_ (.A(_1656_),
    .B(_1657_),
    .Y(_1658_));
 sky130_fd_sc_hd__mux2_1 _3521_ (.A0(_1655_),
    .A1(_1658_),
    .S(net61),
    .X(_1659_));
 sky130_fd_sc_hd__nor2_1 _3522_ (.A(net59),
    .B(_1659_),
    .Y(_1660_));
 sky130_fd_sc_hd__a21o_1 _3523_ (.A1(net470),
    .A2(net59),
    .B1(net489),
    .X(_1661_));
 sky130_fd_sc_hd__o221a_1 _3524_ (.A1(net455),
    .A2(net600),
    .B1(_1660_),
    .B2(_1661_),
    .C1(net96),
    .X(_0348_));
 sky130_fd_sc_hd__xnor2_1 _3525_ (.A(_0436_),
    .B(_0543_),
    .Y(_1662_));
 sky130_fd_sc_hd__o21ba_1 _3526_ (.A1(_1826_),
    .A2(_0561_),
    .B1_N(_1657_),
    .X(_1663_));
 sky130_fd_sc_hd__a21oi_1 _3527_ (.A1(_1826_),
    .A2(_0561_),
    .B1(_1663_),
    .Y(_1664_));
 sky130_fd_sc_hd__xnor2_1 _3528_ (.A(_1662_),
    .B(_1664_),
    .Y(_1665_));
 sky130_fd_sc_hd__xnor2_1 _3529_ (.A(_0436_),
    .B(_0721_),
    .Y(_1666_));
 sky130_fd_sc_hd__o21a_1 _3530_ (.A1(_1651_),
    .A2(_1654_),
    .B1(_1652_),
    .X(_1667_));
 sky130_fd_sc_hd__xnor2_1 _3531_ (.A(_1666_),
    .B(_1667_),
    .Y(_1668_));
 sky130_fd_sc_hd__mux2_1 _3532_ (.A0(_1665_),
    .A1(_1668_),
    .S(net66),
    .X(_1669_));
 sky130_fd_sc_hd__nor2_1 _3533_ (.A(net59),
    .B(_1669_),
    .Y(_1670_));
 sky130_fd_sc_hd__a21o_1 _3534_ (.A1(net750),
    .A2(net59),
    .B1(net489),
    .X(_1671_));
 sky130_fd_sc_hd__o221a_1 _3535_ (.A1(net543),
    .A2(net600),
    .B1(_1670_),
    .B2(_1671_),
    .C1(net103),
    .X(_0349_));
 sky130_fd_sc_hd__o21ba_1 _3536_ (.A1(_0436_),
    .A2(_0721_),
    .B1_N(_1667_),
    .X(_1672_));
 sky130_fd_sc_hd__a21oi_1 _3537_ (.A1(_0436_),
    .A2(_0721_),
    .B1(_1672_),
    .Y(_1673_));
 sky130_fd_sc_hd__xnor2_1 _3538_ (.A(_1820_),
    .B(_1673_),
    .Y(_1674_));
 sky130_fd_sc_hd__xnor2_1 _3539_ (.A(_0709_),
    .B(_1674_),
    .Y(_1675_));
 sky130_fd_sc_hd__xnor2_1 _3540_ (.A(_1820_),
    .B(_0624_),
    .Y(_1676_));
 sky130_fd_sc_hd__o21ba_1 _3541_ (.A1(_0436_),
    .A2(_0543_),
    .B1_N(_1664_),
    .X(_1677_));
 sky130_fd_sc_hd__a21oi_1 _3542_ (.A1(_0436_),
    .A2(_0543_),
    .B1(_1677_),
    .Y(_1678_));
 sky130_fd_sc_hd__xnor2_1 _3543_ (.A(_1676_),
    .B(_1678_),
    .Y(_1679_));
 sky130_fd_sc_hd__mux2_1 _3544_ (.A0(_1675_),
    .A1(_1679_),
    .S(net61),
    .X(_1680_));
 sky130_fd_sc_hd__nor2_1 _3545_ (.A(net59),
    .B(_1680_),
    .Y(_1681_));
 sky130_fd_sc_hd__a21o_1 _3546_ (.A1(net742),
    .A2(net59),
    .B1(net489),
    .X(_1682_));
 sky130_fd_sc_hd__o221a_1 _3547_ (.A1(net483),
    .A2(net600),
    .B1(_1681_),
    .B2(_1682_),
    .C1(net103),
    .X(_0350_));
 sky130_fd_sc_hd__o21ba_1 _3548_ (.A1(_1820_),
    .A2(_0624_),
    .B1_N(_1678_),
    .X(_1683_));
 sky130_fd_sc_hd__a21oi_1 _3549_ (.A1(_1820_),
    .A2(_0624_),
    .B1(_1683_),
    .Y(_1684_));
 sky130_fd_sc_hd__nor2_1 _3550_ (.A(_0606_),
    .B(_0805_),
    .Y(_1685_));
 sky130_fd_sc_hd__nand2_1 _3551_ (.A(_0606_),
    .B(_0805_),
    .Y(_1686_));
 sky130_fd_sc_hd__and2b_1 _3552_ (.A_N(_1685_),
    .B(_1686_),
    .X(_1687_));
 sky130_fd_sc_hd__xnor2_1 _3553_ (.A(_1684_),
    .B(_1687_),
    .Y(_1688_));
 sky130_fd_sc_hd__nor2_1 _3554_ (.A(net66),
    .B(net59),
    .Y(_1689_));
 sky130_fd_sc_hd__a221o_1 _3555_ (.A1(net729),
    .A2(net59),
    .B1(_1688_),
    .B2(_1689_),
    .C1(net489),
    .X(_1690_));
 sky130_fd_sc_hd__o211a_1 _3556_ (.A1(net639),
    .A2(net600),
    .B1(_1690_),
    .C1(net103),
    .X(_0351_));
 sky130_fd_sc_hd__or2_1 _3557_ (.A(_0642_),
    .B(_0793_),
    .X(_1691_));
 sky130_fd_sc_hd__nand2_1 _3558_ (.A(_0642_),
    .B(_0793_),
    .Y(_1692_));
 sky130_fd_sc_hd__nand2_1 _3559_ (.A(_1691_),
    .B(_1692_),
    .Y(_1693_));
 sky130_fd_sc_hd__o21a_1 _3560_ (.A1(_1684_),
    .A2(_1685_),
    .B1(_1686_),
    .X(_1694_));
 sky130_fd_sc_hd__nand2_1 _3561_ (.A(_1693_),
    .B(_1694_),
    .Y(_1695_));
 sky130_fd_sc_hd__or2_1 _3562_ (.A(_1693_),
    .B(_1694_),
    .X(_1696_));
 sky130_fd_sc_hd__a32o_1 _3563_ (.A1(_1689_),
    .A2(_1695_),
    .A3(_1696_),
    .B1(net59),
    .B2(net800),
    .X(_1697_));
 sky130_fd_sc_hd__or2_1 _3564_ (.A(net753),
    .B(net600),
    .X(_1698_));
 sky130_fd_sc_hd__o211a_1 _3565_ (.A1(net489),
    .A2(_1697_),
    .B1(_1698_),
    .C1(net98),
    .X(_0352_));
 sky130_fd_sc_hd__xnor2_1 _3566_ (.A(_0460_),
    .B(_0588_),
    .Y(_1699_));
 sky130_fd_sc_hd__a21o_1 _3567_ (.A1(_1692_),
    .A2(_1696_),
    .B1(_1699_),
    .X(_1700_));
 sky130_fd_sc_hd__a311oi_1 _3568_ (.A1(_1692_),
    .A2(_1696_),
    .A3(_1699_),
    .B1(_0466_),
    .C1(net66),
    .Y(_1701_));
 sky130_fd_sc_hd__a221o_1 _3569_ (.A1(net472),
    .A2(net59),
    .B1(_1700_),
    .B2(_1701_),
    .C1(net489),
    .X(_1702_));
 sky130_fd_sc_hd__o211a_1 _3570_ (.A1(net672),
    .A2(net600),
    .B1(_1702_),
    .C1(net103),
    .X(_0353_));
 sky130_fd_sc_hd__or2_1 _3571_ (.A(net370),
    .B(_0486_),
    .X(_1703_));
 sky130_fd_sc_hd__o211a_1 _3572_ (.A1(net463),
    .A2(net489),
    .B1(_1703_),
    .C1(net103),
    .X(_0354_));
 sky130_fd_sc_hd__or2_1 _3573_ (.A(\S8x305.A[9] ),
    .B(_0486_),
    .X(_1704_));
 sky130_fd_sc_hd__o211a_1 _3574_ (.A1(net441),
    .A2(_0487_),
    .B1(_1704_),
    .C1(net103),
    .X(_0355_));
 sky130_fd_sc_hd__or2_1 _3575_ (.A(net453),
    .B(_0486_),
    .X(_1705_));
 sky130_fd_sc_hd__o211a_1 _3576_ (.A1(net556),
    .A2(net489),
    .B1(net601),
    .C1(net103),
    .X(_0356_));
 sky130_fd_sc_hd__or2_1 _3577_ (.A(\S8x305.A[11] ),
    .B(_0486_),
    .X(_1706_));
 sky130_fd_sc_hd__o211a_1 _3578_ (.A1(net122),
    .A2(_0487_),
    .B1(_1706_),
    .C1(net96),
    .X(_0357_));
 sky130_fd_sc_hd__or2_1 _3579_ (.A(\S8x305.A[12] ),
    .B(_0486_),
    .X(_1707_));
 sky130_fd_sc_hd__o211a_1 _3580_ (.A1(net445),
    .A2(_0487_),
    .B1(_1707_),
    .C1(net103),
    .X(_0358_));
 sky130_fd_sc_hd__nor2_1 _3581_ (.A(_1808_),
    .B(_1080_),
    .Y(_1708_));
 sky130_fd_sc_hd__o21ai_1 _3582_ (.A1(net740),
    .A2(_1079_),
    .B1(_1075_),
    .Y(_1709_));
 sky130_fd_sc_hd__o221a_1 _3583_ (.A1(net740),
    .A2(_1075_),
    .B1(_1708_),
    .B2(_1709_),
    .C1(net96),
    .X(_0359_));
 sky130_fd_sc_hd__nand2_1 _3584_ (.A(net740),
    .B(_1080_),
    .Y(_1710_));
 sky130_fd_sc_hd__a2bb2o_1 _3585_ (.A1_N(net801),
    .A2_N(_1710_),
    .B1(_1079_),
    .B2(_1804_),
    .X(_1711_));
 sky130_fd_sc_hd__a22o_1 _3586_ (.A1(net801),
    .A2(_1709_),
    .B1(_1711_),
    .B2(_1075_),
    .X(_1712_));
 sky130_fd_sc_hd__and2_1 _3587_ (.A(net96),
    .B(_1712_),
    .X(_0360_));
 sky130_fd_sc_hd__a21oi_1 _3588_ (.A1(\S8x305.PC[1] ),
    .A2(\S8x305.PC[0] ),
    .B1(net470),
    .Y(_1713_));
 sky130_fd_sc_hd__nor3_1 _3589_ (.A(_1079_),
    .B(_1081_),
    .C(_1713_),
    .Y(_1714_));
 sky130_fd_sc_hd__a21o_1 _3590_ (.A1(_1826_),
    .A2(_1079_),
    .B1(_1076_),
    .X(_1715_));
 sky130_fd_sc_hd__o221a_1 _3591_ (.A1(net470),
    .A2(_1075_),
    .B1(_1714_),
    .B2(_1715_),
    .C1(net103),
    .X(_0361_));
 sky130_fd_sc_hd__or2_1 _3592_ (.A(net750),
    .B(_1081_),
    .X(_1716_));
 sky130_fd_sc_hd__and3_1 _3593_ (.A(_1080_),
    .B(_1082_),
    .C(_1716_),
    .X(_1717_));
 sky130_fd_sc_hd__a21o_1 _3594_ (.A1(_0436_),
    .A2(_1079_),
    .B1(_1076_),
    .X(_1718_));
 sky130_fd_sc_hd__o221a_1 _3595_ (.A1(net750),
    .A2(_1075_),
    .B1(_1717_),
    .B2(_1718_),
    .C1(net103),
    .X(_0362_));
 sky130_fd_sc_hd__nor2_1 _3596_ (.A(_1819_),
    .B(_1080_),
    .Y(_1719_));
 sky130_fd_sc_hd__a21o_1 _3597_ (.A1(\S8x305.PC[3] ),
    .A2(_1081_),
    .B1(net742),
    .X(_1720_));
 sky130_fd_sc_hd__a31o_1 _3598_ (.A1(_1080_),
    .A2(_1083_),
    .A3(_1720_),
    .B1(_1076_),
    .X(_1721_));
 sky130_fd_sc_hd__o221a_1 _3599_ (.A1(net742),
    .A2(_1075_),
    .B1(_1719_),
    .B2(_1721_),
    .C1(net104),
    .X(_0363_));
 sky130_fd_sc_hd__or2_1 _3600_ (.A(net599),
    .B(net84),
    .X(_1722_));
 sky130_fd_sc_hd__and3_1 _3601_ (.A(net97),
    .B(_1073_),
    .C(_1722_),
    .X(_0364_));
 sky130_fd_sc_hd__nand2_1 _3602_ (.A(net82),
    .B(_1073_),
    .Y(_1723_));
 sky130_fd_sc_hd__a21oi_1 _3603_ (.A1(_1074_),
    .A2(_1723_),
    .B1(_1771_),
    .Y(_0365_));
 sky130_fd_sc_hd__or3_4 _3604_ (.A(\cmdr[3] ),
    .B(\cmdr[2] ),
    .C(_1603_),
    .X(_1724_));
 sky130_fd_sc_hd__mux2_1 _3605_ (.A0(net81),
    .A1(net258),
    .S(_1724_),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_1 _3606_ (.A0(net80),
    .A1(net272),
    .S(_1724_),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _3607_ (.A0(net79),
    .A1(net282),
    .S(_1724_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _3608_ (.A0(net78),
    .A1(net192),
    .S(_1724_),
    .X(_0369_));
 sky130_fd_sc_hd__mux2_1 _3609_ (.A0(net77),
    .A1(net184),
    .S(_1724_),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _3610_ (.A0(net76),
    .A1(net144),
    .S(_1724_),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _3611_ (.A0(net75),
    .A1(net346),
    .S(_1724_),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _3612_ (.A0(net74),
    .A1(net314),
    .S(_1724_),
    .X(_0373_));
 sky130_fd_sc_hd__or3_4 _3613_ (.A(\cmdr[3] ),
    .B(\cmdr[2] ),
    .C(_1606_),
    .X(_1725_));
 sky130_fd_sc_hd__mux2_1 _3614_ (.A0(net81),
    .A1(net384),
    .S(_1725_),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_1 _3615_ (.A0(net80),
    .A1(net366),
    .S(_1725_),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_1 _3616_ (.A0(net52),
    .A1(net356),
    .S(_1725_),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _3617_ (.A0(net78),
    .A1(net304),
    .S(_1725_),
    .X(_0377_));
 sky130_fd_sc_hd__mux2_1 _3618_ (.A0(net77),
    .A1(net380),
    .S(_1725_),
    .X(_0378_));
 sky130_fd_sc_hd__mux2_1 _3619_ (.A0(net55),
    .A1(net270),
    .S(_1725_),
    .X(_0379_));
 sky130_fd_sc_hd__mux2_1 _3620_ (.A0(net75),
    .A1(net354),
    .S(_1725_),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_1 _3621_ (.A0(net74),
    .A1(net266),
    .S(_1725_),
    .X(_0381_));
 sky130_fd_sc_hd__or3_4 _3622_ (.A(\cmdr[3] ),
    .B(\cmdr[2] ),
    .C(_1615_),
    .X(_1726_));
 sky130_fd_sc_hd__mux2_1 _3623_ (.A0(net81),
    .A1(net340),
    .S(_1726_),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _3624_ (.A0(net51),
    .A1(net308),
    .S(_1726_),
    .X(_0383_));
 sky130_fd_sc_hd__mux2_1 _3625_ (.A0(net52),
    .A1(net248),
    .S(_1726_),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _3626_ (.A0(net78),
    .A1(net330),
    .S(_1726_),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _3627_ (.A0(net77),
    .A1(net276),
    .S(_1726_),
    .X(_0386_));
 sky130_fd_sc_hd__mux2_1 _3628_ (.A0(net55),
    .A1(net328),
    .S(_1726_),
    .X(_0387_));
 sky130_fd_sc_hd__mux2_1 _3629_ (.A0(net75),
    .A1(net288),
    .S(_1726_),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _3630_ (.A0(net74),
    .A1(net382),
    .S(_1726_),
    .X(_0389_));
 sky130_fd_sc_hd__or2_4 _3631_ (.A(_1064_),
    .B(_1602_),
    .X(_1727_));
 sky130_fd_sc_hd__mux2_1 _3632_ (.A0(net81),
    .A1(net296),
    .S(_1727_),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _3633_ (.A0(net80),
    .A1(net320),
    .S(_1727_),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_1 _3634_ (.A0(net79),
    .A1(net260),
    .S(_1727_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _3635_ (.A0(net78),
    .A1(net178),
    .S(_1727_),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_1 _3636_ (.A0(net77),
    .A1(net238),
    .S(_1727_),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _3637_ (.A0(net76),
    .A1(net256),
    .S(_1727_),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _3638_ (.A0(net75),
    .A1(net210),
    .S(_1727_),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _3639_ (.A0(net74),
    .A1(net160),
    .S(_1727_),
    .X(_0397_));
 sky130_fd_sc_hd__and3_2 _3640_ (.A(_1107_),
    .B(_1146_),
    .C(_1570_),
    .X(_1728_));
 sky130_fd_sc_hd__or3b_2 _3641_ (.A(_1106_),
    .B(_1147_),
    .C_N(_1570_),
    .X(_1729_));
 sky130_fd_sc_hd__and3_1 _3642_ (.A(net110),
    .B(net789),
    .C(_1729_),
    .X(_1730_));
 sky130_fd_sc_hd__a21o_1 _3643_ (.A1(_1112_),
    .A2(_1728_),
    .B1(_1730_),
    .X(_0398_));
 sky130_fd_sc_hd__and3_1 _3644_ (.A(net111),
    .B(net845),
    .C(_1729_),
    .X(_1731_));
 sky130_fd_sc_hd__a21o_1 _3645_ (.A1(_1114_),
    .A2(_1728_),
    .B1(_1731_),
    .X(_0399_));
 sky130_fd_sc_hd__and3_1 _3646_ (.A(net110),
    .B(net813),
    .C(_1729_),
    .X(_1732_));
 sky130_fd_sc_hd__a21o_1 _3647_ (.A1(_1116_),
    .A2(_1728_),
    .B1(_1732_),
    .X(_0400_));
 sky130_fd_sc_hd__and3_1 _3648_ (.A(net111),
    .B(net814),
    .C(_1729_),
    .X(_1733_));
 sky130_fd_sc_hd__a21o_1 _3649_ (.A1(_1118_),
    .A2(_1728_),
    .B1(_1733_),
    .X(_0401_));
 sky130_fd_sc_hd__and3_1 _3650_ (.A(net111),
    .B(net805),
    .C(_1729_),
    .X(_1734_));
 sky130_fd_sc_hd__a21o_1 _3651_ (.A1(_1120_),
    .A2(_1728_),
    .B1(_1734_),
    .X(_0402_));
 sky130_fd_sc_hd__and3_1 _3652_ (.A(net111),
    .B(net812),
    .C(_1729_),
    .X(_1735_));
 sky130_fd_sc_hd__a21o_1 _3653_ (.A1(_1123_),
    .A2(_1728_),
    .B1(_1735_),
    .X(_0403_));
 sky130_fd_sc_hd__and3_1 _3654_ (.A(net111),
    .B(net788),
    .C(_1729_),
    .X(_1736_));
 sky130_fd_sc_hd__a21o_1 _3655_ (.A1(_1125_),
    .A2(_1728_),
    .B1(_1736_),
    .X(_0404_));
 sky130_fd_sc_hd__and3_1 _3656_ (.A(net110),
    .B(net771),
    .C(_1729_),
    .X(_1737_));
 sky130_fd_sc_hd__a21o_1 _3657_ (.A1(_1128_),
    .A2(_1728_),
    .B1(_1737_),
    .X(_0405_));
 sky130_fd_sc_hd__nand2_8 _3658_ (.A(net599),
    .B(net98),
    .Y(_1738_));
 sky130_fd_sc_hd__mux2_1 _3659_ (.A0(_1807_),
    .A1(net437),
    .S(_1738_),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_1 _3660_ (.A0(_1804_),
    .A1(net390),
    .S(_1738_),
    .X(_0407_));
 sky130_fd_sc_hd__mux2_1 _3661_ (.A0(_1826_),
    .A1(net378),
    .S(_1738_),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_1 _3662_ (.A0(_0436_),
    .A1(net433),
    .S(_1738_),
    .X(_0409_));
 sky130_fd_sc_hd__mux2_1 _3663_ (.A0(_1820_),
    .A1(net757),
    .S(_1738_),
    .X(_0410_));
 sky130_fd_sc_hd__mux2_1 _3664_ (.A0(_0474_),
    .A1(net386),
    .S(_1738_),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _3665_ (.A0(_0469_),
    .A1(net451),
    .S(_1738_),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_1 _3666_ (.A0(_0459_),
    .A1(net710),
    .S(_1738_),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _3667_ (.A0(net71),
    .A1(net407),
    .S(_1738_),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _3668_ (.A0(net73),
    .A1(net686),
    .S(_1738_),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_1 _3669_ (.A0(net60),
    .A1(net713),
    .S(_1738_),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_1 _3670_ (.A0(_0434_),
    .A1(net684),
    .S(_1738_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _3671_ (.A0(net66),
    .A1(net449),
    .S(_1738_),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _3672_ (.A0(_1788_),
    .A1(net459),
    .S(_1738_),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_1 _3673_ (.A0(_1796_),
    .A1(net760),
    .S(_1738_),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _3674_ (.A0(_1792_),
    .A1(net158),
    .S(_1738_),
    .X(_0421_));
 sky130_fd_sc_hd__or2_4 _3675_ (.A(_1604_),
    .B(_1615_),
    .X(_1739_));
 sky130_fd_sc_hd__mux2_1 _3676_ (.A0(net81),
    .A1(net176),
    .S(_1739_),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_1 _3677_ (.A0(net51),
    .A1(net180),
    .S(_1739_),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _3678_ (.A0(net52),
    .A1(net148),
    .S(_1739_),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_1 _3679_ (.A0(net53),
    .A1(net334),
    .S(_1739_),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_1 _3680_ (.A0(net54),
    .A1(net372),
    .S(_1739_),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_1 _3681_ (.A0(net55),
    .A1(net292),
    .S(_1739_),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _3682_ (.A0(net75),
    .A1(net142),
    .S(_1739_),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _3683_ (.A0(net30),
    .A1(net250),
    .S(_1739_),
    .X(_0429_));
 sky130_fd_sc_hd__o211a_1 _3684_ (.A1(net680),
    .A2(_1130_),
    .B1(_1131_),
    .C1(net100),
    .X(_0187_));
 sky130_fd_sc_hd__o211a_1 _3685_ (.A1(net641),
    .A2(_1130_),
    .B1(_1132_),
    .C1(net100),
    .X(_0188_));
 sky130_fd_sc_hd__o211a_1 _3686_ (.A1(net809),
    .A2(_1130_),
    .B1(_1133_),
    .C1(net100),
    .X(_0189_));
 sky130_fd_sc_hd__o211a_1 _3687_ (.A1(net730),
    .A2(_1130_),
    .B1(_1134_),
    .C1(net100),
    .X(_0190_));
 sky130_fd_sc_hd__dfxtp_2 _3688_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0004_),
    .Q(\S8x305.iv_latch[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3689_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0005_),
    .Q(\S8x305.iv_latch[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3690_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0006_),
    .Q(\S8x305.iv_latch[5] ));
 sky130_fd_sc_hd__dfxtp_4 _3691_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0007_),
    .Q(\S8x305.iv_latch[4] ));
 sky130_fd_sc_hd__dfxtp_4 _3692_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0008_),
    .Q(\S8x305.iv_latch[3] ));
 sky130_fd_sc_hd__dfxtp_2 _3693_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0009_),
    .Q(\S8x305.iv_latch[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3694_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0010_),
    .Q(\S8x305.iv_latch[1] ));
 sky130_fd_sc_hd__dfxtp_2 _3695_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net785),
    .Q(\S8x305.iv_latch[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3696_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net375),
    .Q(\memory[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3697_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net339),
    .Q(\memory[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3698_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net311),
    .Q(\memory[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3699_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net377),
    .Q(\memory[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3700_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net363),
    .Q(\memory[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3701_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net301),
    .Q(\memory[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3702_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net303),
    .Q(\memory[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3703_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net323),
    .Q(\memory[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3704_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0020_),
    .Q(\S8x305.PC[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3705_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0021_),
    .Q(\S8x305.PC[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3706_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0022_),
    .Q(\S8x305.PC[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3707_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0023_),
    .Q(\S8x305.PC[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3708_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0024_),
    .Q(\S8x305.PC[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3709_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net623),
    .Q(\S8x305.regs[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3710_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0026_),
    .Q(\S8x305.regs[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3711_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0027_),
    .Q(\S8x305.regs[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3712_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0028_),
    .Q(\S8x305.regs[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3713_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net629),
    .Q(\S8x305.regs[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3714_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0030_),
    .Q(\S8x305.regs[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3715_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0031_),
    .Q(\S8x305.regs[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3716_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0032_),
    .Q(\S8x305.regs[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3717_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net681),
    .Q(_0000_));
 sky130_fd_sc_hd__dfxtp_1 _3718_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net667),
    .Q(_0001_));
 sky130_fd_sc_hd__dfxtp_1 _3719_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0035_),
    .Q(_0002_));
 sky130_fd_sc_hd__dfxtp_4 _3720_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net735),
    .Q(_0003_));
 sky130_fd_sc_hd__dfxtp_1 _3721_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net578),
    .Q(\S8x305.regs[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3722_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0038_),
    .Q(\S8x305.regs[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3723_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0039_),
    .Q(\S8x305.regs[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3724_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0040_),
    .Q(\S8x305.regs[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3725_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0041_),
    .Q(\S8x305.regs[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3726_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0042_),
    .Q(\S8x305.regs[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3727_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0043_),
    .Q(\S8x305.regs[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3728_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0044_),
    .Q(\S8x305.regs[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3729_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net169),
    .Q(\S8x305.regs[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3730_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net147),
    .Q(\S8x305.regs[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3731_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net153),
    .Q(\S8x305.regs[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3732_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net141),
    .Q(\S8x305.regs[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3733_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net209),
    .Q(\S8x305.regs[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3734_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net129),
    .Q(\S8x305.regs[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3735_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net157),
    .Q(\S8x305.regs[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3736_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0052_),
    .Q(\S8x305.PC[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3737_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0053_),
    .Q(\S8x305.PC[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3738_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0054_),
    .Q(\S8x305.PC[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3739_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0055_),
    .Q(\S8x305.regs[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3740_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net574),
    .Q(\S8x305.regs[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3741_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net529),
    .Q(\S8x305.regs[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3742_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0058_),
    .Q(\S8x305.regs[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3743_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0059_),
    .Q(\S8x305.regs[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3744_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net631),
    .Q(\S8x305.regs[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3745_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0061_),
    .Q(\S8x305.regs[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3746_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0062_),
    .Q(\S8x305.regs[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3747_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net508),
    .Q(\S8x305.regs[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3748_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net647),
    .Q(\S8x305.regs[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3749_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net569),
    .Q(\S8x305.regs[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3750_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0066_),
    .Q(\S8x305.regs[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3751_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0067_),
    .Q(\S8x305.regs[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3752_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0068_),
    .Q(\S8x305.regs[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3753_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0069_),
    .Q(\S8x305.regs[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3754_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0070_),
    .Q(\S8x305.regs[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3755_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net603),
    .Q(\S8x305.regs[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3756_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net514),
    .Q(\S8x305.regs[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3757_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net576),
    .Q(\S8x305.regs[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3758_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0074_),
    .Q(\S8x305.regs[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3759_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0075_),
    .Q(\S8x305.regs[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3760_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0076_),
    .Q(\S8x305.regs[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3761_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0077_),
    .Q(\S8x305.regs[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3762_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0078_),
    .Q(\S8x305.regs[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3763_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net546),
    .Q(\S8x305.regs[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3764_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net654),
    .Q(\S8x305.regs[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3765_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net560),
    .Q(\S8x305.regs[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3766_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0082_),
    .Q(\S8x305.regs[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3767_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0083_),
    .Q(\S8x305.regs[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3768_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net607),
    .Q(\S8x305.regs[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3769_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0085_),
    .Q(\S8x305.regs[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3770_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0086_),
    .Q(\S8x305.regs[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3771_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net649),
    .Q(\S8x305.regs[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3772_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net554),
    .Q(\S8x305.regs[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3773_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net512),
    .Q(\S8x305.regs[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3774_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0090_),
    .Q(\S8x305.regs[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3775_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0091_),
    .Q(\S8x305.regs[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3776_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net532),
    .Q(\S8x305.regs[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3777_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0093_),
    .Q(\S8x305.regs[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3778_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0094_),
    .Q(\S8x305.regs[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3779_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net612),
    .Q(\S8x305.regs[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3780_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net707),
    .Q(\S8x305.regs[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3781_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0097_),
    .Q(\S8x305.regs[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3782_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0098_),
    .Q(\S8x305.regs[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3783_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0099_),
    .Q(\S8x305.regs[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3784_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net626),
    .Q(\S8x305.regs[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3785_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0101_),
    .Q(\S8x305.regs[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3786_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0102_),
    .Q(\S8x305.regs[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3787_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0103_),
    .Q(\S8x305.regs[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3788_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net656),
    .Q(\S8x305.regs[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3789_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0105_),
    .Q(\S8x305.regs[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3790_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0106_),
    .Q(\S8x305.regs[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3791_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0107_),
    .Q(\S8x305.regs[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3792_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net605),
    .Q(\S8x305.regs[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3793_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0109_),
    .Q(\S8x305.regs[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3794_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0110_),
    .Q(\S8x305.regs[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3795_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net594),
    .Q(\S8x305.regs[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3796_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net552),
    .Q(\S8x305.regs[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3797_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0113_),
    .Q(\S8x305.regs[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3798_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0114_),
    .Q(\S8x305.regs[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3799_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0115_),
    .Q(\S8x305.regs[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3800_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net580),
    .Q(\S8x305.regs[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3801_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0117_),
    .Q(\S8x305.regs[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3802_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0118_),
    .Q(\S8x305.regs[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3803_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net525),
    .Q(\S8x305.regs[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3804_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net426),
    .Q(\S8x305.I[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3805_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net422),
    .Q(\S8x305.I[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3806_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net406),
    .Q(\S8x305.I[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3807_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net428),
    .Q(\S8x305.I[7] ));
 sky130_fd_sc_hd__dfxtp_2 _3808_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0124_),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_1 _3809_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net634),
    .Q(net43));
 sky130_fd_sc_hd__dfxtp_1 _3810_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net621),
    .Q(net44));
 sky130_fd_sc_hd__dfxtp_1 _3811_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net705),
    .Q(net45));
 sky130_fd_sc_hd__dfxtp_1 _3812_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net658),
    .Q(net46));
 sky130_fd_sc_hd__dfxtp_1 _3813_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net669),
    .Q(net47));
 sky130_fd_sc_hd__dfxtp_2 _3814_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0130_),
    .Q(net48));
 sky130_fd_sc_hd__dfxtp_1 _3815_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0131_),
    .Q(net49));
 sky130_fd_sc_hd__dfxtp_1 _3816_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net765),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_2 _3817_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net728),
    .Q(\ROM_spi_cycle[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3818_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net819),
    .Q(\ROM_spi_cycle[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3819_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net432),
    .Q(\ROM_spi_cycle[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3820_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net695),
    .Q(\ROM_spi_cycle[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3821_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net689),
    .Q(\ROM_spi_cycle[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3822_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net770),
    .Q(\startup_cycle[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3823_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net478),
    .Q(\startup_cycle[1] ));
 sky130_fd_sc_hd__dfxtp_2 _3824_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net808),
    .Q(\startup_cycle[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3825_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net662),
    .Q(\startup_cycle[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3826_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net700),
    .Q(\startup_cycle[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3827_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net723),
    .Q(\startup_cycle[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3828_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net721),
    .Q(\startup_cycle[6] ));
 sky130_fd_sc_hd__dfxtp_2 _3829_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net843),
    .Q(\mem_cycle[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3830_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0146_),
    .Q(\mem_cycle[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3831_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net444),
    .Q(\mem_cycle[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3832_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net832),
    .Q(\mem_cycle[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3833_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0149_),
    .Q(\mem_cycle[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3834_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0150_),
    .Q(\mem_cycle[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3835_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net745),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_1 _3836_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0152_),
    .Q(net42));
 sky130_fd_sc_hd__dfxtp_1 _3837_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0153_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_1 _3838_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net448),
    .Q(ROM_OEB));
 sky130_fd_sc_hd__dfxtp_1 _3839_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net215),
    .Q(ROM_spi_mode));
 sky130_fd_sc_hd__dfxtp_1 _3840_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net393),
    .Q(\ROM_spi_dat_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3841_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net410),
    .Q(\ROM_spi_dat_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3842_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net418),
    .Q(\ROM_spi_dat_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3843_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net414),
    .Q(\ROM_spi_dat_out[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3844_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net420),
    .Q(\ROM_spi_dat_out[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3845_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net416),
    .Q(\ROM_spi_dat_out[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3846_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net502),
    .Q(\ROM_spi_dat_out[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3847_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net424),
    .Q(\ROM_spi_dat_out[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3848_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net125),
    .Q(\last_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3849_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0165_),
    .Q(\last_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3850_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0166_),
    .Q(\last_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3851_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net697),
    .Q(\last_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3852_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net763),
    .Q(\last_addr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3853_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0169_),
    .Q(\last_addr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3854_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0170_),
    .Q(\last_addr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3855_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0171_),
    .Q(\last_addr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3856_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0172_),
    .Q(\last_addr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3857_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0173_),
    .Q(\last_addr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3858_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net683),
    .Q(\last_addr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3859_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net775),
    .Q(\last_addr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3860_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net717),
    .Q(\last_addr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3861_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net739),
    .Q(\last_addr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3862_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(_0178_),
    .Q(spi_clkdiv));
 sky130_fd_sc_hd__dfxtp_1 _3863_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net517),
    .Q(\cmdl[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3864_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net487),
    .Q(\cmdl[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3865_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net462),
    .Q(\cmdl[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3866_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net497),
    .Q(\cmdl[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3867_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net482),
    .Q(\cmdl[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3868_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net458),
    .Q(\cmdl[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3869_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net436),
    .Q(\cmdl[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3870_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net467),
    .Q(\cmdl[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3871_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net691),
    .Q(\cmdr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _3872_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net642),
    .Q(\cmdr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _3873_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net810),
    .Q(\cmdr[2] ));
 sky130_fd_sc_hd__dfxtp_2 _3874_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net731),
    .Q(\cmdr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3875_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net506),
    .Q(\cmdr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3876_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net430),
    .Q(\cmdr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3877_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net440),
    .Q(\cmdr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3878_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net476),
    .Q(\cmdr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3879_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0195_),
    .Q(\last_A[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3880_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0196_),
    .Q(\last_A[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3881_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0197_),
    .Q(\last_A[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3882_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0198_),
    .Q(\last_A[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3883_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0199_),
    .Q(\last_A[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3884_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0200_),
    .Q(\last_A[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3885_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0201_),
    .Q(\last_A[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3886_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0202_),
    .Q(\last_A[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3887_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0203_),
    .Q(\last_A[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3888_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0204_),
    .Q(\last_A[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3889_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0205_),
    .Q(\last_A[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3890_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net195),
    .Q(\memory[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3891_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net369),
    .Q(\memory[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3892_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net299),
    .Q(\memory[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3893_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net135),
    .Q(\memory[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3894_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net139),
    .Q(\memory[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3895_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net151),
    .Q(\memory[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3896_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net241),
    .Q(\memory[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3897_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net255),
    .Q(\memory[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3898_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net562),
    .Q(\S8x305.regs[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3899_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0215_),
    .Q(\S8x305.regs[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3900_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0216_),
    .Q(\S8x305.regs[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3901_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0217_),
    .Q(\S8x305.regs[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3902_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0218_),
    .Q(\S8x305.regs[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3903_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0219_),
    .Q(\S8x305.regs[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3904_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0220_),
    .Q(\S8x305.regs[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3905_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0221_),
    .Q(\S8x305.regs[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3906_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0222_),
    .Q(\S8x305.I[12] ));
 sky130_fd_sc_hd__dfxtp_1 _3907_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0223_),
    .Q(\S8x305.I[13] ));
 sky130_fd_sc_hd__dfxtp_1 _3908_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0224_),
    .Q(\S8x305.I[14] ));
 sky130_fd_sc_hd__dfxtp_1 _3909_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0225_),
    .Q(\S8x305.I[15] ));
 sky130_fd_sc_hd__dfxtp_1 _3910_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0226_),
    .Q(\S8x305.I[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3911_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0227_),
    .Q(\S8x305.I[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3912_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0228_),
    .Q(\S8x305.I[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3913_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0229_),
    .Q(\S8x305.I[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3914_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0230_),
    .Q(\S8x305.I[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3915_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0231_),
    .Q(\S8x305.I[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3916_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0232_),
    .Q(\S8x305.I[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3917_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0233_),
    .Q(\S8x305.I[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3918_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net779),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_1 _3919_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0235_),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_1 _3920_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0236_),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_1 _3921_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net644),
    .Q(\S8x305.regs[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3922_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0238_),
    .Q(\S8x305.regs[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3923_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0239_),
    .Q(\S8x305.regs[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3924_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0240_),
    .Q(\S8x305.regs[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3925_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0241_),
    .Q(\S8x305.regs[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3926_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0242_),
    .Q(\S8x305.regs[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3927_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0243_),
    .Q(\S8x305.regs[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3928_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net660),
    .Q(\S8x305.regs[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3929_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net520),
    .Q(\S8x305.regs[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3930_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0246_),
    .Q(\S8x305.regs[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3931_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0247_),
    .Q(\S8x305.regs[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3932_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0248_),
    .Q(\S8x305.regs[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3933_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0249_),
    .Q(\S8x305.regs[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3934_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0250_),
    .Q(\S8x305.regs[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3935_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0251_),
    .Q(\S8x305.regs[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3936_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net504),
    .Q(\S8x305.regs[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3937_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net542),
    .Q(\S8x305.regs[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3938_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0254_),
    .Q(\S8x305.regs[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3939_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0255_),
    .Q(\S8x305.regs[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3940_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0256_),
    .Q(\S8x305.regs[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3941_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0257_),
    .Q(\S8x305.regs[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3942_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0258_),
    .Q(\S8x305.regs[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3943_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0259_),
    .Q(\S8x305.regs[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3944_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0260_),
    .Q(\S8x305.regs[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3945_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net361),
    .Q(\memory[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3946_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net343),
    .Q(\memory[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3947_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net285),
    .Q(\memory[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3948_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net349),
    .Q(\memory[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3949_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net365),
    .Q(\memory[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3950_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net279),
    .Q(\memory[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3951_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net205),
    .Q(\memory[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3952_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net221),
    .Q(\memory[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3953_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net197),
    .Q(\memory[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3954_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net291),
    .Q(\memory[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3955_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net133),
    .Q(\memory[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3956_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net219),
    .Q(\memory[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3957_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net223),
    .Q(\memory[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3958_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net233),
    .Q(\memory[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3959_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net137),
    .Q(\memory[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3960_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net253),
    .Q(\memory[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3961_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net307),
    .Q(\memory[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3962_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net269),
    .Q(\memory[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3963_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net173),
    .Q(\memory[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3964_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net313),
    .Q(\memory[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3965_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net351),
    .Q(\memory[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3966_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net319),
    .Q(\memory[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3967_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net265),
    .Q(\memory[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3968_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net295),
    .Q(\memory[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3969_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net287),
    .Q(\memory[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3970_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net225),
    .Q(\memory[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3971_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net389),
    .Q(\memory[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3972_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net187),
    .Q(\memory[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3973_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net359),
    .Q(\memory[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3974_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net275),
    .Q(\memory[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3975_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net345),
    .Q(\memory[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3976_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net333),
    .Q(\memory[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3977_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net227),
    .Q(\memory[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3978_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net281),
    .Q(\memory[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3979_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net213),
    .Q(\memory[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3980_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net163),
    .Q(\memory[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3981_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net263),
    .Q(\memory[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3982_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net207),
    .Q(\memory[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3983_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net245),
    .Q(\memory[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3984_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net217),
    .Q(\memory[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3985_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net171),
    .Q(\memory[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3986_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net229),
    .Q(\memory[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3987_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net201),
    .Q(\memory[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3988_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net183),
    .Q(\memory[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3989_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net175),
    .Q(\memory[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3990_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net337),
    .Q(\memory[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3991_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net189),
    .Q(\memory[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3992_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net203),
    .Q(\memory[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3993_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net353),
    .Q(\memory[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3994_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net243),
    .Q(\memory[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3995_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net167),
    .Q(\memory[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3996_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net235),
    .Q(\memory[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3997_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net327),
    .Q(\memory[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3998_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net237),
    .Q(\memory[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3999_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net247),
    .Q(\memory[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4000_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net199),
    .Q(\memory[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4001_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net317),
    .Q(\memory[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4002_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net155),
    .Q(\memory[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4003_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net131),
    .Q(\memory[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4004_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net165),
    .Q(\memory[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4005_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net231),
    .Q(\memory[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4006_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net325),
    .Q(\memory[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4007_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net127),
    .Q(\memory[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4008_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net191),
    .Q(\memory[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4009_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0325_),
    .Q(\memory[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4010_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net402),
    .Q(\memory[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4011_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net395),
    .Q(\memory[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4012_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net412),
    .Q(\memory[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4013_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net397),
    .Q(\memory[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4014_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0330_),
    .Q(\memory[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4015_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net399),
    .Q(\memory[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4016_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net404),
    .Q(\memory[5][7] ));
 sky130_fd_sc_hd__dfxtp_2 _4017_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net703),
    .Q(\ROM_addr_buff[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4018_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0334_),
    .Q(\ROM_addr_buff[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4019_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0335_),
    .Q(\ROM_addr_buff[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4020_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0336_),
    .Q(\ROM_addr_buff[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4021_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0337_),
    .Q(\ROM_addr_buff[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4022_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0338_),
    .Q(\ROM_addr_buff[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4023_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0339_),
    .Q(\ROM_addr_buff[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4024_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0340_),
    .Q(\ROM_addr_buff[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4025_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net371),
    .Q(\ROM_addr_buff[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4026_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0342_),
    .Q(\ROM_addr_buff[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4027_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0343_),
    .Q(\ROM_addr_buff[11] ));
 sky130_fd_sc_hd__dfxtp_1 _4028_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0344_),
    .Q(\ROM_addr_buff[12] ));
 sky130_fd_sc_hd__dfxtp_1 _4029_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0345_),
    .Q(\ROM_addr_buff[13] ));
 sky130_fd_sc_hd__dfxtp_1 _4030_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net741),
    .Q(\S8x305.A[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4031_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net787),
    .Q(\S8x305.A[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4032_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0348_),
    .Q(\S8x305.A[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4033_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0349_),
    .Q(\S8x305.A[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4034_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0350_),
    .Q(\S8x305.A[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4035_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0351_),
    .Q(\S8x305.A[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4036_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0352_),
    .Q(\S8x305.A[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4037_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0353_),
    .Q(\S8x305.A[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4038_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net490),
    .Q(\S8x305.A[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4039_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net442),
    .Q(\S8x305.A[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4040_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0356_),
    .Q(\S8x305.A[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4041_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net123),
    .Q(\S8x305.A[11] ));
 sky130_fd_sc_hd__dfxtp_1 _4042_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net446),
    .Q(\S8x305.A[12] ));
 sky130_fd_sc_hd__dfxtp_1 _4043_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0359_),
    .Q(\S8x305.PC[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4044_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0360_),
    .Q(\S8x305.PC[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4045_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net471),
    .Q(\S8x305.PC[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4046_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0362_),
    .Q(\S8x305.PC[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4047_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net743),
    .Q(\S8x305.PC[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4048_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0364_),
    .Q(\S8x305.cycle[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4049_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0365_),
    .Q(\S8x305.cycle[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4050_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net259),
    .Q(\memory[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4051_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net273),
    .Q(\memory[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4052_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net283),
    .Q(\memory[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4053_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net193),
    .Q(\memory[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4054_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net185),
    .Q(\memory[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4055_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net145),
    .Q(\memory[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4056_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net347),
    .Q(\memory[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4057_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net315),
    .Q(\memory[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4058_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net385),
    .Q(\memory[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4059_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net367),
    .Q(\memory[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4060_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net357),
    .Q(\memory[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4061_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net305),
    .Q(\memory[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4062_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net381),
    .Q(\memory[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4063_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net271),
    .Q(\memory[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4064_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net355),
    .Q(\memory[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4065_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net267),
    .Q(\memory[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4066_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net341),
    .Q(\memory[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4067_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net309),
    .Q(\memory[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4068_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net249),
    .Q(\memory[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4069_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net331),
    .Q(\memory[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4070_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net277),
    .Q(\memory[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4071_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net329),
    .Q(\memory[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4072_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net289),
    .Q(\memory[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4073_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net383),
    .Q(\memory[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4074_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net297),
    .Q(\memory[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4075_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net321),
    .Q(\memory[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4076_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net261),
    .Q(\memory[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4077_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net179),
    .Q(\memory[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4078_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net239),
    .Q(\memory[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4079_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net257),
    .Q(\memory[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4080_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net211),
    .Q(\memory[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4081_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net161),
    .Q(\memory[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4082_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0398_),
    .Q(\S8x305.ALU_in1[0] ));
 sky130_fd_sc_hd__dfxtp_2 _4083_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0399_),
    .Q(\S8x305.ALU_in1[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4084_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0400_),
    .Q(\S8x305.ALU_in1[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4085_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0401_),
    .Q(\S8x305.ALU_in1[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4086_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0402_),
    .Q(\S8x305.ALU_in1[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4087_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0403_),
    .Q(\S8x305.ALU_in1[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4088_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0404_),
    .Q(\S8x305.ALU_in1[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4089_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0405_),
    .Q(\S8x305.ALU_in1[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4090_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net438),
    .Q(\S8x305.i_latch[0] ));
 sky130_fd_sc_hd__dfxtp_1 _4091_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net391),
    .Q(\S8x305.i_latch[1] ));
 sky130_fd_sc_hd__dfxtp_1 _4092_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net379),
    .Q(\S8x305.i_latch[2] ));
 sky130_fd_sc_hd__dfxtp_1 _4093_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net434),
    .Q(\S8x305.i_latch[3] ));
 sky130_fd_sc_hd__dfxtp_1 _4094_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0410_),
    .Q(\S8x305.i_latch[4] ));
 sky130_fd_sc_hd__dfxtp_1 _4095_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net387),
    .Q(\S8x305.i_latch[5] ));
 sky130_fd_sc_hd__dfxtp_1 _4096_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net452),
    .Q(\S8x305.i_latch[6] ));
 sky130_fd_sc_hd__dfxtp_1 _4097_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0413_),
    .Q(\S8x305.i_latch[7] ));
 sky130_fd_sc_hd__dfxtp_1 _4098_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net408),
    .Q(\S8x305.i_latch[8] ));
 sky130_fd_sc_hd__dfxtp_1 _4099_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net687),
    .Q(\S8x305.i_latch[9] ));
 sky130_fd_sc_hd__dfxtp_1 _4100_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net714),
    .Q(\S8x305.i_latch[10] ));
 sky130_fd_sc_hd__dfxtp_1 _4101_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net685),
    .Q(\S8x305.i_latch[11] ));
 sky130_fd_sc_hd__dfxtp_1 _4102_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net450),
    .Q(\S8x305.i_latch[12] ));
 sky130_fd_sc_hd__dfxtp_1 _4103_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net460),
    .Q(\S8x305.i_latch[13] ));
 sky130_fd_sc_hd__dfxtp_1 _4104_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0420_),
    .Q(\S8x305.i_latch[14] ));
 sky130_fd_sc_hd__dfxtp_1 _4105_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net159),
    .Q(\S8x305.i_latch[15] ));
 sky130_fd_sc_hd__dfxtp_1 _4106_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net177),
    .Q(\memory[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4107_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net181),
    .Q(\memory[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4108_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net149),
    .Q(\memory[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4109_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net335),
    .Q(\memory[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4110_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net373),
    .Q(\memory[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4111_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net293),
    .Q(\memory[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4112_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net143),
    .Q(\memory[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4113_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net251),
    .Q(\memory[9][7] ));
 sky130_fd_sc_hd__buf_1 _4122_ (.A(net28),
    .X(net25));
 sky130_fd_sc_hd__buf_1 _4123_ (.A(net28),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_4 fanout100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_4 fanout101 (.A(net102),
    .X(net101));
 sky130_fd_sc_hd__buf_2 fanout102 (.A(net23),
    .X(net102));
 sky130_fd_sc_hd__buf_4 fanout103 (.A(net104),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_4 fanout104 (.A(net113),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_4 fanout105 (.A(net113),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_2 fanout106 (.A(net113),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_4 fanout107 (.A(net108),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_4 fanout108 (.A(net113),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_4 fanout109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_4 fanout110 (.A(net112),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_4 fanout111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_2 fanout112 (.A(net113),
    .X(net112));
 sky130_fd_sc_hd__buf_4 fanout113 (.A(net23),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_8 fanout57 (.A(net58),
    .X(net57));
 sky130_fd_sc_hd__buf_4 fanout58 (.A(_1295_),
    .X(net58));
 sky130_fd_sc_hd__buf_4 fanout59 (.A(_0466_),
    .X(net59));
 sky130_fd_sc_hd__buf_6 fanout60 (.A(_1829_),
    .X(net60));
 sky130_fd_sc_hd__buf_4 fanout61 (.A(_1823_),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_8 fanout62 (.A(_1802_),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_8 fanout63 (.A(_1798_),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_8 fanout64 (.A(net821),
    .X(net64));
 sky130_fd_sc_hd__buf_6 fanout65 (.A(net66),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_8 fanout66 (.A(_1824_),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_8 fanout67 (.A(net68),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_8 fanout68 (.A(net71),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_8 fanout69 (.A(net71),
    .X(net69));
 sky130_fd_sc_hd__buf_4 fanout70 (.A(net71),
    .X(net70));
 sky130_fd_sc_hd__buf_4 fanout71 (.A(_1812_),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_8 fanout72 (.A(net73),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_8 fanout73 (.A(_1801_),
    .X(net73));
 sky130_fd_sc_hd__buf_4 fanout74 (.A(net30),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_8 fanout75 (.A(net56),
    .X(net75));
 sky130_fd_sc_hd__buf_4 fanout76 (.A(net55),
    .X(net76));
 sky130_fd_sc_hd__buf_4 fanout77 (.A(net54),
    .X(net77));
 sky130_fd_sc_hd__buf_4 fanout78 (.A(net53),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_8 fanout79 (.A(net52),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_8 fanout80 (.A(net51),
    .X(net80));
 sky130_fd_sc_hd__buf_4 fanout81 (.A(net50),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_8 fanout82 (.A(net784),
    .X(net82));
 sky130_fd_sc_hd__buf_2 fanout83 (.A(net784),
    .X(net83));
 sky130_fd_sc_hd__buf_6 fanout84 (.A(net488),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_4 fanout85 (.A(net86),
    .X(net85));
 sky130_fd_sc_hd__buf_4 fanout86 (.A(_0002_),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_8 fanout87 (.A(net88),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_8 fanout88 (.A(_0001_),
    .X(net88));
 sky130_fd_sc_hd__buf_6 fanout89 (.A(net90),
    .X(net89));
 sky130_fd_sc_hd__buf_8 fanout90 (.A(_0000_),
    .X(net90));
 sky130_fd_sc_hd__buf_4 fanout91 (.A(_1771_),
    .X(net91));
 sky130_fd_sc_hd__buf_2 fanout92 (.A(_1771_),
    .X(net92));
 sky130_fd_sc_hd__buf_4 fanout93 (.A(net94),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_4 fanout94 (.A(net98),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_4 fanout95 (.A(net98),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_4 fanout96 (.A(net98),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_4 fanout97 (.A(net98),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_4 fanout98 (.A(net23),
    .X(net98));
 sky130_fd_sc_hd__buf_4 fanout99 (.A(net100),
    .X(net99));
 sky130_fd_sc_hd__buf_1 hold1 (.A(net869),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0319_),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_0268_),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\memory[11][4] ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_0273_),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\memory[0][1] ),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_0286_),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\memory[8][0] ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_0293_),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\memory[7][1] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_0302_),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\memory[4][4] ),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\memory[11][2] ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_0321_),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\memory[11][5] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_0274_),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\memory[6][3] ),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_0312_),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\memory[6][5] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_0314_),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\memory[15][4] ),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_0394_),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\memory[13][6] ),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0271_),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_0212_),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\memory[6][1] ),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_0310_),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\memory[8][6] ),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_0299_),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\memory[6][6] ),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(_0315_),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\memory[1][2] ),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(_0384_),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\memory[9][7] ),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\memory[13][3] ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_0429_),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\memory[11][7] ),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_0276_),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\memory[13][7] ),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(_0213_),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\memory[15][5] ),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_0395_),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\memory[3][0] ),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_0366_),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\memory[15][2] ),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0209_),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(_0392_),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\memory[8][4] ),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_0297_),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\memory[10][6] ),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_0283_),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\memory[2][7] ),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_0381_),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\memory[10][1] ),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_0278_),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\memory[2][5] ),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\memory[11][6] ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(_0379_),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\memory[3][1] ),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_0367_),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\memory[0][5] ),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(_0290_),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\memory[1][4] ),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_0386_),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\memory[12][5] ),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_0266_),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\memory[8][1] ),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_0275_),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(_0294_),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\memory[3][2] ),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_0368_),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\memory[12][2] ),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_0263_),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\memory[0][0] ),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_0285_),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\memory[1][6] ),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(_0388_),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\memory[11][1] ),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\memory[13][4] ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_0270_),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\memory[9][5] ),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_0427_),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\memory[10][7] ),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(_0284_),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\memory[15][0] ),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(_0390_),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\memory[13][2] ),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_0208_),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\memory[14][5] ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_0210_),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(_0017_),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\memory[14][6] ),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(_0018_),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\memory[2][3] ),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(_0377_),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\memory[10][0] ),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(_0277_),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\memory[1][1] ),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(_0383_),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\memory[14][2] ),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\S8x305.regs[8][4] ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(_0014_),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\memory[10][3] ),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(_0280_),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\memory[3][7] ),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(_0373_),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\memory[4][0] ),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(_0317_),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\memory[10][5] ),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(_0282_),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\memory[15][1] ),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0357_),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_0048_),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(_0391_),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\memory[14][7] ),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_0019_),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\memory[4][5] ),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(_0322_),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\memory[6][4] ),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(_0313_),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\memory[1][5] ),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_0387_),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\memory[1][3] ),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\memory[9][6] ),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_0385_),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\memory[0][7] ),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(_0292_),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\memory[9][3] ),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(_0425_),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\memory[7][5] ),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(_0306_),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\memory[14][1] ),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(_0013_),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\memory[1][0] ),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0428_),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(_0382_),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\memory[12][1] ),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(_0262_),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\memory[0][6] ),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(_0291_),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\memory[3][6] ),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(_0372_),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\memory[12][3] ),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(_0264_),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\memory[10][4] ),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\memory[3][5] ),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(_0281_),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\memory[6][0] ),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_0309_),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\memory[2][6] ),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(_0380_),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\memory[2][2] ),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(_0376_),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\memory[0][4] ),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(_0289_),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\memory[12][0] ),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_0371_),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(_0261_),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\memory[14][4] ),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(_0016_),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\memory[12][4] ),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(_0265_),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\memory[2][1] ),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(_0375_),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\memory[13][1] ),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(_0207_),
    .X(net369));
 sky130_fd_sc_hd__buf_1 hold249 (.A(\S8x305.A[8] ),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\S8x305.regs[8][2] ),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(_0341_),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\memory[9][4] ),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(_0426_),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\memory[14][0] ),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(_0012_),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\memory[14][3] ),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(_0015_),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\S8x305.i_latch[2] ),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(_0408_),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\memory[2][4] ),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_0046_),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(_0378_),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\memory[1][7] ),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(_0389_),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\memory[2][0] ),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(_0374_),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\S8x305.i_latch[5] ),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(_0411_),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\memory[0][2] ),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(_0287_),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\S8x305.i_latch[1] ),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\memory[9][2] ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(_0407_),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\ROM_spi_dat_out[0] ),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(_0156_),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\memory[5][2] ),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(_0327_),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\memory[5][4] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(_0329_),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\memory[5][6] ),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_0331_),
    .X(net399));
 sky130_fd_sc_hd__buf_2 hold279 (.A(\S8x305.iv_latch[6] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0424_),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(_1618_),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(_0326_),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\memory[5][7] ),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(_0332_),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\S8x305.I[6] ),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(_0122_),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\S8x305.i_latch[8] ),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(_0414_),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\ROM_spi_dat_out[1] ),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(_0157_),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\memory[13][5] ),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\memory[5][3] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(_0328_),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\ROM_spi_dat_out[3] ),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(_0159_),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\ROM_spi_dat_out[5] ),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(_0161_),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\ROM_spi_dat_out[2] ),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(_0158_),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\ROM_spi_dat_out[4] ),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(_0160_),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\last_addr[0] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0211_),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\S8x305.I[5] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(_0121_),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\ROM_spi_dat_out[7] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(_0163_),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\S8x305.I[4] ),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(_0120_),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\S8x305.I[7] ),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(_0123_),
    .X(net428));
 sky130_fd_sc_hd__buf_2 hold308 (.A(\S8x305.iv_latch[5] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(_0192_),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\S8x305.regs[8][3] ),
    .X(net152));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold310 (.A(\ROM_spi_cycle[2] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(_0135_),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\S8x305.i_latch[3] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(_0409_),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\cmdl[6] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(_0185_),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\S8x305.i_latch[0] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(_0406_),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\cmdr[6] ),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(_0193_),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0047_),
    .X(net153));
 sky130_fd_sc_hd__buf_1 hold320 (.A(net855),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(_0355_),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_2 hold322 (.A(\mem_cycle[2] ),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(_0147_),
    .X(net444));
 sky130_fd_sc_hd__buf_1 hold324 (.A(net857),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(_0358_),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(ROM_OEB),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(_0154_),
    .X(net448));
 sky130_fd_sc_hd__buf_1 hold328 (.A(\S8x305.i_latch[12] ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(_0418_),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\memory[4][1] ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\S8x305.i_latch[6] ),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(_0412_),
    .X(net452));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold332 (.A(net860),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(_1525_),
    .X(net454));
 sky130_fd_sc_hd__buf_1 hold334 (.A(net867),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(_1518_),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(\cmdl[5] ),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(_0184_),
    .X(net458));
 sky130_fd_sc_hd__buf_1 hold338 (.A(\S8x305.i_latch[13] ),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(_0419_),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0318_),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\cmdl[2] ),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(_0181_),
    .X(net462));
 sky130_fd_sc_hd__buf_1 hold342 (.A(net856),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(_1086_),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(_1092_),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\cmdl[7] ),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(_0186_),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\memory[5][5] ),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(_1622_),
    .X(net469));
 sky130_fd_sc_hd__buf_1 hold349 (.A(\S8x305.PC[2] ),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\S8x305.regs[8][7] ),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(_0361_),
    .X(net471));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold351 (.A(\S8x305.PC[7] ),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(_1087_),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(_1088_),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(\cmdr[7] ),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(_0194_),
    .X(net476));
 sky130_fd_sc_hd__clkbuf_2 hold356 (.A(\startup_cycle[1] ),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(_0139_),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\memory[5][0] ),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(_1617_),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_0051_),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\cmdl[4] ),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(_0183_),
    .X(net482));
 sky130_fd_sc_hd__buf_1 hold362 (.A(net865),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(_1520_),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\S8x305.regs[2][3] ),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\cmdl[1] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(_0180_),
    .X(net487));
 sky130_fd_sc_hd__clkbuf_2 hold367 (.A(\S8x305.cycle[0] ),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_4 hold368 (.A(_0487_),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(_0354_),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\S8x305.i_latch[15] ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\S8x305.regs[12][6] ),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\S8x305.regs[6][5] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\S8x305.regs[10][2] ),
    .X(net493));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold373 (.A(\S8x305.A[9] ),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(_1524_),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\cmdl[3] ),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(_0182_),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\S8x305.regs[6][7] ),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\S8x305.regs[1][7] ),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\ROM_spi_dat_out[6] ),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_0421_),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(_1485_),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(_0162_),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\S8x305.regs[2][7] ),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(_0252_),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\cmdr[4] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(_0191_),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\S8x305.regs[10][7] ),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(_0063_),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\S8x305.regs[9][6] ),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\S8x305.regs[11][3] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\memory[15][7] ),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\S8x305.regs[12][1] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(_0089_),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\S8x305.regs[11][0] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(_0072_),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\S8x305.regs[11][5] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\cmdl[0] ),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(_0179_),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\S8x305.regs[13][2] ),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(\S8x305.regs[2][0] ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(_0245_),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0164_),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_0397_),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(\S8x305.regs[11][2] ),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\S8x305.regs[4][1] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(\S8x305.regs[2][1] ),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\S8x305.regs[9][7] ),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(_0119_),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\S8x305.regs[1][6] ),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\S8x305.regs[9][5] ),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\S8x305.regs[10][1] ),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(_0057_),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\S8x305.regs[1][2] ),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\memory[8][3] ),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(\S8x305.regs[12][4] ),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(_0092_),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(\S8x305.regs[9][1] ),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\S8x305.regs[15][2] ),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(\S8x305.regs[12][3] ),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\S8x305.regs[3][4] ),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(\S8x305.regs[7][2] ),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\S8x305.regs[14][6] ),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(\S8x305.regs[7][6] ),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\S8x305.regs[1][1] ),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0296_),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(\S8x305.regs[1][0] ),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(_0253_),
    .X(net542));
 sky130_fd_sc_hd__buf_1 hold422 (.A(net862),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(_1519_),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(\S8x305.regs[11][7] ),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(_0079_),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(\S8x305.regs[2][5] ),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\S8x305.regs[6][6] ),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(\S8x305.regs[2][6] ),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\S8x305.regs[13][3] ),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\memory[4][3] ),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(\S8x305.regs[9][0] ),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(_0112_),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(\S8x305.regs[12][0] ),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(_0088_),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\S8x305.regs[11][4] ),
    .X(net555));
 sky130_fd_sc_hd__clkbuf_2 hold435 (.A(net854),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\S8x305.regs[4][7] ),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\S8x305.regs[5][7] ),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\S8x305.regs[14][1] ),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(_0081_),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_0320_),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\S8x305.regs[4][0] ),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(_0214_),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(\S8x305.regs[10][5] ),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\S8x305.regs[4][5] ),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(\S8x305.regs[1][5] ),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\S8x305.regs[6][2] ),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(\S8x305.regs[14][2] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\S8x305.regs[15][1] ),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(_0065_),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\S8x305.regs[3][6] ),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\memory[6][2] ),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\S8x305.regs[15][3] ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\S8x305.regs[1][3] ),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\S8x305.regs[10][0] ),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(_0056_),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\S8x305.regs[11][1] ),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(_0073_),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\S8x305.regs[7][0] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(_0037_),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\S8x305.regs[9][4] ),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(_0116_),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_0311_),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(\S8x305.regs[12][2] ),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\S8x305.regs[3][5] ),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\S8x305.regs[5][2] ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\S8x305.regs[9][3] ),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\S8x305.regs[5][6] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\S8x305.regs[6][3] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\S8x305.regs[3][3] ),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\S8x305.regs[5][3] ),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\S8x305.regs[14][3] ),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\S8x305.regs[7][3] ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\S8x305.regs[8][1] ),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(\S8x305.regs[15][6] ),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\S8x305.regs[1][4] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\S8x305.regs[13][7] ),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(_0111_),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\S8x305.regs[4][4] ),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\S8x305.regs[10][6] ),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\S8x305.regs[13][6] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\S8x305.regs[7][4] ),
    .X(net598));
 sky130_fd_sc_hd__clkbuf_4 hold478 (.A(net40),
    .X(net599));
 sky130_fd_sc_hd__buf_2 hold479 (.A(_0486_),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_0045_),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(_1705_),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\S8x305.regs[15][7] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(_0071_),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\S8x305.regs[13][4] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(_0108_),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\S8x305.regs[14][4] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(_0084_),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\S8x305.regs[11][6] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\S8x305.regs[5][1] ),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\S8x305.regs[2][2] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\memory[7][0] ),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\S8x305.regs[12][7] ),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(_0095_),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\S8x305.regs[6][1] ),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\S8x305.regs[4][6] ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\S8x305.regs[7][7] ),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\S8x305.regs[14][5] ),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(\S8x305.regs[2][4] ),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\S8x305.regs[12][5] ),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(\S8x305.regs[7][1] ),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(net44),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\memory[4][6] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_0301_),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(_0126_),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\S8x305.regs[6][0] ),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(_0025_),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\S8x305.regs[5][5] ),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(\S8x305.regs[5][4] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(_0100_),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(\S8x305.regs[3][1] ),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\S8x305.regs[6][4] ),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(_0029_),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\S8x305.regs[10][4] ),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\memory[10][2] ),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(_0060_),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\S8x305.regs[3][2] ),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(net43),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(_0125_),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(\S8x305.regs[15][5] ),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\S8x305.regs[10][3] ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(\S8x305.regs[4][3] ),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\S8x305.regs[13][5] ),
    .X(net638));
 sky130_fd_sc_hd__buf_1 hold518 (.A(net863),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(_1521_),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_0279_),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_2 hold520 (.A(\S8x305.iv_latch[1] ),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(_0188_),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(\S8x305.regs[3][0] ),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(_0237_),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(\S8x305.regs[4][2] ),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\S8x305.regs[15][0] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(_0064_),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\S8x305.regs[14][7] ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(_0087_),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\S8x305.regs[13][1] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\memory[7][4] ),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(\S8x305.regs[15][4] ),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\S8x305.regs[7][5] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(\S8x305.regs[14][0] ),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(_0080_),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(\S8x305.regs[13][0] ),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(_0104_),
    .X(net656));
 sky130_fd_sc_hd__buf_1 hold536 (.A(net46),
    .X(net657));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold537 (.A(_0128_),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(\S8x305.regs[3][7] ),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(_0244_),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_0305_),
    .X(net175));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold540 (.A(\startup_cycle[3] ),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(_0141_),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(\S8x305.I[14] ),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(_1543_),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(net48),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\cmdr[1] ),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(_0034_),
    .X(net667));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold547 (.A(net47),
    .X(net668));
 sky130_fd_sc_hd__buf_1 hold548 (.A(_0129_),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(\last_addr[9] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\memory[9][0] ),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(_1498_),
    .X(net671));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold551 (.A(net859),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(_1523_),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(\last_addr[5] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(_1494_),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(\S8x305.I[10] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(_1548_),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\S8x305.I[8] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(_1546_),
    .X(net679));
 sky130_fd_sc_hd__clkbuf_2 hold559 (.A(\S8x305.iv_latch[0] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_0422_),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(_0033_),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\last_addr[10] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(_0174_),
    .X(net683));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold563 (.A(\S8x305.i_latch[11] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(_0417_),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\S8x305.i_latch[9] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(_0415_),
    .X(net687));
 sky130_fd_sc_hd__buf_1 hold567 (.A(\ROM_spi_cycle[4] ),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(_0137_),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\cmdr[0] ),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\memory[15][3] ),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(_0187_),
    .X(net691));
 sky130_fd_sc_hd__buf_1 hold571 (.A(\ROM_addr_buff[3] ),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(\ROM_spi_cycle[3] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(_1328_),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(_0136_),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\last_addr[3] ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(_0167_),
    .X(net697));
 sky130_fd_sc_hd__buf_2 hold577 (.A(\startup_cycle[4] ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(_1340_),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(_0142_),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_0393_),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(\S8x305.i_latch[6] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\S8x305.A[0] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(_0333_),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(net45),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(_0127_),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\S8x305.regs[5][0] ),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(_0096_),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\last_A[12] ),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(_1527_),
    .X(net709));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold589 (.A(net858),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\memory[9][1] ),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(\last_addr[7] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(_1496_),
    .X(net712));
 sky130_fd_sc_hd__buf_1 hold592 (.A(\S8x305.i_latch[10] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(_0416_),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(\S8x305.regs[9][2] ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\last_addr[12] ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(_0176_),
    .X(net717));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold597 (.A(\ROM_addr_buff[11] ),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(net49),
    .X(net719));
 sky130_fd_sc_hd__clkbuf_2 hold599 (.A(\startup_cycle[6] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0323_),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_0423_),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(_0144_),
    .X(net721));
 sky130_fd_sc_hd__buf_2 hold601 (.A(\startup_cycle[5] ),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(_0143_),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\last_A[11] ),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(_1526_),
    .X(net725));
 sky130_fd_sc_hd__clkbuf_2 hold605 (.A(net861),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(_1321_),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(_0133_),
    .X(net728));
 sky130_fd_sc_hd__buf_1 hold608 (.A(\S8x305.PC[5] ),
    .X(net729));
 sky130_fd_sc_hd__clkbuf_2 hold609 (.A(\S8x305.iv_latch[3] ),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\memory[7][3] ),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(_0190_),
    .X(net731));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold611 (.A(\S8x305.I[2] ),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(_1553_),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\cmdr[3] ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(_0036_),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\ROM_addr_buff[8] ),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(\S8x305.PC[7] ),
    .X(net737));
 sky130_fd_sc_hd__clkbuf_2 hold617 (.A(net866),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(_0177_),
    .X(net739));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold619 (.A(net868),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_0304_),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(_0346_),
    .X(net741));
 sky130_fd_sc_hd__buf_1 hold621 (.A(\S8x305.PC[4] ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(_0363_),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(net41),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(_0151_),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\S8x305.I[1] ),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(_1552_),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\S8x305.I[9] ),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(_1547_),
    .X(net749));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold629 (.A(\S8x305.PC[3] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\memory[3][4] ),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(\last_A[1] ),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(_1517_),
    .X(net752));
 sky130_fd_sc_hd__buf_1 hold632 (.A(net864),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(_1522_),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(\S8x305.I[13] ),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(_1542_),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(\S8x305.i_latch[4] ),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\ROM_addr_buff[4] ),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(\S8x305.iv_latch[4] ),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\S8x305.i_latch[14] ),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_0370_),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(\ROM_addr_buff[5] ),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\last_addr[4] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(_0168_),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(net29),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(_0132_),
    .X(net765));
 sky130_fd_sc_hd__buf_1 hold645 (.A(\ROM_addr_buff[6] ),
    .X(net766));
 sky130_fd_sc_hd__buf_1 hold646 (.A(\ROM_addr_buff[10] ),
    .X(net767));
 sky130_fd_sc_hd__clkbuf_2 hold647 (.A(\startup_cycle[0] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(_1336_),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(_0138_),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\memory[0][3] ),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(\S8x305.ALU_in1[7] ),
    .X(net771));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold651 (.A(\S8x305.I[0] ),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(\S8x305.A[12] ),
    .X(net773));
 sky130_fd_sc_hd__buf_1 hold653 (.A(\last_addr[11] ),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(_0175_),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\S8x305.I[11] ),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(_1549_),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(net37),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(_0234_),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(\ROM_addr_buff[1] ),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_0288_),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(_1490_),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(\S8x305.I[15] ),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(_1544_),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\S8x305.cycle[1] ),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(_0011_),
    .X(net785));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold665 (.A(\S8x305.A[1] ),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(_0347_),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(\S8x305.ALU_in1[6] ),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(\S8x305.ALU_in1[0] ),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(\ROM_addr_buff[7] ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\memory[7][6] ),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(\last_addr[8] ),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(_1497_),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(\S8x305.iv_latch[7] ),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(\S8x305.I[3] ),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(_1554_),
    .X(net795));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold675 (.A(\mem_cycle[1] ),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(_1430_),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(\last_addr[6] ),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(_1495_),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(\S8x305.PC[6] ),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_0307_),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(\S8x305.PC[1] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(\last_addr[2] ),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(_1491_),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(\S8x305.I[12] ),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(\S8x305.ALU_in1[4] ),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(\startup_cycle[2] ),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(_1339_),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(_0140_),
    .X(net808));
 sky130_fd_sc_hd__buf_1 hold688 (.A(\S8x305.iv_latch[2] ),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(_0189_),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\memory[4][7] ),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(\cmdr[2] ),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(\S8x305.ALU_in1[5] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(\S8x305.ALU_in1[2] ),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(\S8x305.ALU_in1[3] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(\S8x305.A[11] ),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(_1636_),
    .X(net816));
 sky130_fd_sc_hd__buf_1 hold696 (.A(\ROM_spi_cycle[1] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(_1323_),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(_0134_),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(\ROM_spi_cycle[0] ),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\S8x305.regs[8][6] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_0324_),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(_1252_),
    .X(net821));
 sky130_fd_sc_hd__buf_1 hold701 (.A(\mem_cycle[4] ),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(_1402_),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(_1403_),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(\S8x305.regs[8][0] ),
    .X(net825));
 sky130_fd_sc_hd__clkbuf_2 hold705 (.A(\mem_cycle[5] ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(_1293_),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(net38),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(_1565_),
    .X(net829));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold709 (.A(\mem_cycle[3] ),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\memory[3][3] ),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(_1399_),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(_0148_),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(net36),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(_1459_),
    .X(net834));
 sky130_fd_sc_hd__clkbuf_2 hold714 (.A(\mem_cycle[0] ),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(\last_A[10] ),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(_1274_),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(_1282_),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(net39),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(_1569_),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_0369_),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(\ROM_addr_buff[12] ),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(_1394_),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(_0145_),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(\ROM_addr_buff[2] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(\S8x305.ALU_in1[1] ),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(net42),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(_1443_),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(\mem_cycle[1] ),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(\memory[5][1] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(\ROM_addr_buff[10] ),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\memory[13][0] ),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(\S8x305.iv_latch[1] ),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(\S8x305.iv_latch[1] ),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(\S8x305.PC[10] ),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(\S8x305.PC[9] ),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(\S8x305.PC[8] ),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(\S8x305.PC[12] ),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(\S8x305.i_latch[7] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(\S8x305.A[7] ),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(\S8x305.A[10] ),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(spi_clkdiv),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_0206_),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(\S8x305.A[3] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(\S8x305.A[5] ),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(\S8x305.A[6] ),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(\S8x305.A[4] ),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(\ROM_addr_buff[13] ),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(\S8x305.A[2] ),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(\S8x305.PC[0] ),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(\S8x305.PC[11] ),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\memory[11][0] ),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_0269_),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\memory[6][7] ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_0316_),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\memory[7][2] ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0050_),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_0303_),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\memory[7][7] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0308_),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\memory[12][6] ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0267_),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\memory[8][5] ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_0298_),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\S8x305.regs[8][5] ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(_0049_),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\memory[15][6] ),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\memory[4][2] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_0396_),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\memory[8][2] ),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_0295_),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(ROM_spi_mode),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_0155_),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\memory[8][7] ),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_0300_),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\memory[11][3] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_0272_),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\memory[12][7] ),
    .X(net220));
 sky130_fd_sc_hd__buf_1 input1 (.A(custom_settings[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(io_in[24]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(io_in[25]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(io_in[26]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(io_in[27]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(io_in[28]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(io_in[2]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(io_in[3]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(io_in[4]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(io_in[5]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(io_in[6]),
    .X(net19));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(custom_settings[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(io_in[7]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(io_in[8]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(io_in[9]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(rst_n),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(io_in[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(io_in[16]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(io_in[17]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(io_in[18]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(io_in[19]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(io_in[22]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(io_in[23]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 load_slew1 (.A(_1793_),
    .X(net853));
 sky130_fd_sc_hd__buf_12 output24 (.A(net24),
    .X(io_oeb[0]));
 sky130_fd_sc_hd__buf_12 output25 (.A(net25),
    .X(io_oeb[1]));
 sky130_fd_sc_hd__buf_12 output26 (.A(net26),
    .X(io_oeb[2]));
 sky130_fd_sc_hd__buf_12 output27 (.A(net27),
    .X(io_oeb[3]));
 sky130_fd_sc_hd__buf_12 output28 (.A(net28),
    .X(io_oeb[4]));
 sky130_fd_sc_hd__buf_12 output29 (.A(net29),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_12 output30 (.A(net74),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_12 output31 (.A(net31),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_12 output32 (.A(net32),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_12 output33 (.A(net33),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_12 output34 (.A(net34),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_12 output35 (.A(net35),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_12 output36 (.A(net36),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_12 output37 (.A(net37),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_12 output38 (.A(net38),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_12 output39 (.A(net39),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_12 output40 (.A(net40),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_12 output41 (.A(net41),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_12 output42 (.A(net42),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_12 output43 (.A(net43),
    .X(io_out[29]));
 sky130_fd_sc_hd__buf_12 output44 (.A(net44),
    .X(io_out[30]));
 sky130_fd_sc_hd__buf_12 output45 (.A(net45),
    .X(io_out[31]));
 sky130_fd_sc_hd__buf_12 output46 (.A(net46),
    .X(io_out[32]));
 sky130_fd_sc_hd__buf_12 output47 (.A(net47),
    .X(io_out[33]));
 sky130_fd_sc_hd__buf_12 output48 (.A(net48),
    .X(io_out[34]));
 sky130_fd_sc_hd__buf_12 output49 (.A(net49),
    .X(io_out[35]));
 sky130_fd_sc_hd__buf_12 output50 (.A(net81),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_12 output51 (.A(net80),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_12 output52 (.A(net79),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_12 output53 (.A(net78),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_12 output54 (.A(net77),
    .X(io_out[7]));
 sky130_fd_sc_hd__buf_12 output55 (.A(net76),
    .X(io_out[8]));
 sky130_fd_sc_hd__buf_12 output56 (.A(net75),
    .X(io_out[9]));
 sky130_fd_sc_hd__conb_1 wrapped_8x305_114 (.LO(net114));
 sky130_fd_sc_hd__conb_1 wrapped_8x305_115 (.LO(net115));
 sky130_fd_sc_hd__conb_1 wrapped_8x305_116 (.LO(net116));
 sky130_fd_sc_hd__conb_1 wrapped_8x305_117 (.LO(net117));
 sky130_fd_sc_hd__conb_1 wrapped_8x305_118 (.LO(net118));
 sky130_fd_sc_hd__conb_1 wrapped_8x305_119 (.LO(net119));
 sky130_fd_sc_hd__conb_1 wrapped_8x305_120 (.LO(net120));
 sky130_fd_sc_hd__conb_1 wrapped_8x305_121 (.HI(net121));
 assign io_out[22] = net114;
 assign io_out[23] = net115;
 assign io_out[24] = net116;
 assign io_out[25] = net117;
 assign io_out[26] = net118;
 assign io_out[27] = net119;
 assign io_out[28] = net120;
 assign io_out[2] = net121;
endmodule

