* NGSPICE file created from execution_unit.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_2 abstract view
.subckt sky130_fd_sc_hd__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt execution_unit busy curr_PC[0] curr_PC[10] curr_PC[11] curr_PC[12] curr_PC[13]
+ curr_PC[14] curr_PC[15] curr_PC[16] curr_PC[17] curr_PC[18] curr_PC[19] curr_PC[1]
+ curr_PC[20] curr_PC[21] curr_PC[22] curr_PC[23] curr_PC[24] curr_PC[25] curr_PC[26]
+ curr_PC[27] curr_PC[2] curr_PC[3] curr_PC[4] curr_PC[5] curr_PC[6] curr_PC[7] curr_PC[8]
+ curr_PC[9] dest_idx[0] dest_idx[1] dest_idx[2] dest_idx[3] dest_idx[4] dest_idx[5]
+ dest_mask[0] dest_mask[1] dest_pred[0] dest_pred[1] dest_pred[2] dest_pred_val dest_val[0]
+ dest_val[10] dest_val[11] dest_val[12] dest_val[13] dest_val[14] dest_val[15] dest_val[16]
+ dest_val[17] dest_val[18] dest_val[19] dest_val[1] dest_val[20] dest_val[21] dest_val[22]
+ dest_val[23] dest_val[24] dest_val[25] dest_val[26] dest_val[27] dest_val[28] dest_val[29]
+ dest_val[2] dest_val[30] dest_val[31] dest_val[3] dest_val[4] dest_val[5] dest_val[6]
+ dest_val[7] dest_val[8] dest_val[9] instruction[0] instruction[10] instruction[11]
+ instruction[12] instruction[13] instruction[14] instruction[15] instruction[16]
+ instruction[17] instruction[18] instruction[19] instruction[1] instruction[20] instruction[21]
+ instruction[22] instruction[23] instruction[24] instruction[25] instruction[26]
+ instruction[27] instruction[28] instruction[29] instruction[2] instruction[30] instruction[31]
+ instruction[32] instruction[33] instruction[34] instruction[35] instruction[36]
+ instruction[37] instruction[38] instruction[39] instruction[3] instruction[40] instruction[41]
+ instruction[4] instruction[5] instruction[6] instruction[7] instruction[8] instruction[9]
+ int_return is_load is_store loadstore_address[0] loadstore_address[10] loadstore_address[11]
+ loadstore_address[12] loadstore_address[13] loadstore_address[14] loadstore_address[15]
+ loadstore_address[16] loadstore_address[17] loadstore_address[18] loadstore_address[19]
+ loadstore_address[1] loadstore_address[20] loadstore_address[21] loadstore_address[22]
+ loadstore_address[23] loadstore_address[24] loadstore_address[25] loadstore_address[26]
+ loadstore_address[27] loadstore_address[28] loadstore_address[29] loadstore_address[2]
+ loadstore_address[30] loadstore_address[31] loadstore_address[3] loadstore_address[4]
+ loadstore_address[5] loadstore_address[6] loadstore_address[7] loadstore_address[8]
+ loadstore_address[9] loadstore_size[0] loadstore_size[1] new_PC[0] new_PC[10] new_PC[11]
+ new_PC[12] new_PC[13] new_PC[14] new_PC[15] new_PC[16] new_PC[17] new_PC[18] new_PC[19]
+ new_PC[1] new_PC[20] new_PC[21] new_PC[22] new_PC[23] new_PC[24] new_PC[25] new_PC[26]
+ new_PC[27] new_PC[2] new_PC[3] new_PC[4] new_PC[5] new_PC[6] new_PC[7] new_PC[8]
+ new_PC[9] pred_idx[0] pred_idx[1] pred_idx[2] pred_val reg1_idx[0] reg1_idx[1] reg1_idx[2]
+ reg1_idx[3] reg1_idx[4] reg1_idx[5] reg1_val[0] reg1_val[10] reg1_val[11] reg1_val[12]
+ reg1_val[13] reg1_val[14] reg1_val[15] reg1_val[16] reg1_val[17] reg1_val[18] reg1_val[19]
+ reg1_val[1] reg1_val[20] reg1_val[21] reg1_val[22] reg1_val[23] reg1_val[24] reg1_val[25]
+ reg1_val[26] reg1_val[27] reg1_val[28] reg1_val[29] reg1_val[2] reg1_val[30] reg1_val[31]
+ reg1_val[3] reg1_val[4] reg1_val[5] reg1_val[6] reg1_val[7] reg1_val[8] reg1_val[9]
+ reg2_idx[0] reg2_idx[1] reg2_idx[2] reg2_idx[3] reg2_idx[4] reg2_idx[5] reg2_val[0]
+ reg2_val[10] reg2_val[11] reg2_val[12] reg2_val[13] reg2_val[14] reg2_val[15] reg2_val[16]
+ reg2_val[17] reg2_val[18] reg2_val[19] reg2_val[1] reg2_val[20] reg2_val[21] reg2_val[22]
+ reg2_val[23] reg2_val[24] reg2_val[25] reg2_val[26] reg2_val[27] reg2_val[28] reg2_val[29]
+ reg2_val[2] reg2_val[30] reg2_val[31] reg2_val[3] reg2_val[4] reg2_val[5] reg2_val[6]
+ reg2_val[7] reg2_val[8] reg2_val[9] rst sign_extend take_branch vccd1 vssd1 wb_clk_i
XANTENNA__12658__A2 _09520_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09671_ _09453_/X _09455_/X _09671_/S vssd1 vssd1 vccd1 vccd1 _09671_/X sky130_fd_sc_hd__mux2_1
X_06883_ _07281_/A reg1_val[19] vssd1 vssd1 vccd1 vccd1 _06884_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_94_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08622_ _08622_/A _08622_/B vssd1 vssd1 vccd1 vccd1 _08653_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08553_ _08553_/A _08553_/B vssd1 vssd1 vccd1 vccd1 _08555_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout162_A _13196_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07504_ _07504_/A _07653_/A _07504_/C vssd1 vssd1 vccd1 vccd1 _07505_/B sky130_fd_sc_hd__and3_1
XANTENNA__07298__B1 _07521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08484_ _08480_/A _08480_/B _08552_/A vssd1 vssd1 vccd1 vccd1 _08498_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07435_ _07634_/B _07435_/B vssd1 vssd1 vccd1 vccd1 _07435_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07366_ _07367_/A _07367_/B vssd1 vssd1 vccd1 vccd1 _07366_/X sky130_fd_sc_hd__and2_4
XANTENNA__11397__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09105_ _10119_/A _09105_/B vssd1 vssd1 vccd1 vccd1 _09108_/A sky130_fd_sc_hd__xnor2_1
X_07297_ _07297_/A _07521_/A vssd1 vssd1 vccd1 vccd1 _07297_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_32_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09036_ _09031_/A _09031_/B _09035_/X vssd1 vssd1 vccd1 vccd1 _09044_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_115_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07470__B1 _07476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09275__A _09275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07222__B1 _07521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12413__B _12764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09938_ _09938_/A vssd1 vssd1 vccd1 vccd1 _09946_/A sky130_fd_sc_hd__inv_2
XANTENNA__07507__B _07572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09869_ hold262/A hold245/A _12314_/A vssd1 vssd1 vccd1 vccd1 _09870_/B sky130_fd_sc_hd__o21a_1
X_11900_ _07230_/Y _07642_/X fanout13/X _12189_/A vssd1 vssd1 vccd1 vccd1 _11901_/B
+ sky130_fd_sc_hd__a22o_1
X_12880_ _12886_/B _12880_/B vssd1 vssd1 vccd1 vccd1 new_PC[11] sky130_fd_sc_hd__and2_4
X_11831_ _11832_/A _11832_/B vssd1 vssd1 vccd1 vccd1 _11833_/A sky130_fd_sc_hd__or2_1
XFILLER_0_68_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _11553_/X _11950_/A _11760_/X vssd1 vssd1 vccd1 vccd1 _11762_/X sky130_fd_sc_hd__a21o_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ hold291/X _13506_/A2 _13500_/X _13506_/B2 vssd1 vssd1 vccd1 vccd1 _13502_/B
+ sky130_fd_sc_hd__a22o_1
X_10713_ _10713_/A _10713_/B vssd1 vssd1 vccd1 vccd1 _10715_/B sky130_fd_sc_hd__xor2_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ hold231/A _11693_/A2 _11878_/C _12533_/B1 vssd1 vssd1 vccd1 vccd1 _11693_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13432_ hold130/A _13142_/A _13444_/B1 hold95/X _13568_/A vssd1 vssd1 vccd1 vccd1
+ hold96/A sky130_fd_sc_hd__o221a_1
X_10644_ _10780_/B _10644_/B vssd1 vssd1 vccd1 vccd1 _10669_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10575_ _10575_/A _10575_/B vssd1 vssd1 vccd1 vccd1 _10981_/B sky130_fd_sc_hd__xnor2_4
X_13363_ _13543_/A hold175/X vssd1 vssd1 vccd1 vccd1 hold176/A sky130_fd_sc_hd__and2_1
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09450__A1 _10004_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12314_ _12314_/A _12390_/B vssd1 vssd1 vccd1 vccd1 _12314_/X sky130_fd_sc_hd__and2_1
XFILLER_0_106_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13294_ _13498_/B _13499_/A _13259_/X vssd1 vssd1 vccd1 vccd1 _13504_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_51_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12337__A1 _12614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12337__B2 _07257_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12245_ curr_PC[22] _12325_/C _12244_/Y vssd1 vssd1 vccd1 vccd1 _12245_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10348__B1 _10349_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10899__A1 _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12176_ _12420_/A _12176_/B vssd1 vssd1 vccd1 vccd1 _12180_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07764__A1 fanout39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07764__B2 _08118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11127_ _11124_/X _11126_/Y _10995_/X _10999_/X vssd1 vssd1 vccd1 vccd1 _11127_/X
+ sky130_fd_sc_hd__a211o_1
X_11058_ _11059_/A _11059_/B vssd1 vssd1 vccd1 vccd1 _11058_/X sky130_fd_sc_hd__and2_1
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07136__C _13744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10009_ _10006_/X _10008_/X _11472_/S vssd1 vssd1 vccd1 vccd1 _10009_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09269__A1 _09604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09269__B2 _09161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11615__A3 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08492__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07220_ _07213_/A _07213_/B _07521_/A vssd1 vssd1 vccd1 vccd1 _07220_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08264__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07151_ instruction[3] _13748_/A _12738_/S _09520_/B vssd1 vssd1 vccd1 vccd1 _07151_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_14_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08244__A2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10587__B1 _11866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11784__C1 _11783_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07082_ _07082_/A _07082_/B vssd1 vssd1 vccd1 vccd1 _07082_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_124_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout105 _07276_/X vssd1 vssd1 vccd1 vccd1 _10235_/A1 sky130_fd_sc_hd__clkbuf_8
XANTENNA__07755__A1 _08395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout116 _11508_/A vssd1 vssd1 vccd1 vccd1 _09591_/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__07755__B2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout127 _07311_/Y vssd1 vssd1 vccd1 vccd1 _10536_/B2 sky130_fd_sc_hd__buf_4
XANTENNA__10354__A3 _10787_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout138 _11231_/A vssd1 vssd1 vccd1 vccd1 _12695_/A sky130_fd_sc_hd__buf_4
Xfanout149 _13151_/A vssd1 vssd1 vccd1 vccd1 _08923_/B1 sky130_fd_sc_hd__buf_6
X_07984_ _09950_/A _07984_/B vssd1 vssd1 vccd1 vccd1 _07989_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09823__A _09824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09723_ _09656_/B _09656_/C _12742_/A vssd1 vssd1 vccd1 vccd1 _09723_/Y sky130_fd_sc_hd__a21oi_1
X_06935_ _07094_/C vssd1 vssd1 vccd1 vccd1 _11356_/A sky130_fd_sc_hd__inv_2
XANTENNA__13345__A _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09542__B _12825_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09654_ _09654_/A _09654_/B vssd1 vssd1 vccd1 vccd1 _09655_/B sky130_fd_sc_hd__nand2_1
X_06866_ reg2_val[20] _06873_/B1 _06872_/B1 _06865_/Y vssd1 vssd1 vccd1 vccd1 _07201_/A
+ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__08180__A1 _08866_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08180__B2 _09216_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08605_ _08613_/B _08613_/A vssd1 vssd1 vccd1 vccd1 _08605_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__13064__B _13129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09585_ _09948_/A _09585_/B _09585_/C vssd1 vssd1 vccd1 vccd1 _09586_/C sky130_fd_sc_hd__nand3_1
X_06797_ reg2_val[27] _06873_/B1 _06872_/B1 _06796_/Y vssd1 vssd1 vccd1 vccd1 _07251_/A
+ sky130_fd_sc_hd__o2bb2a_2
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08536_ _08608_/A _08548_/B vssd1 vssd1 vccd1 vccd1 _08536_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12264__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10814__A1 _10814_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08467_ _08470_/A _08470_/B vssd1 vssd1 vccd1 vccd1 _08467_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_64_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10814__B2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07418_ _10456_/S _10004_/S _09703_/B _07398_/B _11463_/A vssd1 vssd1 vccd1 vccd1
+ _07420_/B sky130_fd_sc_hd__o311a_4
XFILLER_0_80_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07691__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08398_ _08417_/A _08417_/B _08392_/X vssd1 vssd1 vccd1 vccd1 _08408_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_123_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07349_ reg1_val[20] _07634_/B _13082_/B vssd1 vssd1 vccd1 vccd1 _07349_/X sky130_fd_sc_hd__or3_1
X_10360_ _10360_/A _10360_/B vssd1 vssd1 vccd1 vccd1 _10363_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_33_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09019_ _09019_/A _09019_/B vssd1 vssd1 vccd1 vccd1 _10731_/C sky130_fd_sc_hd__xnor2_1
X_10291_ _10292_/A _10292_/B vssd1 vssd1 vccd1 vccd1 _10291_/X sky130_fd_sc_hd__and2_1
X_12030_ _12120_/B _12030_/B vssd1 vssd1 vccd1 vccd1 _12032_/C sky130_fd_sc_hd__and2_1
XANTENNA__07518__A _11281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold170 hold170/A vssd1 vssd1 vccd1 vccd1 hold170/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 hold181/A vssd1 vssd1 vccd1 vccd1 hold181/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 hold192/A vssd1 vssd1 vccd1 vccd1 hold192/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12932_ _12937_/C _12932_/B vssd1 vssd1 vccd1 vccd1 new_PC[19] sky130_fd_sc_hd__xnor2_4
XFILLER_0_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12863_ _12872_/A _12863_/B vssd1 vssd1 vccd1 vccd1 _12865_/C sky130_fd_sc_hd__nand2_1
X_11814_ _12092_/A _11814_/B vssd1 vssd1 vccd1 vccd1 _11816_/B sky130_fd_sc_hd__xnor2_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _09839_/A _09499_/Y _09860_/A _12783_/A _12793_/Y vssd1 vssd1 vccd1 vccd1
+ _12794_/X sky130_fd_sc_hd__o221a_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _11745_/A _11745_/B vssd1 vssd1 vccd1 vccd1 _11746_/B sky130_fd_sc_hd__xnor2_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12007__B1 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08084__A _10266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11676_ _11674_/X _11675_/X _07092_/D vssd1 vssd1 vccd1 vccd1 _11676_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10018__C1 _12760_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13415_ _07467_/B _13419_/A2 hold108/X vssd1 vssd1 vccd1 vccd1 _13689_/D sky130_fd_sc_hd__o21a_1
X_10627_ _10342_/A _10625_/Y _10626_/X _10624_/X vssd1 vssd1 vccd1 vccd1 dest_val[7]
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_70_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07029__A3 _12806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10119__A _10119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10033__A2 _12314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13346_ hold297/X _13506_/B2 _13506_/A2 hold193/X vssd1 vssd1 vccd1 vccd1 hold194/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10558_ _10415_/A _10415_/B _10398_/A vssd1 vssd1 vccd1 vccd1 _10569_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_106_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06788__A2 _13082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13277_ hold7/X hold285/A vssd1 vssd1 vccd1 vccd1 _13277_/X sky130_fd_sc_hd__and2b_1
X_10489_ _12093_/A _10489_/B vssd1 vssd1 vccd1 vccd1 _10497_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_121_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12228_ _12311_/B1 _12393_/C _13663_/Q vssd1 vssd1 vccd1 vccd1 _12230_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__13149__B _13193_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07737__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07737__B2 _08821_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12159_ _07201_/B _11793_/B _07152_/X _12158_/X vssd1 vssd1 vccd1 vccd1 _12159_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_75_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06986__B _07556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09370_ _07238_/X _12667_/A _10536_/A2 _07239_/Y vssd1 vssd1 vccd1 vccd1 _09371_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12797__A1 _09529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08321_ _08321_/A vssd1 vssd1 vccd1 vccd1 _08401_/A sky130_fd_sc_hd__inv_2
XFILLER_0_46_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08252_ _08252_/A _08252_/B vssd1 vssd1 vccd1 vccd1 _08347_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07673__B1 _08486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10272__A2 _10518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07203_ _07203_/A _07204_/B vssd1 vssd1 vccd1 vccd1 _07203_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_27_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08183_ _10266_/A _08183_/B vssd1 vssd1 vccd1 vccd1 _08186_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout125_A _07347_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07134_ instruction[29] instruction[22] _07135_/S vssd1 vssd1 vccd1 vccd1 reg2_idx[4]
+ sky130_fd_sc_hd__mux2_8
XANTENNA__07976__A1 _08806_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07976__B2 _08806_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07065_ reg1_val[25] _07223_/A vssd1 vssd1 vccd1 vccd1 _07079_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_100_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10980__B1 _10978_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13059__B _13059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07728__A1 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07728__B2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09553__A _12092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07967_ _08033_/A _08033_/B vssd1 vssd1 vccd1 vccd1 _07967_/X sky130_fd_sc_hd__and2_1
XANTENNA__06896__B _12990_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ hold245/A _12314_/A hold262/A vssd1 vssd1 vccd1 vccd1 _09706_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_4_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06918_ _11586_/A _06919_/B vssd1 vssd1 vccd1 vccd1 _06918_/X sky130_fd_sc_hd__and2_1
X_07898_ _07897_/B _07897_/C _07897_/A vssd1 vssd1 vccd1 vccd1 _07899_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__09350__B1 _10536_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09637_ _09340_/A _09340_/B _09341_/X vssd1 vssd1 vccd1 vccd1 _09642_/A sky130_fd_sc_hd__o21bai_2
XANTENNA__11307__B _11307_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06849_ _12778_/A _12452_/A _06849_/C _12382_/A vssd1 vssd1 vccd1 vccd1 _06850_/B
+ sky130_fd_sc_hd__or4_1
XANTENNA__12237__B1 _11688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09568_ _09568_/A _09568_/B vssd1 vssd1 vccd1 vccd1 _09613_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13434__C1 _13568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09102__B1 _07833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout38_A fanout39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08519_ _08520_/A _08520_/B vssd1 vssd1 vccd1 vccd1 _08519_/Y sky130_fd_sc_hd__nand2_1
X_09499_ _11576_/A _09497_/X _09498_/X vssd1 vssd1 vccd1 vccd1 _09499_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__10799__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12419__A _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11530_ _11530_/A _11530_/B vssd1 vssd1 vccd1 vccd1 _11531_/B sky130_fd_sc_hd__and2_1
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11461_ _11461_/A _11461_/B vssd1 vssd1 vccd1 vccd1 _11461_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__12853__S _12867_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13200_ _07257_/X _13598_/C hold43/X _13605_/A vssd1 vssd1 vccd1 vccd1 _13636_/D
+ sky130_fd_sc_hd__o211a_1
X_10412_ _10412_/A _10412_/B vssd1 vssd1 vccd1 vccd1 _10414_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__09728__A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11392_ _11392_/A _11392_/B vssd1 vssd1 vccd1 vccd1 _11430_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13131_ _13131_/A _13131_/B vssd1 vssd1 vccd1 vccd1 _13133_/A sky130_fd_sc_hd__nand2_2
X_10343_ _10480_/B _10342_/Y _12825_/S _10339_/X vssd1 vssd1 vccd1 vccd1 dest_val[5]
+ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__11696__C _11696_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07431__A3 _07435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07248__A _08951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13062_ _13062_/A _13062_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[15] sky130_fd_sc_hd__nor2_8
X_10274_ _10274_/A _10274_/B vssd1 vssd1 vccd1 vccd1 _10275_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12013_ _12016_/B _11916_/B _11924_/B _11925_/B _11925_/A vssd1 vssd1 vccd1 vccd1
+ _12025_/A sky130_fd_sc_hd__a32o_1
XANTENNA__07195__A2 _07213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08144__A1 _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08144__B2 wire122/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12915_ _12956_/A _12915_/B vssd1 vssd1 vccd1 vccd1 _12922_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12846_ _13015_/A curr_PC[7] _12867_/S vssd1 vssd1 vccd1 vccd1 _12848_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_75_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08807__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12777_ _10734_/A _07085_/Y _12740_/Y _12776_/Y vssd1 vssd1 vccd1 vccd1 _12778_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13440__A2 _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11728_ _11922_/A fanout8/X fanout3/X wire101/X vssd1 vssd1 vccd1 vccd1 _11729_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11659_ _11660_/A _11660_/B _11660_/C vssd1 vssd1 vccd1 vccd1 _11659_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_3_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09947__A2 _10536_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13329_ _13359_/A hold183/X vssd1 vssd1 vccd1 vccd1 hold184/A sky130_fd_sc_hd__and2_1
XFILLER_0_12_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07158__A _12982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11506__A2 _07597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08870_ _07175_/X _09910_/A1 _07420_/Y _08933_/B vssd1 vssd1 vccd1 vccd1 _08871_/B
+ sky130_fd_sc_hd__a22o_1
X_07821_ fanout24/X _10522_/A _09885_/B1 _08486_/B vssd1 vssd1 vccd1 vccd1 _07822_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09580__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09373__A _09373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10190__A1 _07363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07752_ _10049_/A2 _08486_/B _09885_/B1 fanout24/X vssd1 vssd1 vccd1 vccd1 _07753_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09332__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07683_ _07683_/A _07683_/B _07715_/A vssd1 vssd1 vccd1 vccd1 _07684_/B sky130_fd_sc_hd__and3_1
X_09422_ _09423_/A _09423_/B vssd1 vssd1 vccd1 vccd1 _09422_/X sky130_fd_sc_hd__and2_1
XFILLER_0_66_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10528__A1_N _07472_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09353_ _10095_/A _09353_/B vssd1 vssd1 vccd1 vccd1 _09357_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13431__A2 _13598_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08304_ _08873_/A2 _11047_/A fanout85/X _08891_/B vssd1 vssd1 vccd1 vccd1 _08305_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10245__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09284_ _11507_/A _09284_/B vssd1 vssd1 vccd1 vccd1 _09286_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08235_ _08235_/A _08235_/B vssd1 vssd1 vccd1 vccd1 _08236_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_90_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08166_ _08166_/A _08166_/B vssd1 vssd1 vccd1 vccd1 _08167_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_43_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07117_ _13142_/A _13141_/B vssd1 vssd1 vccd1 vccd1 _07117_/Y sky130_fd_sc_hd__nand2_1
X_08097_ _08168_/A _08168_/B _08094_/X vssd1 vssd1 vccd1 vccd1 _08109_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07048_ _11867_/B _11867_/C _07092_/B vssd1 vssd1 vccd1 vccd1 _11958_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_100_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08374__A1 _09501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08374__B2 _08271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ _08999_/A _08999_/B vssd1 vssd1 vccd1 vccd1 _09318_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_97_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10961_ _10841_/A _10841_/B _10839_/X vssd1 vssd1 vccd1 vccd1 _10968_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09874__A1 _12648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12700_ _12782_/C _12699_/Y _12782_/B vssd1 vssd1 vccd1 vccd1 _12700_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07885__B1 _08950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13680_ _13693_/CLK hold6/X vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08627__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10892_ _06966_/B _11587_/A2 _09520_/X _06963_/Y _10890_/X vssd1 vssd1 vccd1 vccd1
+ _10893_/B sky130_fd_sc_hd__o221a_1
XFILLER_0_78_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12631_ _12368_/X _12508_/X _12730_/B _12628_/Y _12630_/X vssd1 vssd1 vccd1 vccd1
+ _12632_/B sky130_fd_sc_hd__o311a_1
XANTENNA__08429__A2 wire122/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13422__A2 _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11053__A _11913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12562_ _12562_/A _12562_/B vssd1 vssd1 vccd1 vccd1 _12563_/B sky130_fd_sc_hd__and2_1
XFILLER_0_93_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11984__A2 _11793_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11513_ fanout54/X _07416_/X _07422_/Y _12268_/A vssd1 vssd1 vccd1 vccd1 _11514_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire122 wire122/A vssd1 vssd1 vccd1 vccd1 wire122/X sky130_fd_sc_hd__clkbuf_8
X_12493_ _12494_/A _12494_/B vssd1 vssd1 vccd1 vccd1 _12565_/B sky130_fd_sc_hd__and2_1
XFILLER_0_18_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13186__A1 _11997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11444_ _11445_/A _11445_/B vssd1 vssd1 vccd1 vccd1 _11551_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_34_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11375_ _07094_/C _09509_/X _11587_/A2 _06934_/B _11374_/X vssd1 vssd1 vccd1 vccd1
+ _11375_/X sky130_fd_sc_hd__o221a_1
X_13114_ _13121_/A _13114_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[26] sky130_fd_sc_hd__xnor2_4
X_10326_ _12314_/A _10325_/X hold294/A vssd1 vssd1 vccd1 vccd1 _10326_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_21_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _13045_/A _13045_/B _13045_/C vssd1 vssd1 vccd1 vccd1 _13046_/B sky130_fd_sc_hd__nand3_1
X_10257_ _10257_/A _10257_/B vssd1 vssd1 vccd1 vccd1 _10258_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_56_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10188_ hold283/A _12314_/A _10463_/C _12748_/B1 vssd1 vssd1 vccd1 vccd1 _10188_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12331__B _12764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08668__A2 _10049_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12829_ _12830_/A _12830_/B _12830_/C vssd1 vssd1 vccd1 vccd1 _12837_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_29_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11888__A1_N _12710_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08020_ _08018_/A _08018_/B _08019_/X vssd1 vssd1 vccd1 vccd1 _08030_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_21_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08272__A _09659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11188__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11410__B fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout7 fanout7/A vssd1 vssd1 vccd1 vccd1 fanout7/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_12_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09971_ _09789_/A _09789_/B _09787_/Y vssd1 vssd1 vccd1 vccd1 _09974_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_40_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08922_ _09371_/A _08922_/B vssd1 vssd1 vccd1 vccd1 _08931_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12152__A2 _09520_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08853_ _09371_/A _08853_/B vssd1 vssd1 vccd1 vccd1 _08887_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10163__A1 _10734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07804_ _10235_/A1 _11732_/A _10814_/A1 _10235_/B2 vssd1 vssd1 vccd1 vccd1 _07805_/B
+ sky130_fd_sc_hd__o22a_1
X_08784_ _08784_/A _08784_/B vssd1 vssd1 vccd1 vccd1 _08788_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_79_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07735_ _07300_/Y _10536_/B2 _11638_/A _08806_/A2 vssd1 vssd1 vccd1 vccd1 _07736_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11112__B1 _11342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07666_ _10507_/A _07666_/B vssd1 vssd1 vccd1 vccd1 _07749_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09405_ _09405_/A _09405_/B vssd1 vssd1 vccd1 vccd1 _09406_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13072__B _13129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10871__C1 _09507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07597_ _10787_/B _10787_/C vssd1 vssd1 vccd1 vccd1 _07597_/X sky130_fd_sc_hd__or2_4
X_09336_ _09337_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09336_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_63_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09267_ _11958_/A _12656_/A reg1_val[29] _13129_/A _13135_/A vssd1 vssd1 vccd1 vccd1
+ _12718_/B sky130_fd_sc_hd__a2111o_1
XANTENNA__08831__A2 _08873_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11601__A _12372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13168__A1 _13168_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08218_ _08290_/A _08290_/B _08290_/C vssd1 vssd1 vccd1 vccd1 _08291_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09198_ _09198_/A _09198_/B vssd1 vssd1 vccd1 vccd1 _09200_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11179__B1 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11718__A2 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08149_ _08173_/A vssd1 vssd1 vccd1 vccd1 _08225_/A sky130_fd_sc_hd__inv_2
XFILLER_0_120_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08595__A1 _08873_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08595__B2 _08891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11160_ _11161_/A _11161_/B _11161_/C vssd1 vssd1 vccd1 vccd1 _11162_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10111_ _10112_/A _10112_/B vssd1 vssd1 vccd1 vccd1 _10111_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11091_ _11091_/A _11091_/B vssd1 vssd1 vccd1 vccd1 _11092_/B sky130_fd_sc_hd__xnor2_1
X_10042_ _10041_/A _10041_/B _12825_/S vssd1 vssd1 vccd1 vccd1 _10042_/X sky130_fd_sc_hd__a21o_1
XANTENNA__11351__B1 _10866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
X_11993_ _11994_/A _11994_/B vssd1 vssd1 vccd1 vccd1 _12107_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12300__C1 _12578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13732_ _13735_/CLK _13732_/D vssd1 vssd1 vccd1 vccd1 hold249/A sky130_fd_sc_hd__dfxtp_1
X_10944_ _10944_/A _10944_/B vssd1 vssd1 vccd1 vccd1 _10952_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13663_ _13719_/CLK hold176/X vssd1 vssd1 vccd1 vccd1 _13663_/Q sky130_fd_sc_hd__dfxtp_1
X_10875_ _10873_/Y _10875_/B vssd1 vssd1 vccd1 vccd1 _10876_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_38_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10209__A2 _11423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12614_ _12614_/A _12764_/B _12614_/C vssd1 vssd1 vccd1 vccd1 _12675_/B sky130_fd_sc_hd__and3_1
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13594_ _13592_/X _13594_/B _13605_/A vssd1 vssd1 vccd1 vccd1 _13737_/D sky130_fd_sc_hd__and3b_1
XFILLER_0_93_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12545_ _07108_/D _12541_/X _12544_/X vssd1 vssd1 vccd1 vccd1 dest_val[26] sky130_fd_sc_hd__o21ai_4
XFILLER_0_81_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12476_ _12476_/A _12476_/B _12476_/C _12475_/X vssd1 vssd1 vccd1 vccd1 _12476_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_34_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_5 _06989_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ _11427_/A _11427_/B vssd1 vssd1 vccd1 vccd1 _11428_/B sky130_fd_sc_hd__or2_1
XFILLER_0_22_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11358_ reg1_val[13] curr_PC[13] vssd1 vssd1 vccd1 vccd1 _11360_/A sky130_fd_sc_hd__or2_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10309_ _07003_/B _10308_/X _10734_/A vssd1 vssd1 vccd1 vccd1 _10309_/Y sky130_fd_sc_hd__a21oi_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11884__C _12235_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11289_ _11288_/B _11288_/C _11288_/A vssd1 vssd1 vccd1 vccd1 _11290_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__12342__A _12417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08338__A1 _09671_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08338__B2 _08873_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13028_ reg1_val[10] _13029_/B vssd1 vssd1 vccd1 vccd1 _13030_/A sky130_fd_sc_hd__or2_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13157__B _13191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07561__A2 _08395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07520_ _07524_/A _11410_/A _11281_/A vssd1 vssd1 vccd1 vccd1 _07520_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07313__A2 _10536_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07171__A _08203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07451_ _10889_/A _07452_/B vssd1 vssd1 vccd1 vccd1 _07451_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_119_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07382_ _07641_/A _07641_/B vssd1 vssd1 vccd1 vccd1 _12551_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_17_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09121_ _09121_/A _09121_/B vssd1 vssd1 vccd1 vccd1 _09169_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09052_ _09052_/A _09052_/B vssd1 vssd1 vccd1 vccd1 _09055_/B sky130_fd_sc_hd__or2_1
X_08003_ _08006_/A _08006_/B vssd1 vssd1 vccd1 vccd1 _08003_/X sky130_fd_sc_hd__or2_1
XFILLER_0_115_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09954_ _09954_/A _09954_/B vssd1 vssd1 vccd1 vccd1 _09963_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_110_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12252__A _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09526__B1 _09521_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08905_ _09371_/A _08905_/B vssd1 vssd1 vccd1 vccd1 _08910_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ _07699_/B _07451_/X _09885_/B1 fanout35/X vssd1 vssd1 vccd1 vccd1 _09886_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _08836_/A _08836_/B vssd1 vssd1 vccd1 vccd1 _08847_/B sky130_fd_sc_hd__xnor2_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08767_ _08806_/A2 _07399_/Y _09910_/A1 _08806_/B1 vssd1 vssd1 vccd1 vccd1 _08768_/B
+ sky130_fd_sc_hd__a22o_1
X_07718_ _07718_/A _07718_/B vssd1 vssd1 vccd1 vccd1 _07842_/A sky130_fd_sc_hd__nand2_1
X_08698_ _08698_/A _08698_/B vssd1 vssd1 vccd1 vccd1 _08700_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_73_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10857__D _10981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07649_ _07649_/A _07649_/B vssd1 vssd1 vccd1 vccd1 _07650_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13389__A1 _09371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10660_ _11603_/A _10660_/B vssd1 vssd1 vccd1 vccd1 _10664_/A sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout20_A fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08905__A _09371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12597__C1 _12748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09319_ _09089_/A _09318_/Y _09317_/Y _09314_/Y vssd1 vssd1 vccd1 vccd1 _10579_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_118_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08265__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12061__A1 _07201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10591_ _12515_/S _10590_/Y _10588_/X vssd1 vssd1 vccd1 vccd1 _10592_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_106_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10072__B1 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12330_ _07415_/Y fanout7/X _12329_/Y _12421_/A vssd1 vssd1 vccd1 vccd1 _12411_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_23_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12261_ _12260_/A _12260_/B _12260_/C vssd1 vssd1 vccd1 vccd1 _12262_/B sky130_fd_sc_hd__a21o_1
X_11212_ _11092_/A _11092_/B _11090_/X vssd1 vssd1 vccd1 vccd1 _11213_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08640__A _10944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12192_ _12192_/A _12192_/B _12192_/C vssd1 vssd1 vccd1 vccd1 _12193_/B sky130_fd_sc_hd__or3_1
X_11143_ _10458_/S _10179_/X _09537_/B vssd1 vssd1 vccd1 vccd1 _11143_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07791__A2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09517__B1 _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11074_ _11281_/A _11074_/B vssd1 vssd1 vccd1 vccd1 _11076_/B sky130_fd_sc_hd__xnor2_1
X_10025_ _10734_/A _07014_/Y _07032_/X _10024_/Y vssd1 vssd1 vccd1 vccd1 _10026_/B
+ sky130_fd_sc_hd__a31oi_1
X_11976_ reg1_val[19] _11688_/B _09515_/Y _06884_/B vssd1 vssd1 vccd1 vccd1 _11980_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_86_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13715_ _13719_/CLK _13715_/D vssd1 vssd1 vccd1 vccd1 hold280/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11225__B _11342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10927_ _10927_/A _10927_/B vssd1 vssd1 vccd1 vccd1 _10929_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_86_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13646_ _13649_/CLK hold184/X vssd1 vssd1 vccd1 vccd1 hold182/A sky130_fd_sc_hd__dfxtp_1
X_10858_ _09654_/A _09654_/B _10298_/X _10857_/X vssd1 vssd1 vccd1 vccd1 _10858_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_27_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13577_ hold247/X _13584_/B _13576_/X _13599_/D vssd1 vssd1 vccd1 vccd1 hold248/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10789_ _10790_/B _10790_/C _11286_/A vssd1 vssd1 vccd1 vccd1 _10791_/B sky130_fd_sc_hd__a21o_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12528_ _12786_/B1 _12595_/B hold273/A vssd1 vssd1 vccd1 vccd1 _12528_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12056__B _12056_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12459_ reg1_val[25] curr_PC[25] vssd1 vssd1 vccd1 vccd1 _12460_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09756__B1 _10536_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11563__B1 _11866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07231__A1 _12982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10118__A1 fanout39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06951_ _07093_/A vssd1 vssd1 vccd1 vccd1 _11122_/A sky130_fd_sc_hd__inv_2
XANTENNA__06990__B1 _12782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10118__B2 _08118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09670_ _09452_/X _09478_/X _09703_/B vssd1 vssd1 vccd1 vccd1 _09670_/X sky130_fd_sc_hd__mux2_1
X_06882_ reg1_val[19] _07281_/A vssd1 vssd1 vccd1 vccd1 _06884_/A sky130_fd_sc_hd__and2b_1
XANTENNA__09381__A _09381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08621_ _08621_/A _08621_/B vssd1 vssd1 vccd1 vccd1 _08653_/A sky130_fd_sc_hd__nand2_1
X_08552_ _08552_/A _08552_/B vssd1 vssd1 vccd1 vccd1 _08555_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_89_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07503_ _07504_/A _07653_/A _07504_/C vssd1 vssd1 vccd1 vccd1 _07505_/A sky130_fd_sc_hd__a21oi_1
X_08483_ _08551_/A _08551_/B vssd1 vssd1 vccd1 vccd1 _08552_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_43_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout155_A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07434_ reg1_val[17] _07865_/B vssd1 vssd1 vccd1 vccd1 _07445_/A sky130_fd_sc_hd__or2_2
XFILLER_0_43_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07365_ _07476_/B _07186_/B _07363_/X _06995_/B vssd1 vssd1 vccd1 vccd1 _07367_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_128_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09104_ fanout39/X _10522_/A _09885_/B1 _08118_/B vssd1 vssd1 vccd1 vccd1 _09105_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11151__A _11151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10054__B1 _07477_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07296_ _07192_/A _07192_/B _07521_/A vssd1 vssd1 vccd1 vccd1 _07296_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09035_ _08788_/A _08788_/B _08976_/B vssd1 vssd1 vccd1 vccd1 _09035_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_4_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11003__C1 _12760_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06899__B _11793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09937_ _11281_/A _09937_/B vssd1 vssd1 vccd1 vccd1 _09938_/A sky130_fd_sc_hd__xnor2_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09868_ _07015_/Y _12793_/A2 _11586_/B vssd1 vssd1 vccd1 vccd1 _09868_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout68_A _10538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08819_ _08838_/A _08838_/B vssd1 vssd1 vccd1 vccd1 _08843_/B sky130_fd_sc_hd__nor2_1
X_09799_ _09797_/X _09799_/B vssd1 vssd1 vccd1 vccd1 _09800_/B sky130_fd_sc_hd__nand2b_1
X_11830_ _11830_/A _11830_/B vssd1 vssd1 vccd1 vccd1 _11832_/B sky130_fd_sc_hd__xnor2_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _11761_/A _11856_/A vssd1 vssd1 vccd1 vccd1 _11950_/A sky130_fd_sc_hd__nor2_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13500_ hold280/X _13499_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13500_/X sky130_fd_sc_hd__mux2_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _10565_/A _10565_/B _10563_/Y vssd1 vssd1 vccd1 vccd1 _10713_/B sky130_fd_sc_hd__a21oi_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _11693_/A2 _11878_/C hold231/A vssd1 vssd1 vccd1 vccd1 _11692_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13431_ _07412_/B _13598_/C hold131/X vssd1 vssd1 vccd1 vccd1 _13697_/D sky130_fd_sc_hd__o21a_1
X_10643_ _10643_/A _10643_/B vssd1 vssd1 vccd1 vccd1 _10644_/B sky130_fd_sc_hd__or2_1
XFILLER_0_125_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13362_ hold174/X _13542_/B2 _13555_/A2 _13663_/Q vssd1 vssd1 vccd1 vccd1 hold175/A
+ sky130_fd_sc_hd__a22o_1
X_10574_ _10575_/A _10575_/B vssd1 vssd1 vccd1 vccd1 _10574_/X sky130_fd_sc_hd__and2_1
XFILLER_0_106_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12313_ hold255/A _12313_/B vssd1 vssd1 vccd1 vccd1 _12390_/B sky130_fd_sc_hd__or2_1
X_13293_ _13493_/B _13494_/A _13261_/X vssd1 vssd1 vccd1 vccd1 _13499_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12337__A2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12244_ curr_PC[22] _12325_/C _12406_/B1 vssd1 vssd1 vccd1 vccd1 _12244_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12175_ fanout15/X _12667_/A _09145_/Y fanout31/X vssd1 vssd1 vccd1 vccd1 _12176_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10405__A _12092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07764__A2 _13149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08961__A1 _08951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11126_ _11126_/A curr_PC[11] vssd1 vssd1 vccd1 vccd1 _11126_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_101_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11057_ _11709_/A _11057_/B vssd1 vssd1 vccd1 vccd1 _11059_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10008_ _10601_/B _10007_/X _10176_/A vssd1 vssd1 vccd1 vccd1 _10008_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_64_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09269__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11959_ _07092_/B _11868_/X _06893_/B vssd1 vssd1 vccd1 vccd1 _11959_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_58_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13629_ _13725_/CLK _13629_/D vssd1 vssd1 vccd1 vccd1 hold134/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07150_ _13744_/A instruction[5] _12578_/A _09525_/C vssd1 vssd1 vccd1 vccd1 _10889_/B
+ sky130_fd_sc_hd__and4b_4
XFILLER_0_14_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07081_ _12578_/B _12578_/C _12581_/A vssd1 vssd1 vccd1 vccd1 _07082_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_89_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09729__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13525__B2 _13542_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10339__A1 _11866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13688__CLK _13701_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout106 _07557_/Y vssd1 vssd1 vccd1 vccd1 _08868_/B1 sky130_fd_sc_hd__buf_6
XANTENNA__07755__A2 _10522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout117 _11508_/A vssd1 vssd1 vccd1 vccd1 _11281_/A sky130_fd_sc_hd__clkbuf_16
Xfanout128 _07308_/X vssd1 vssd1 vccd1 vccd1 _08806_/A2 sky130_fd_sc_hd__clkbuf_8
X_07983_ fanout53/X _08907_/A fanout47/X _08328_/B2 vssd1 vssd1 vccd1 vccd1 _07984_/B
+ sky130_fd_sc_hd__o22a_1
Xfanout139 _12311_/B1 vssd1 vssd1 vccd1 vccd1 _11693_/A2 sky130_fd_sc_hd__buf_4
X_09722_ _10342_/A _09720_/X _09721_/Y _09719_/X vssd1 vssd1 vccd1 vccd1 dest_val[1]
+ sky130_fd_sc_hd__a31o_4
X_06934_ _11373_/A _06934_/B vssd1 vssd1 vccd1 vccd1 _07094_/C sky130_fd_sc_hd__nand2_1
XANTENNA__09823__B _09824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07624__A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ _09986_/A _09315_/X _10150_/A _09989_/C _09989_/A vssd1 vssd1 vccd1 vccd1
+ _09654_/B sky130_fd_sc_hd__o32a_1
X_06865_ _06886_/A _13005_/B vssd1 vssd1 vccd1 vccd1 _06865_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout272_A _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08180__A2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08604_ _08602_/Y _08642_/B _08592_/Y vssd1 vssd1 vccd1 vccd1 _08613_/B sky130_fd_sc_hd__o21a_1
XANTENNA__10050__A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09584_ _09585_/B _09585_/C _09948_/A vssd1 vssd1 vccd1 vccd1 _09586_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_49_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06796_ _06928_/B _13042_/B vssd1 vssd1 vccd1 vccd1 _06796_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_54_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08535_ _08606_/A _08606_/B _08531_/Y vssd1 vssd1 vccd1 vccd1 _08548_/B sky130_fd_sc_hd__o21a_1
XANTENNA__12264__A1 _12413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12264__B2 _12331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13361__A _13543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08466_ _08466_/A _08466_/B vssd1 vssd1 vccd1 vccd1 _08470_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_64_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10814__A2 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13080__B _13129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07417_ _12421_/A _12329_/A _07415_/Y vssd1 vssd1 vccd1 vccd1 _07417_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07691__A1 _08328_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07691__B2 _08907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08397_ _08397_/A _08397_/B vssd1 vssd1 vccd1 vccd1 _08417_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07348_ _07348_/A _07637_/B vssd1 vssd1 vccd1 vccd1 _07360_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_116_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07279_ _07309_/A _07476_/B vssd1 vssd1 vccd1 vccd1 _07281_/C sky130_fd_sc_hd__nor2_1
X_09018_ _09018_/A _09018_/B vssd1 vssd1 vccd1 vccd1 _10731_/B sky130_fd_sc_hd__and2_1
XFILLER_0_60_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12319__A2 _12793_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13516__B2 _13542_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10290_ _10290_/A _10290_/B vssd1 vssd1 vccd1 vccd1 _10292_/B sky130_fd_sc_hd__xnor2_2
Xhold160 hold160/A vssd1 vssd1 vccd1 vccd1 hold160/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10225__A _10225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold171 hold171/A vssd1 vssd1 vccd1 vccd1 hold171/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 hold182/A vssd1 vssd1 vccd1 vccd1 hold182/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 hold193/A vssd1 vssd1 vccd1 vccd1 hold193/X sky130_fd_sc_hd__dlygate4sd3_1
X_12931_ _12938_/A _12931_/B vssd1 vssd1 vccd1 vccd1 _12932_/B sky130_fd_sc_hd__nand2_2
X_12862_ _13025_/B _12862_/B vssd1 vssd1 vccd1 vccd1 _12863_/B sky130_fd_sc_hd__or2_1
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11813_ _12413_/A fanout15/X fanout31/X _12496_/A vssd1 vssd1 vccd1 vccd1 _11814_/B
+ sky130_fd_sc_hd__a22o_1
X_12793_ _12778_/A _12793_/A2 _12792_/X vssd1 vssd1 vccd1 vccd1 _12793_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _11743_/A _11743_/B _11745_/A vssd1 vssd1 vccd1 vccd1 _11744_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_56_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12007__A1 _07257_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11675_ _11958_/A _11675_/B _11675_/C vssd1 vssd1 vccd1 vccd1 _11675_/X sky130_fd_sc_hd__and3_1
XANTENNA__12007__B2 _12614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13414_ hold107/X _13416_/A2 _13420_/B1 hold22/X _13383_/A vssd1 vssd1 vccd1 vccd1
+ hold108/A sky130_fd_sc_hd__o221a_1
X_10626_ curr_PC[7] _10763_/C vssd1 vssd1 vccd1 vccd1 _10626_/X sky130_fd_sc_hd__or2_1
XFILLER_0_36_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13345_ _13459_/A hold236/X vssd1 vssd1 vccd1 vccd1 _13654_/D sky130_fd_sc_hd__and2_1
XANTENNA__11230__A2 _12372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10557_ _10557_/A _10557_/B vssd1 vssd1 vccd1 vccd1 _10571_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_59_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13276_ _13274_/X _13276_/B vssd1 vssd1 vccd1 vccd1 _13465_/A sky130_fd_sc_hd__nand2b_1
X_10488_ _07310_/Y fanout20/X fanout18/X fanout42/X vssd1 vssd1 vccd1 vccd1 _10489_/B
+ sky130_fd_sc_hd__o22a_2
XANTENNA__12715__C1 _12971_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12227_ hold174/A _12227_/B vssd1 vssd1 vccd1 vccd1 _12393_/C sky130_fd_sc_hd__or2_1
XANTENNA__07737__A2 _08821_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08934__A1 _09948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12158_ _11955_/A _12128_/X _12129_/Y _12132_/X _12157_/X vssd1 vssd1 vccd1 vccd1
+ _12158_/X sky130_fd_sc_hd__o311a_1
X_11109_ _10851_/X _10977_/A _10977_/B vssd1 vssd1 vccd1 vccd1 _11109_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_0_75_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_12_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13705_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12089_ fanout38/X fanout10/X fanout5/X fanout36/X vssd1 vssd1 vccd1 vccd1 _12090_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13165__B _13191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08320_ _11286_/A _08320_/B vssd1 vssd1 vccd1 vccd1 _08321_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08251_ _08251_/A _08251_/B vssd1 vssd1 vccd1 vccd1 _08252_/B sky130_fd_sc_hd__and2_1
XANTENNA__11413__B _11413_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07673__A1 _07451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08870__B1 _07420_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07673__B2 _09173_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07202_ _07213_/A _07212_/C _07521_/A vssd1 vssd1 vccd1 vccd1 _07204_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08182_ _09671_/S fanout21/X _08246_/B _08873_/B2 vssd1 vssd1 vccd1 vccd1 _08183_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07133_ instruction[28] instruction[21] _07135_/S vssd1 vssd1 vccd1 vccd1 reg2_idx[3]
+ sky130_fd_sc_hd__mux2_8
XFILLER_0_15_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12525__A _12525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07976__A2 _13174_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07064_ reg1_val[26] _07217_/A vssd1 vssd1 vccd1 vccd1 _12578_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10980__A1 _10628_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07338__B _13082_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07728__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07966_ _07966_/A _07966_/B vssd1 vssd1 vccd1 vccd1 _08033_/B sky130_fd_sc_hd__xnor2_2
X_09705_ hold17/A _12578_/A vssd1 vssd1 vccd1 vccd1 _09705_/X sky130_fd_sc_hd__and2_1
X_06917_ reg1_val[15] _07544_/A vssd1 vssd1 vccd1 vccd1 _06919_/B sky130_fd_sc_hd__nand2_1
X_07897_ _07897_/A _07897_/B _07897_/C vssd1 vssd1 vccd1 vccd1 _07899_/A sky130_fd_sc_hd__and3_1
XFILLER_0_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09350__A1 _07230_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09636_ _09410_/A _09410_/B _09409_/A vssd1 vssd1 vccd1 vccd1 _09646_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09350__B2 _12331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06848_ _12581_/A _12740_/A _12693_/A _06848_/D vssd1 vssd1 vccd1 vccd1 _06850_/A
+ sky130_fd_sc_hd__or4_1
X_09567_ _09567_/A _09567_/B vssd1 vssd1 vccd1 vccd1 _09568_/B sky130_fd_sc_hd__xor2_2
X_06779_ instruction[0] instruction[1] instruction[2] pred_val vssd1 vssd1 vccd1 vccd1
+ _06894_/B sky130_fd_sc_hd__o31a_1
XANTENNA__13434__B1 _13444_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09102__A1 _10225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09102__B2 _10349_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08518_ _08518_/A _08518_/B vssd1 vssd1 vccd1 vccd1 _08520_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08185__A _10263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09498_ _11472_/S _09466_/X _09451_/X _10603_/S vssd1 vssd1 vccd1 vccd1 _09498_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_93_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10799__A1 _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10799__B2 _07477_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11996__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08449_ _08449_/A _08449_/B vssd1 vssd1 vccd1 vccd1 _08506_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_93_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13198__C1 _13568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11460_ _11864_/A _11460_/B vssd1 vssd1 vccd1 vccd1 _11461_/B sky130_fd_sc_hd__and2_1
XFILLER_0_92_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10411_ _10224_/A _10223_/B _10221_/X vssd1 vssd1 vccd1 vccd1 _10412_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_61_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11391_ _11391_/A _11391_/B vssd1 vssd1 vccd1 vccd1 _11392_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13130_ reg1_val[30] _13136_/A vssd1 vssd1 vccd1 vccd1 _13131_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07529__A _09591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10342_ _10342_/A _10342_/B vssd1 vssd1 vccd1 vccd1 _10342_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_104_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13061_ _13061_/A _13061_/B _13061_/C vssd1 vssd1 vccd1 vccd1 _13062_/B sky130_fd_sc_hd__and3_2
XFILLER_0_103_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10273_ _10274_/A _10274_/B vssd1 vssd1 vccd1 vccd1 _10273_/Y sky130_fd_sc_hd__nand2_1
X_12012_ _12012_/A _12012_/B vssd1 vssd1 vccd1 vccd1 _12027_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10184__C1 _12533_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12170__A _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08144__A2 _07541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12914_ reg1_val[17] curr_PC[17] _12978_/S vssd1 vssd1 vccd1 vccd1 _12915_/B sky130_fd_sc_hd__mux2_2
XANTENNA__11684__C1 _12760_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12845_ _12851_/B _12845_/B vssd1 vssd1 vccd1 vccd1 new_PC[6] sky130_fd_sc_hd__and2_4
XFILLER_0_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11514__A _11514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12776_ _13129_/A _09254_/A _10734_/A vssd1 vssd1 vccd1 vccd1 _12776_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12329__B fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _11727_/A _11727_/B vssd1 vssd1 vccd1 vccd1 _11737_/B sky130_fd_sc_hd__or2_1
XFILLER_0_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08852__B1 _10225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07430__C _07435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11658_ _11758_/B _11658_/B vssd1 vssd1 vccd1 vccd1 _11660_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_4_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10609_ _07492_/A _10889_/B _07266_/X _12754_/C _10608_/Y vssd1 vssd1 vccd1 vccd1
+ _10609_/X sky130_fd_sc_hd__a221o_2
XFILLER_0_52_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11589_ _11583_/Y _11584_/X _11588_/X vssd1 vssd1 vccd1 vccd1 _11589_/X sky130_fd_sc_hd__o21a_1
XANTENNA__12400__B2 _12710_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13328_ hold238/A _13506_/B2 _13506_/A2 hold182/X vssd1 vssd1 vccd1 vccd1 hold183/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07158__B _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13259_ hold62/X hold280/X vssd1 vssd1 vccd1 vccd1 _13259_/X sky130_fd_sc_hd__and2b_1
XANTENNA__12999__B _13000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06997__B _07110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07820_ _07830_/A _07830_/B vssd1 vssd1 vccd1 vccd1 _07836_/A sky130_fd_sc_hd__or2_1
XANTENNA__09580__A1 _07238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09580__B2 _07239_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12080__A _12417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07591__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10190__A2 _11793_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07751_ _10266_/A _07751_/B vssd1 vssd1 vccd1 vccd1 _07757_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09332__A1 _10104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09332__B2 _09955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07682_ _07683_/B _07715_/A _07683_/A vssd1 vssd1 vccd1 vccd1 _07780_/A sky130_fd_sc_hd__a21oi_1
X_09421_ _09421_/A _09421_/B vssd1 vssd1 vccd1 vccd1 _09423_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07902__A _10078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09352_ fanout49/X _10235_/A1 _10235_/B2 fanout51/X vssd1 vssd1 vccd1 vccd1 _09353_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08303_ _08358_/A _08358_/B vssd1 vssd1 vccd1 vccd1 _08303_/Y sky130_fd_sc_hd__nor2_1
X_09283_ fanout28/X fanout85/X fanout82/X _08395_/B vssd1 vssd1 vccd1 vccd1 _09284_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout235_A _09429_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08234_ _08234_/A _08234_/B _08234_/C vssd1 vssd1 vccd1 vccd1 _08235_/B sky130_fd_sc_hd__or3_1
XFILLER_0_51_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08733__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08165_ _08234_/A _08234_/B _08234_/C vssd1 vssd1 vccd1 vccd1 _08235_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10402__B1 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07116_ _13141_/A _13142_/B vssd1 vssd1 vccd1 vccd1 _07118_/B sky130_fd_sc_hd__nor2_4
X_08096_ _08096_/A _08096_/B vssd1 vssd1 vccd1 vccd1 _08168_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07047_ _11772_/B _11772_/C _11774_/A vssd1 vssd1 vccd1 vccd1 _11867_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_30_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08374__A2 _07300_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08998_ _08035_/X _08998_/B vssd1 vssd1 vccd1 vccd1 _09094_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_76_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07949_ _07647_/A _07647_/B _07632_/Y vssd1 vssd1 vccd1 vccd1 _07951_/B sky130_fd_sc_hd__a21oi_2
X_10960_ _10832_/A _10832_/C _10832_/B vssd1 vssd1 vccd1 vccd1 _10970_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__08908__A _09659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09619_ _12094_/A _09619_/B vssd1 vssd1 vccd1 vccd1 _09627_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07885__A1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07885__B2 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10891_ _07095_/A _12793_/A2 _12754_/C _07294_/X vssd1 vssd1 vccd1 vccd1 _10891_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12630_ _12507_/Y _12629_/Y _12730_/B vssd1 vssd1 vccd1 vccd1 _12630_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_78_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12561_ _12562_/A _12562_/B vssd1 vssd1 vccd1 vccd1 _12625_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_38_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11512_ _11512_/A _11512_/B vssd1 vssd1 vccd1 vccd1 _11516_/A sky130_fd_sc_hd__xnor2_2
Xwire101 wire101/A vssd1 vssd1 vccd1 vccd1 wire101/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__11988__B _12164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12492_ _12565_/A _12492_/B vssd1 vssd1 vccd1 vccd1 _12494_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_18_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11443_ _11443_/A _11443_/B vssd1 vssd1 vccd1 vccd1 _11445_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13186__A2 _13194_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11197__A1 _07477_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07259__A _09950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11374_ _07523_/A _11793_/B _12657_/B1 reg1_val[13] _11373_/Y vssd1 vssd1 vccd1 vccd1
+ _11374_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_0_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13113_ _13136_/A _07378_/D _13112_/X vssd1 vssd1 vccd1 vccd1 _13114_/B sky130_fd_sc_hd__a21bo_2
X_10325_ hold283/A _10463_/C vssd1 vssd1 vccd1 vccd1 _10325_/X sky130_fd_sc_hd__or2_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ _13045_/A _13045_/B _13045_/C vssd1 vssd1 vccd1 vccd1 _13051_/B sky130_fd_sc_hd__a21o_1
X_10256_ _10257_/A _10257_/B vssd1 vssd1 vccd1 vccd1 _10256_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10187_ _12314_/A _10463_/C hold283/A vssd1 vssd1 vccd1 vccd1 _10187_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12828_ _12837_/A _12828_/B vssd1 vssd1 vccd1 vccd1 _12830_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_56_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _12759_/A1 _09692_/X _12749_/Y _12754_/X _12758_/X vssd1 vssd1 vccd1 vccd1
+ _12759_/X sky130_fd_sc_hd__a2111o_1
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06772__S _07135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08272__B _08272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11188__A1 _07526_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11188__B2 _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09250__B1 _12667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout8 fanout9/X vssd1 vssd1 vccd1 vccd1 fanout8/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_12_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10935__B2 _11076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09970_ _09738_/A _09738_/B _09739_/Y vssd1 vssd1 vccd1 vccd1 _09975_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_0_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12137__B1 _09507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08921_ _07238_/X _07399_/Y _09910_/A1 _07239_/Y vssd1 vssd1 vccd1 vccd1 _08922_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09384__A _10522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08852_ _07238_/X _10104_/A _10225_/A _07239_/Y vssd1 vssd1 vccd1 vccd1 _08853_/B
+ sky130_fd_sc_hd__a22o_1
X_07803_ _07807_/A _07807_/B vssd1 vssd1 vccd1 vccd1 _08021_/B sky130_fd_sc_hd__and2_1
X_08783_ _08789_/A _08789_/B _08763_/Y vssd1 vssd1 vccd1 vccd1 _08788_/A sky130_fd_sc_hd__a21o_1
XANTENNA__11138__B _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07335__C _13082_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07734_ _07744_/B _07744_/C _07744_/A vssd1 vssd1 vccd1 vccd1 _07747_/A sky130_fd_sc_hd__a21oi_1
X_07665_ fanout82/X fanout75/X _08704_/B fanout76/X vssd1 vssd1 vccd1 vccd1 _07666_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09404_ _09405_/A _09405_/B vssd1 vssd1 vccd1 vccd1 _09404_/Y sky130_fd_sc_hd__nor2_1
X_07596_ _10787_/B _10787_/C vssd1 vssd1 vccd1 vccd1 _12614_/A sky130_fd_sc_hd__nor2_8
X_09335_ _12092_/A _09335_/B vssd1 vssd1 vccd1 vccd1 _09337_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_118_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09266_ _11958_/A _12754_/A _13135_/A vssd1 vssd1 vccd1 vccd1 _09266_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_62_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08217_ _08256_/A _08217_/B vssd1 vssd1 vccd1 vccd1 _08290_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__13168__A2 _13194_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09197_ _09197_/A _09197_/B vssd1 vssd1 vccd1 vccd1 _09198_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11179__A1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11179__B2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08148_ _08172_/A _08172_/B vssd1 vssd1 vccd1 vccd1 _08173_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08595__A2 _10522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08079_ _08115_/A vssd1 vssd1 vccd1 vccd1 _08079_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_31_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10110_ _10110_/A _10110_/B vssd1 vssd1 vccd1 vccd1 _10112_/B sky130_fd_sc_hd__xnor2_4
XANTENNA_fanout98_A _10119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11090_ _10928_/Y _10932_/A _11091_/B vssd1 vssd1 vccd1 vccd1 _11090_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_101_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10041_ _10041_/A _10041_/B vssd1 vssd1 vccd1 vccd1 _10340_/C sky130_fd_sc_hd__nor2_2
XANTENNA__13340__A2 _13506_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold88/X vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ _07487_/Y fanout7/X _11991_/X _12094_/A vssd1 vssd1 vccd1 vccd1 _11994_/B
+ sky130_fd_sc_hd__a22o_1
X_10943_ _12557_/B fanout83/X fanout79/X _07597_/X vssd1 vssd1 vccd1 vccd1 _10944_/B
+ sky130_fd_sc_hd__o22a_1
X_13731_ _13731_/CLK _13731_/D vssd1 vssd1 vccd1 vccd1 hold273/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10874_ reg1_val[9] curr_PC[9] vssd1 vssd1 vccd1 vccd1 _10875_/B sky130_fd_sc_hd__nand2_1
X_13662_ _13717_/CLK _13662_/D vssd1 vssd1 vccd1 vccd1 hold174/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12613_ _12675_/A _12613_/B vssd1 vssd1 vccd1 vccd1 _12614_/C sky130_fd_sc_hd__and2b_1
X_13593_ hold191/X _13599_/D vssd1 vssd1 vccd1 vccd1 _13594_/B sky130_fd_sc_hd__or2_1
XFILLER_0_53_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12544_ _12971_/S _12544_/B _12546_/B vssd1 vssd1 vccd1 vccd1 _12544_/X sky130_fd_sc_hd__or3b_1
XANTENNA__08373__A _08951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12475_ _12475_/A _12475_/B _12475_/C _12475_/D vssd1 vssd1 vccd1 vccd1 _12475_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_123_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11426_ _11426_/A _11426_/B vssd1 vssd1 vccd1 vccd1 _11427_/B sky130_fd_sc_hd__and2_1
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_6 _07203_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11357_ _11356_/A _11356_/B _09507_/X vssd1 vssd1 vccd1 vccd1 _11357_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07794__B1 _08704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11590__A1 _12748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10308_ _07010_/B _10161_/X _07001_/Y vssd1 vssd1 vccd1 vccd1 _10308_/X sky130_fd_sc_hd__a21o_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11288_ _11288_/A _11288_/B _11288_/C vssd1 vssd1 vccd1 vccd1 _11290_/B sky130_fd_sc_hd__and3_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13027_ _13027_/A _13027_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[9] sky130_fd_sc_hd__xor2_4
XANTENNA__08338__A2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10239_ _10239_/A _10240_/B vssd1 vssd1 vccd1 vccd1 _10239_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_83_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06767__S _07135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07452__A _10889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13173__B _13191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07450_ _07449_/A _07186_/B _07186_/C _07476_/B vssd1 vssd1 vccd1 vccd1 _07452_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07381_ _07641_/A _07641_/B vssd1 vssd1 vccd1 vccd1 _07381_/X sky130_fd_sc_hd__and2_1
XFILLER_0_8_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09120_ _09121_/B _09121_/A vssd1 vssd1 vccd1 vccd1 _09120_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_29_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09471__A0 _11126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09051_ _08983_/A _09051_/B vssd1 vssd1 vccd1 vccd1 _09052_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08002_ _11286_/A _08002_/B vssd1 vssd1 vccd1 vccd1 _08006_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout100_A _07310_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09953_ _09953_/A _09953_/B vssd1 vssd1 vccd1 vccd1 _09954_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08904_ _07238_/X _09910_/A1 _07420_/Y _07239_/Y vssd1 vssd1 vccd1 vccd1 _08905_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13322__A2 _13463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10053__A _11731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ _09766_/A _09766_/B _09786_/B _09784_/Y vssd1 vssd1 vccd1 vccd1 _09898_/A
+ sky130_fd_sc_hd__a31oi_4
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ _08862_/A _08862_/B vssd1 vssd1 vccd1 vccd1 _08863_/A sky130_fd_sc_hd__nor2_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08766_ _08766_/A _08766_/B vssd1 vssd1 vccd1 vccd1 _08776_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07717_ _07717_/A _07717_/B vssd1 vssd1 vccd1 vccd1 _07718_/B sky130_fd_sc_hd__or2_1
XANTENNA__10199__S _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08697_ _08697_/A _08697_/B vssd1 vssd1 vccd1 vccd1 _08698_/B sky130_fd_sc_hd__nand2_1
X_07648_ _07649_/A _07649_/B vssd1 vssd1 vccd1 vccd1 _07648_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_95_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07579_ _09575_/A _07579_/B vssd1 vssd1 vccd1 vccd1 _07583_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09318_ _09318_/A _09318_/B _09318_/C _09825_/A vssd1 vssd1 vccd1 vccd1 _09318_/Y
+ sky130_fd_sc_hd__nor4_1
XFILLER_0_48_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08265__A1 _08873_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08193__A _11286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08265__B2 _08891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10590_ _10590_/A _10590_/B vssd1 vssd1 vccd1 vccd1 _10590_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12061__A2 _12799_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10072__A1 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09249_ _09249_/A _09249_/B vssd1 vssd1 vccd1 vccd1 _09262_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10072__B2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12260_ _12260_/A _12260_/B _12260_/C vssd1 vssd1 vccd1 vccd1 _12336_/B sky130_fd_sc_hd__nand3_1
XANTENNA__09214__B1 _09885_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11211_ _11211_/A _11211_/B vssd1 vssd1 vccd1 vccd1 _11213_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12191_ _12192_/A _12192_/B _12192_/C vssd1 vssd1 vccd1 vccd1 _12283_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07537__A _11076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11142_ _11134_/Y _11135_/X _11141_/X vssd1 vssd1 vccd1 vccd1 _11142_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09517__A1 _10866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11073_ fanout84/X _07597_/X _07891_/X _08580_/B vssd1 vssd1 vccd1 vccd1 _11074_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07528__B1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ _07015_/Y _09865_/B _07016_/Y _10734_/A vssd1 vssd1 vccd1 vccd1 _10024_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11975_ _11975_/A _11975_/B vssd1 vssd1 vccd1 vccd1 _11975_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13714_ _13719_/CLK _13714_/D vssd1 vssd1 vccd1 vccd1 hold253/A sky130_fd_sc_hd__dfxtp_1
X_10926_ _10924_/X _10926_/B vssd1 vssd1 vccd1 vccd1 _10927_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_58_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10857_ _10857_/A _10981_/A _10981_/B _10981_/C vssd1 vssd1 vccd1 vccd1 _10857_/X
+ sky130_fd_sc_hd__or4_1
X_13645_ _13649_/CLK _13645_/D vssd1 vssd1 vccd1 vccd1 hold238/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ _07892_/A _07892_/B _07546_/X vssd1 vssd1 vccd1 vccd1 _10790_/C sky130_fd_sc_hd__a21o_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13576_ hold249/A _13575_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13576_/X sky130_fd_sc_hd__mux2_1
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12527_ hold278/A _12527_/B vssd1 vssd1 vccd1 vccd1 _12595_/B sky130_fd_sc_hd__or2_1
XFILLER_0_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09927__A _11076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12458_ reg1_val[25] curr_PC[25] vssd1 vssd1 vccd1 vccd1 _12458_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_112_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11012__B1 _09520_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09756__A1 _12413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09756__B2 _12496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11409_ _11709_/A _11409_/B vssd1 vssd1 vccd1 vccd1 _11413_/A sky130_fd_sc_hd__xnor2_1
X_12389_ _10596_/Y _12388_/Y _12782_/B vssd1 vssd1 vccd1 vccd1 _12389_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07767__B1 _07833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07231__A2 _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06950_ _11138_/A _06950_/B vssd1 vssd1 vccd1 vccd1 _07093_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_94_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10118__A2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06881_ reg1_val[19] _07281_/A vssd1 vssd1 vccd1 vccd1 _07050_/A sky130_fd_sc_hd__and2_1
XFILLER_0_27_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08192__B1 _07545_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08620_ _08620_/A _08620_/B vssd1 vssd1 vccd1 vccd1 _08621_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09381__B _10522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_10_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08551_ _08551_/A _08551_/B vssd1 vssd1 vccd1 vccd1 _08552_/B sky130_fd_sc_hd__and2_1
X_07502_ _07502_/A _07502_/B vssd1 vssd1 vccd1 vccd1 _07504_/C sky130_fd_sc_hd__xor2_1
X_08482_ _10542_/A _08482_/B vssd1 vssd1 vccd1 vccd1 _08551_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07433_ _07486_/A _07486_/B vssd1 vssd1 vccd1 vccd1 _07433_/X sky130_fd_sc_hd__and2_1
XFILLER_0_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07364_ _07363_/B _07186_/B _07476_/B _06995_/B vssd1 vssd1 vccd1 vccd1 _07367_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09103_ _12421_/A _09103_/B vssd1 vssd1 vccd1 vccd1 _09110_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10054__A1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10054__B2 _07833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07295_ reg1_val[9] _07294_/X _07572_/S vssd1 vssd1 vccd1 vccd1 _07295_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09034_ _09034_/A _11233_/A _09034_/C _11117_/B vssd1 vssd1 vccd1 vccd1 _11460_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_115_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13078__B _13129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07222__A2 _07213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09936_ fanout40/X fanout83/X fanout79/X fanout56/X vssd1 vssd1 vccd1 vccd1 _09937_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_110_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06981__A1 _06936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09867_ _07097_/B _09864_/X _09865_/Y _09507_/X vssd1 vssd1 vccd1 vccd1 _09867_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08818_ _08818_/A _08818_/B vssd1 vssd1 vccd1 vccd1 _08838_/B sky130_fd_sc_hd__and2_1
XFILLER_0_99_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09798_ _09798_/A _09798_/B vssd1 vssd1 vccd1 vccd1 _09799_/B sky130_fd_sc_hd__or2_1
X_08749_ _09371_/A _08749_/B vssd1 vssd1 vccd1 vccd1 _08777_/A sky130_fd_sc_hd__xnor2_2
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _11550_/Y _11659_/Y _11661_/B vssd1 vssd1 vccd1 vccd1 _11760_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_67_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _10711_/A _10711_/B vssd1 vssd1 vccd1 vccd1 _10713_/A sky130_fd_sc_hd__xnor2_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11691_ hold195/A _11691_/B vssd1 vssd1 vccd1 vccd1 _11878_/C sky130_fd_sc_hd__or2_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11342__A _11342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10642_ _10643_/A _10643_/B vssd1 vssd1 vccd1 vccd1 _10780_/B sky130_fd_sc_hd__nand2_1
X_13430_ hold70/X _06744_/Y _13444_/B1 hold130/X _13430_/C1 vssd1 vssd1 vccd1 vccd1
+ hold131/A sky130_fd_sc_hd__o221a_1
XFILLER_0_125_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13361_ _13543_/A hold213/X vssd1 vssd1 vccd1 vccd1 _13662_/D sky130_fd_sc_hd__and2_1
XFILLER_0_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10573_ _10575_/A _10575_/B vssd1 vssd1 vccd1 vccd1 _10573_/X sky130_fd_sc_hd__or2_1
XFILLER_0_51_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12312_ hold229/A _12312_/B vssd1 vssd1 vccd1 vccd1 _12312_/Y sky130_fd_sc_hd__xnor2_1
X_13292_ _13488_/B _13489_/A _13263_/X vssd1 vssd1 vccd1 vccd1 _13494_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_51_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12243_ _12211_/Y _12212_/X _12214_/Y _10866_/B _12242_/Y vssd1 vssd1 vccd1 vccd1
+ _12243_/X sky130_fd_sc_hd__o221a_1
X_12174_ _12174_/A _12174_/B vssd1 vssd1 vccd1 vccd1 _12182_/A sky130_fd_sc_hd__nand2_1
X_11125_ _11126_/A curr_PC[11] vssd1 vssd1 vccd1 vccd1 _11125_/X sky130_fd_sc_hd__and2_1
X_11056_ fanout51/X fanout25/X fanout23/X _12557_/B vssd1 vssd1 vccd1 vccd1 _11057_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09910__A1 _09910_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10007_ _09685_/X _09687_/X _10007_/S vssd1 vssd1 vccd1 vccd1 _10007_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_98_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11958_ _11958_/A _11958_/B _11958_/C vssd1 vssd1 vccd1 vccd1 _11958_/X sky130_fd_sc_hd__and3_1
XFILLER_0_80_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11481__B1 _11587_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10909_ _10909_/A _10909_/B vssd1 vssd1 vccd1 vccd1 _10910_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11889_ _11887_/X _11889_/B _11889_/C _11889_/D vssd1 vssd1 vccd1 vccd1 _11889_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_117_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13628_ _13725_/CLK _13628_/D vssd1 vssd1 vccd1 vccd1 hold116/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13559_ hold269/X _13584_/B _13558_/X _13563_/B2 vssd1 vssd1 vccd1 vccd1 hold270/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11784__A1 _12710_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11784__B2 _12537_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07080_ _07079_/A _07079_/B _06849_/C vssd1 vssd1 vccd1 vccd1 _12578_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09729__A1 _10349_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09729__B2 _10225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13525__A2 _13555_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout118 _07460_/X vssd1 vssd1 vccd1 vccd1 _11508_/A sky130_fd_sc_hd__buf_8
X_07982_ _09948_/A _07982_/B vssd1 vssd1 vccd1 vccd1 _07989_/A sky130_fd_sc_hd__xnor2_2
Xfanout129 _07308_/X vssd1 vssd1 vccd1 vccd1 _10536_/A1 sky130_fd_sc_hd__clkbuf_4
X_09721_ curr_PC[0] curr_PC[1] vssd1 vssd1 vccd1 vccd1 _09721_/Y sky130_fd_sc_hd__nand2_1
X_06933_ reg1_val[13] _07522_/A vssd1 vssd1 vccd1 vccd1 _06934_/B sky130_fd_sc_hd__nand2_1
X_09652_ _09313_/A _09313_/B _09426_/A _09426_/B vssd1 vssd1 vccd1 vccd1 _09989_/C
+ sky130_fd_sc_hd__o2bb2a_1
X_06864_ instruction[30] _12981_/C vssd1 vssd1 vccd1 vccd1 _13005_/B sky130_fd_sc_hd__and2_4
X_08603_ _08645_/A _08603_/B vssd1 vssd1 vccd1 vccd1 _08642_/B sky130_fd_sc_hd__xnor2_2
X_09583_ _07892_/A _07892_/B _07200_/Y vssd1 vssd1 vccd1 vccd1 _09585_/C sky130_fd_sc_hd__a21o_1
X_06795_ instruction[37] _12981_/C vssd1 vssd1 vccd1 vccd1 _13042_/B sky130_fd_sc_hd__and2_4
XFILLER_0_89_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout265_A _13082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08534_ _08951_/A _08534_/B vssd1 vssd1 vccd1 vccd1 _08606_/B sky130_fd_sc_hd__xnor2_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12264__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08465_ _08463_/A _08463_/B _08464_/Y vssd1 vssd1 vccd1 vccd1 _08470_/A sky130_fd_sc_hd__o21ai_4
X_07416_ _07422_/A _07422_/B _12420_/A vssd1 vssd1 vccd1 vccd1 _07416_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08396_ _10263_/A _08457_/A _08457_/B vssd1 vssd1 vccd1 vccd1 _08417_/A sky130_fd_sc_hd__mux2_4
XANTENNA__07691__A2 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07347_ _08907_/B _08907_/C vssd1 vssd1 vccd1 vccd1 _07347_/X sky130_fd_sc_hd__or2_4
XFILLER_0_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07278_ _07193_/A _07193_/B _07190_/Y _07594_/B vssd1 vssd1 vccd1 vccd1 _07310_/B
+ sky130_fd_sc_hd__o31a_4
XFILLER_0_60_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09017_ _09017_/A _09017_/B vssd1 vssd1 vccd1 vccd1 _09018_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_103_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13516__A2 _13555_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold150 hold150/A vssd1 vssd1 vccd1 vccd1 hold150/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold161 hold161/A vssd1 vssd1 vccd1 vccd1 hold161/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10225__B _10518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold172 hold172/A vssd1 vssd1 vccd1 vccd1 hold172/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 hold183/A vssd1 vssd1 vccd1 vccd1 hold183/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 hold194/A vssd1 vssd1 vccd1 vccd1 hold194/X sky130_fd_sc_hd__dlygate4sd3_1
X_09919_ _09919_/A _09919_/B vssd1 vssd1 vccd1 vccd1 _09922_/B sky130_fd_sc_hd__xor2_1
X_12930_ _12938_/C _12930_/B vssd1 vssd1 vccd1 vccd1 _12937_/C sky130_fd_sc_hd__nand2_2
XANTENNA__07903__B1 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12867__S _12867_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12861_ _13025_/B _12862_/B vssd1 vssd1 vccd1 vccd1 _12872_/A sky130_fd_sc_hd__nand2_1
X_11812_ _12094_/A _11812_/B vssd1 vssd1 vccd1 vccd1 _11816_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ reg1_val[31] _07398_/B _09515_/Y _12790_/Y _12791_/X vssd1 vssd1 vccd1 vccd1
+ _12792_/X sky130_fd_sc_hd__a311o_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07550__A _11286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _11743_/A _11743_/B vssd1 vssd1 vccd1 vccd1 _11745_/B sky130_fd_sc_hd__nor2_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12168__A _12417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11072__A _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13204__A1 _12667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12007__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11674_ _12515_/S _11674_/B vssd1 vssd1 vccd1 vccd1 _11674_/X sky130_fd_sc_hd__and2_1
XFILLER_0_126_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10018__A1 _12525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13413_ _11281_/A _13419_/A2 hold137/X vssd1 vssd1 vccd1 vccd1 _13688_/D sky130_fd_sc_hd__o21a_1
X_10625_ curr_PC[7] _10763_/C vssd1 vssd1 vccd1 vccd1 _10625_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_107_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10556_ _10556_/A _10556_/B vssd1 vssd1 vccd1 vccd1 _10557_/B sky130_fd_sc_hd__nor2_2
X_13344_ hold214/X _13506_/B2 _13506_/A2 hold235/X vssd1 vssd1 vccd1 vccd1 hold236/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10487_ _10351_/A _10350_/B _10348_/X vssd1 vssd1 vccd1 vccd1 _10499_/A sky130_fd_sc_hd__a21o_2
X_13275_ hold264/X hold83/X vssd1 vssd1 vccd1 vccd1 _13276_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12226_ _12225_/A _12224_/X _12225_/Y _07137_/Y vssd1 vssd1 vccd1 vccd1 _12241_/A
+ sky130_fd_sc_hd__o211a_1
X_12157_ _12136_/Y _12137_/X _12144_/X _12156_/X vssd1 vssd1 vccd1 vccd1 _12157_/X
+ sky130_fd_sc_hd__o211a_1
X_11108_ _10578_/X _10579_/X _10581_/Y _11107_/Y vssd1 vssd1 vccd1 vccd1 _11113_/B
+ sky130_fd_sc_hd__a31o_1
X_12088_ _12088_/A _12088_/B vssd1 vssd1 vccd1 vccd1 _12099_/A sky130_fd_sc_hd__xor2_1
X_11039_ _11161_/A _11039_/B vssd1 vssd1 vccd1 vccd1 _11041_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_79_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09940__A _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13181__B _13191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12078__A _12666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08250_ _10263_/A _08250_/B vssd1 vssd1 vccd1 vccd1 _08347_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08870__A1 _07175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07673__A2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08870__B2 _08933_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07201_ _07201_/A _07201_/B vssd1 vssd1 vccd1 vccd1 _07212_/C sky130_fd_sc_hd__and2_2
XFILLER_0_7_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08181_ _09940_/A _08181_/B vssd1 vssd1 vccd1 vccd1 _08186_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12806__A _12806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07132_ instruction[27] instruction[20] _07135_/S vssd1 vssd1 vccd1 vccd1 reg2_idx[2]
+ sky130_fd_sc_hd__mux2_8
XFILLER_0_70_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06804__A _06886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07063_ reg1_val[27] _07251_/A vssd1 vssd1 vccd1 vccd1 _07082_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_23_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07965_ _07965_/A _07965_/B vssd1 vssd1 vccd1 vccd1 _08033_/A sky130_fd_sc_hd__and2_2
XANTENNA__08138__B1 _13172_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09704_ _07026_/A _09509_/X _09520_/X vssd1 vssd1 vccd1 vccd1 _09704_/X sky130_fd_sc_hd__o21a_1
X_06916_ reg1_val[15] _07544_/A vssd1 vssd1 vccd1 vccd1 _11586_/A sky130_fd_sc_hd__or2_1
X_07896_ _07895_/B _07895_/C _09949_/A vssd1 vssd1 vccd1 vccd1 _07897_/C sky130_fd_sc_hd__a21o_1
X_09635_ _09635_/A _09635_/B vssd1 vssd1 vccd1 vccd1 _09648_/A sky130_fd_sc_hd__xor2_4
XANTENNA__09350__A2 _10536_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11693__B1 _12533_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06847_ _06847_/A _06847_/B vssd1 vssd1 vccd1 vccd1 _12382_/A sky130_fd_sc_hd__nor2_2
X_09566_ _09567_/A _09567_/B vssd1 vssd1 vccd1 vccd1 _09566_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12237__A2 _12799_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06778_ reg2_val[31] _07110_/A vssd1 vssd1 vccd1 vccd1 _06778_/X sky130_fd_sc_hd__and2_1
XFILLER_0_77_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09102__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07370__A _10119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08517_ _08517_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08520_/A sky130_fd_sc_hd__nor2_1
XANTENNA__13091__B _13129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09497_ _09481_/X _09496_/X _11575_/S vssd1 vssd1 vccd1 vccd1 _09497_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10799__A2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11996__A1 _12189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10000__S _10004_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11996__B2 _07198_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08448_ _08448_/A _08448_/B vssd1 vssd1 vccd1 vccd1 _08449_/B sky130_fd_sc_hd__or2_1
XFILLER_0_108_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08379_ _08379_/A _08379_/B vssd1 vssd1 vccd1 vccd1 _08453_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_46_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10410_ _10410_/A _10410_/B vssd1 vssd1 vccd1 vccd1 _10412_/A sky130_fd_sc_hd__xor2_4
X_11390_ _11388_/A _11388_/B _11391_/B vssd1 vssd1 vccd1 vccd1 _11390_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_33_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10341_ curr_PC[4] _10340_/C curr_PC[5] vssd1 vssd1 vccd1 vccd1 _10342_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_104_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10236__A _10236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13060_ _13061_/A _13061_/B _13061_/C vssd1 vssd1 vccd1 vccd1 _13062_/A sky130_fd_sc_hd__a21oi_4
X_10272_ _10104_/A _10518_/A _10110_/B _10108_/X vssd1 vssd1 vccd1 vccd1 _10274_/B
+ sky130_fd_sc_hd__a31o_1
X_12011_ _12011_/A _12011_/B vssd1 vssd1 vccd1 vccd1 _12012_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13370__B1 _13584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09877__B1 _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12913_ _12922_/A _12913_/B vssd1 vssd1 vccd1 vccd1 new_PC[16] sky130_fd_sc_hd__and2_4
X_12844_ _12844_/A _12844_/B _12844_/C vssd1 vssd1 vccd1 vccd1 _12845_/B sky130_fd_sc_hd__nand3_1
XANTENNA__13425__A1 _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _12763_/Y _12771_/Y _12773_/X _12774_/X _09429_/X vssd1 vssd1 vccd1 vccd1
+ _12775_/Y sky130_fd_sc_hd__a311oi_4
XANTENNA__11987__A1 _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _11727_/A _11727_/B vssd1 vssd1 vccd1 vccd1 _11737_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08852__A1 _07238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08852__B2 _07239_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11657_ _11657_/A _11657_/B vssd1 vssd1 vccd1 vccd1 _11658_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_36_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10608_ reg1_val[7] _11688_/B vssd1 vssd1 vccd1 vccd1 _10608_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_4_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11588_ _07094_/A _09509_/X _11585_/Y _11587_/X vssd1 vssd1 vccd1 vccd1 _11588_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13327_ _13459_/A hold239/X vssd1 vssd1 vccd1 vccd1 _13645_/D sky130_fd_sc_hd__and2_1
X_10539_ _07892_/A _07892_/B _07577_/X vssd1 vssd1 vccd1 vccd1 _10541_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_24_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13258_ hold291/A hold51/X vssd1 vssd1 vccd1 vccd1 _13503_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_122_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12209_ _12035_/A _11861_/B _12035_/B _12368_/B _12208_/X vssd1 vssd1 vccd1 vccd1
+ _12210_/B sky130_fd_sc_hd__o41a_2
XFILLER_0_110_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13189_ hold48/X _13191_/B vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__or2_1
XANTENNA__09580__A2 _10536_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07591__A1 _08821_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07591__B2 _08821_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07750_ _08866_/A2 fanout21/X _08246_/B _07366_/X vssd1 vssd1 vccd1 vccd1 _07751_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09868__B1 _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09332__A2 _07643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07681_ _07714_/A _07714_/B vssd1 vssd1 vccd1 vccd1 _07715_/A sky130_fd_sc_hd__or2_1
XANTENNA__10478__B2 _11866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09420_ _09421_/B _09421_/A vssd1 vssd1 vccd1 vccd1 _09420_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__11705__A _11913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07190__A _11793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09351_ _10078_/A _09351_/B vssd1 vssd1 vccd1 vccd1 _09359_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08302_ _08302_/A _08302_/B vssd1 vssd1 vccd1 vccd1 _08358_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09282_ _10266_/A _09282_/B vssd1 vssd1 vccd1 vccd1 _09286_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08233_ _08297_/A _08297_/B vssd1 vssd1 vccd1 vccd1 _08236_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_74_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout130_A _07285_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10034__A2_N _12235_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08164_ _08164_/A _08164_/B vssd1 vssd1 vccd1 vccd1 _08234_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_15_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10402__A1 _07299_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07115_ _07123_/B _09524_/B vssd1 vssd1 vccd1 vccd1 _13141_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_43_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08095_ _08095_/A _08095_/B vssd1 vssd1 vccd1 vccd1 _08168_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10402__B2 _10814_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07046_ _11675_/B _11675_/C _07092_/D vssd1 vssd1 vccd1 vccd1 _11772_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13352__B1 _13506_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11902__A1 _12557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07031__B1 _09703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11902__B2 _12557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13086__B _13129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ _08997_/A _08997_/B vssd1 vssd1 vccd1 vccd1 _09318_/B sky130_fd_sc_hd__xnor2_4
X_07948_ _07948_/A _07948_/B vssd1 vssd1 vccd1 vccd1 _07951_/A sky130_fd_sc_hd__or2_2
XANTENNA__09859__B1 _09529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07879_ _09604_/A _07643_/B fanout13/X _09161_/A vssd1 vssd1 vccd1 vccd1 _07880_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09618_ fanout85/X fanout21/X _08246_/B _07522_/Y vssd1 vssd1 vccd1 vccd1 _09619_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07885__A2 _08866_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08196__A _09948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10890_ reg1_val[9] _11688_/B _10889_/Y _12327_/A vssd1 vssd1 vccd1 vccd1 _10890_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout43_A fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09549_ _10050_/A _09549_/B vssd1 vssd1 vccd1 vccd1 _09557_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12560_ _12560_/A _12560_/B vssd1 vssd1 vccd1 vccd1 _12562_/B sky130_fd_sc_hd__xor2_1
XANTENNA__12091__B1 _12667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08924__A _09659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11511_ _12557_/A fanout20/X fanout18/X _12557_/B vssd1 vssd1 vccd1 vccd1 _11512_/B
+ sky130_fd_sc_hd__o22a_1
X_12491_ _12491_/A _12491_/B _12491_/C vssd1 vssd1 vccd1 vccd1 _12492_/B sky130_fd_sc_hd__and3_1
X_11442_ _11443_/B _11443_/A vssd1 vssd1 vccd1 vccd1 _11442_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_123_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08598__B1 _07556_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11197__A2 _11802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11373_ _11373_/A _11586_/B vssd1 vssd1 vccd1 vccd1 _11373_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_33_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13112_ _13112_/A _13112_/B vssd1 vssd1 vccd1 vccd1 _13112_/X sky130_fd_sc_hd__or2_1
X_10324_ _06994_/A _12793_/A2 _11586_/B vssd1 vssd1 vccd1 vccd1 _10324_/Y sky130_fd_sc_hd__a21oi_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13043_ _13043_/A _13051_/A vssd1 vssd1 vccd1 vccd1 _13045_/C sky130_fd_sc_hd__nand2_1
X_10255_ _10255_/A _10255_/B vssd1 vssd1 vccd1 vccd1 _10257_/B sky130_fd_sc_hd__xor2_1
XANTENNA__10157__B1 _10730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07275__A _10095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10186_ hold264/A hold285/A hold262/A hold245/A vssd1 vssd1 vccd1 vccd1 _10463_/C
+ sky130_fd_sc_hd__or4_2
XFILLER_0_100_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout290 reg1_val[11] vssd1 vssd1 vccd1 vccd1 _11126_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08522__B1 _07545_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_15_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12827_ _13000_/B _12827_/B vssd1 vssd1 vccd1 vccd1 _12828_/B sky130_fd_sc_hd__or2_1
XFILLER_0_8_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12758_ _12740_/A _12793_/A2 _09716_/Y _09504_/Y _12757_/X vssd1 vssd1 vccd1 vccd1
+ _12758_/X sky130_fd_sc_hd__a221o_1
XANTENNA__08834__A _10078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11709_ _11709_/A _11709_/B vssd1 vssd1 vccd1 vccd1 _11710_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12689_ _12733_/C _12688_/X _10730_/B vssd1 vssd1 vccd1 vccd1 _12689_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08589__B1 _07477_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11188__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09250__A1 _07238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09250__B2 _07239_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout9 fanout9/A vssd1 vssd1 vccd1 vccd1 fanout9/X sky130_fd_sc_hd__buf_6
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10935__A2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13334__B1 _13506_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08920_ _08920_/A _08920_/B _08920_/C vssd1 vssd1 vccd1 vccd1 _08929_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_110_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08851_ _08857_/A _08857_/B vssd1 vssd1 vccd1 vccd1 _08851_/Y sky130_fd_sc_hd__nand2_1
X_07802_ _10078_/A _07802_/B vssd1 vssd1 vccd1 vccd1 _07807_/B sky130_fd_sc_hd__xor2_1
X_08782_ _08755_/B _08765_/Y _08776_/B _08781_/X vssd1 vssd1 vccd1 vccd1 _08789_/B
+ sky130_fd_sc_hd__a31o_1
X_07733_ _07733_/A _07811_/B vssd1 vssd1 vccd1 vccd1 _07744_/C sky130_fd_sc_hd__or2_1
X_07664_ _07667_/A _07667_/B vssd1 vssd1 vccd1 vccd1 _07668_/A sky130_fd_sc_hd__and2_1
X_09403_ _09276_/A _09276_/B _09274_/Y vssd1 vssd1 vccd1 vccd1 _09405_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07595_ _07595_/A _07595_/B vssd1 vssd1 vccd1 vccd1 _10787_/C sky130_fd_sc_hd__nor2_8
XFILLER_0_1_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09334_ fanout14/X _10374_/B2 _10637_/A _07833_/B vssd1 vssd1 vccd1 vccd1 _09335_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12073__B1 _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11977__A2_N _09520_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06827__B1 _07110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09265_ _11958_/A _12754_/A _13135_/A vssd1 vssd1 vccd1 vccd1 _09265_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08216_ _08258_/A _08216_/B vssd1 vssd1 vccd1 vccd1 _08290_/B sky130_fd_sc_hd__nand2_1
X_09196_ _09197_/B _09197_/A vssd1 vssd1 vccd1 vccd1 _09196_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_105_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11179__A2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08147_ _09591_/A _08147_/B vssd1 vssd1 vccd1 vccd1 _08172_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10387__B1 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09575__A _09575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08078_ _09591_/A _08078_/B vssd1 vssd1 vccd1 vccd1 _08115_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07029_ _06928_/A _06928_/B _12806_/A _07027_/X vssd1 vssd1 vccd1 vccd1 _07029_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10040_ _09992_/Y _09993_/X _10039_/X vssd1 vssd1 vccd1 vccd1 _10040_/Y sky130_fd_sc_hd__o21bai_2
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08919__A _09948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ _11991_/A fanout5/X vssd1 vssd1 vccd1 vccd1 _11991_/X sky130_fd_sc_hd__or2_1
XFILLER_0_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13730_ _13731_/CLK _13730_/D vssd1 vssd1 vccd1 vccd1 hold278/A sky130_fd_sc_hd__dfxtp_1
X_10942_ _10811_/A _10811_/B _10812_/Y vssd1 vssd1 vccd1 vccd1 _10958_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_98_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13661_ _13717_/CLK hold179/X vssd1 vssd1 vccd1 vccd1 hold212/A sky130_fd_sc_hd__dfxtp_1
X_10873_ reg1_val[9] curr_PC[9] vssd1 vssd1 vccd1 vccd1 _10873_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_39_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ _12612_/A _12612_/B vssd1 vssd1 vccd1 vccd1 _12613_/B sky130_fd_sc_hd__or2_1
X_13592_ hold191/X _13599_/D _13207_/B vssd1 vssd1 vccd1 vccd1 _13592_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_66_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12543_ curr_PC[26] _12543_/B vssd1 vssd1 vccd1 vccd1 _12546_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11811__B1 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12176__A _12420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12474_ _07386_/Y _12754_/C _12473_/X vssd1 vssd1 vccd1 vccd1 _12475_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11425_ _11426_/A _11426_/B vssd1 vssd1 vccd1 vccd1 _11427_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_124_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12904__A _13059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_7 instruction[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07243__B1 _08950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11356_ _11356_/A _11356_/B vssd1 vssd1 vccd1 vccd1 _11356_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_104_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07794__A1 _11047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07794__B2 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10307_ _11864_/A _10306_/B _10306_/C vssd1 vssd1 vccd1 vccd1 _10307_/X sky130_fd_sc_hd__a21o_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11287_ _11286_/B _11286_/C _11286_/A vssd1 vssd1 vccd1 vccd1 _11288_/C sky130_fd_sc_hd__a21o_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13026_ _13031_/B _13033_/A vssd1 vssd1 vccd1 vccd1 _13027_/B sky130_fd_sc_hd__nand2_2
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10238_ _10537_/A _10238_/B vssd1 vssd1 vccd1 vccd1 _10240_/B sky130_fd_sc_hd__xnor2_1
X_10169_ _10167_/Y _10169_/B vssd1 vssd1 vccd1 vccd1 _10170_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_89_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07380_ _12598_/A _12598_/B _07865_/B vssd1 vssd1 vccd1 vccd1 _07641_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_45_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09050_ _09047_/A _09047_/B _09049_/Y _09048_/B _11562_/B vssd1 vssd1 vccd1 vccd1
+ _11864_/B sky130_fd_sc_hd__o2111ai_4
X_08001_ _09173_/B2 fanout75/X _08704_/B _11047_/A vssd1 vssd1 vccd1 vccd1 _08002_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09952_ _09953_/A _09953_/B vssd1 vssd1 vccd1 vccd1 _09952_/X sky130_fd_sc_hd__or2_1
X_08903_ _08911_/B _08911_/A vssd1 vssd1 vccd1 vccd1 _08903_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_110_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09883_ _09817_/A _09817_/B _09818_/Y vssd1 vssd1 vccd1 vccd1 _09982_/A sky130_fd_sc_hd__a21bo_2
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08734__B1 _08868_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout295_A _12578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08834_ _10078_/A _08834_/B vssd1 vssd1 vccd1 vccd1 _08862_/B sky130_fd_sc_hd__xnor2_2
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07643__A _09161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08765_ _08766_/A _08766_/B vssd1 vssd1 vccd1 vccd1 _08765_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11165__A _12092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07716_ _07719_/A _07719_/B vssd1 vssd1 vccd1 vccd1 _07716_/X sky130_fd_sc_hd__or2_1
X_08696_ _08724_/A _08724_/B vssd1 vssd1 vccd1 vccd1 _09051_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_67_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07647_ _07647_/A _07647_/B vssd1 vssd1 vccd1 vccd1 _07649_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07578_ fanout70/X fanout68/X fanout66/X _11732_/A vssd1 vssd1 vccd1 vccd1 _07579_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09317_ _08105_/Y _08998_/B _09825_/A _08035_/X _09318_/A vssd1 vssd1 vccd1 vccd1
+ _09317_/Y sky130_fd_sc_hd__a2111oi_2
XFILLER_0_118_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08265__A2 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11075__A_N _11076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09248_ _09248_/A _09248_/B vssd1 vssd1 vccd1 vccd1 _09249_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10072__A2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09214__A1 _08118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09179_ _09179_/A _09179_/B _09179_/C vssd1 vssd1 vccd1 vccd1 _09180_/B sky130_fd_sc_hd__and3_1
XFILLER_0_16_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09214__B2 fanout39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07225__B1 _08907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11210_ _11210_/A _11210_/B vssd1 vssd1 vccd1 vccd1 _11211_/B sky130_fd_sc_hd__nor2_1
X_12190_ _12190_/A _12190_/B vssd1 vssd1 vccd1 vccd1 _12192_/C sky130_fd_sc_hd__xnor2_1
X_11141_ _07531_/Y _12598_/C _12796_/A1 _11137_/Y _11140_/X vssd1 vssd1 vccd1 vccd1
+ _11141_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09517__A2 _11587_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11072_ _11072_/A _11072_/B vssd1 vssd1 vccd1 vccd1 _11078_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07528__A1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07528__B2 _11423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10023_ _12537_/B2 _10010_/X _10022_/Y _12759_/A1 vssd1 vssd1 vccd1 vccd1 _10023_/X
+ sky130_fd_sc_hd__a22o_1
X_11974_ _13660_/Q _12311_/B1 _12148_/C _12533_/B1 vssd1 vssd1 vccd1 vccd1 _11975_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_98_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13713_ _13725_/CLK _13713_/D vssd1 vssd1 vccd1 vccd1 hold295/A sky130_fd_sc_hd__dfxtp_1
X_10925_ _10925_/A _10925_/B vssd1 vssd1 vccd1 vccd1 _10926_/B sky130_fd_sc_hd__or2_1
XFILLER_0_58_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11803__A _11920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13644_ _13649_/CLK hold228/X vssd1 vssd1 vccd1 vccd1 hold226/A sky130_fd_sc_hd__dfxtp_1
X_10856_ _10580_/Y _11107_/A _10854_/Y vssd1 vssd1 vccd1 vccd1 _10856_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13575_ _13579_/C _13575_/B vssd1 vssd1 vccd1 vccd1 _13575_/Y sky130_fd_sc_hd__nor2_1
X_10787_ _10787_/A _10787_/B _10787_/C vssd1 vssd1 vccd1 vccd1 _10790_/B sky130_fd_sc_hd__or3_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12526_ _12525_/A _12524_/Y _12525_/Y _09529_/B vssd1 vssd1 vccd1 vccd1 _12526_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11260__B2 _12710_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12457_ _12388_/A _12385_/Y _12387_/B vssd1 vssd1 vccd1 vccd1 _12461_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_112_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09756__A2 _10536_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11408_ fanout25/X _07891_/X _09146_/Y fanout23/X vssd1 vssd1 vccd1 vccd1 _11409_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_112_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12388_ _12388_/A _12388_/B vssd1 vssd1 vccd1 vccd1 _12388_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__07767__A1 _09161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07767__B2 _09604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12760__A1 _12760_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11339_ _11340_/A _11340_/B _11340_/C vssd1 vssd1 vccd1 vccd1 _11339_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10771__B1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06990__A2 _07110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13009_ reg1_val[6] _13010_/B vssd1 vssd1 vccd1 vccd1 _13009_/Y sky130_fd_sc_hd__nor2_1
X_06880_ reg2_val[19] _06873_/B1 _06906_/B1 _06879_/Y vssd1 vssd1 vccd1 vccd1 _07281_/A
+ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__08192__A1 _07492_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08192__B2 _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08550_ _08560_/B _08560_/A vssd1 vssd1 vccd1 vccd1 _08562_/A sky130_fd_sc_hd__nand2b_1
X_07501_ _07502_/B vssd1 vssd1 vccd1 vccd1 _07501_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08481_ _08873_/A2 _10049_/A2 _09173_/B2 _08891_/B vssd1 vssd1 vccd1 vccd1 _08482_/B
+ sky130_fd_sc_hd__o22a_1
X_07432_ _07337_/Y _07431_/Y _07637_/B vssd1 vssd1 vccd1 vccd1 _07486_/B sky130_fd_sc_hd__a21o_1
XANTENNA__06807__A _13129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07363_ _12515_/S _07363_/B _07398_/B vssd1 vssd1 vccd1 vccd1 _07363_/X sky130_fd_sc_hd__or3b_1
X_09102_ _10225_/A fanout14/X _07833_/B _10349_/A1 vssd1 vssd1 vccd1 vccd1 _09103_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10054__A2 _07472_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07294_ reg1_val[9] _10750_/A vssd1 vssd1 vccd1 vccd1 _07294_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_127_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09033_ _09033_/A _09033_/B vssd1 vssd1 vccd1 vccd1 _09034_/C sky130_fd_sc_hd__xor2_2
XFILLER_0_60_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout210_A _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12544__A _12971_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11003__A1 _12525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08955__B1 _13147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07357__B _07535_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09935_ _09935_/A _09935_/B vssd1 vssd1 vccd1 vccd1 _09954_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08707__B1 _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11306__A2 _11307_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06981__A2 _06928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09866_ _09864_/X _09865_/Y _07097_/B vssd1 vssd1 vccd1 vccd1 _09866_/Y sky130_fd_sc_hd__a21oi_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08817_ _09671_/S _08778_/B _08778_/C vssd1 vssd1 vccd1 vccd1 _08818_/B sky130_fd_sc_hd__o21ai_1
X_09797_ _09798_/A _09798_/B vssd1 vssd1 vccd1 vccd1 _09797_/X sky130_fd_sc_hd__and2_1
XFILLER_0_84_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08748_ _07238_/X _07492_/Y _10637_/A _07239_/Y vssd1 vssd1 vccd1 vccd1 _08749_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _08690_/A _08690_/B vssd1 vssd1 vccd1 vccd1 _08679_/X sky130_fd_sc_hd__and2_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _10710_/A _10710_/B vssd1 vssd1 vccd1 vccd1 _10711_/B sky130_fd_sc_hd__xor2_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _07092_/D _12709_/A2 _12754_/C _07462_/Y _11689_/X vssd1 vssd1 vccd1 vccd1
+ _11696_/C sky130_fd_sc_hd__a221o_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10641_ _10641_/A _10641_/B vssd1 vssd1 vccd1 vccd1 _10643_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11342__B _11452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10239__A _10239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13360_ hold177/X _13463_/B2 _13450_/B hold174/X vssd1 vssd1 vccd1 vccd1 hold213/A
+ sky130_fd_sc_hd__a22o_1
X_10572_ _10572_/A _10572_/B vssd1 vssd1 vccd1 vccd1 _10575_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__08932__A _09703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12311_ _13663_/Q _12393_/C _12311_/B1 vssd1 vssd1 vccd1 vccd1 _12312_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13291_ _13483_/B _13484_/A _13265_/X vssd1 vssd1 vccd1 vccd1 _13489_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_16_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12242_ _12218_/Y _12219_/X _12241_/X vssd1 vssd1 vccd1 vccd1 _12242_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12173_ _12173_/A _12173_/B _12173_/C vssd1 vssd1 vccd1 vccd1 _12174_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_31_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11124_ _11126_/A curr_PC[11] vssd1 vssd1 vccd1 vccd1 _11124_/X sky130_fd_sc_hd__or2_1
XFILLER_0_101_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11055_ _12094_/A _11055_/B vssd1 vssd1 vccd1 vccd1 _11059_/A sky130_fd_sc_hd__xnor2_1
X_10006_ _10004_/X _10005_/X _10176_/A vssd1 vssd1 vccd1 vccd1 _10006_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09910__A2 _10518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap55_A _07203_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11957_ _12742_/A _11957_/B _11957_/C vssd1 vssd1 vccd1 vccd1 _11957_/Y sky130_fd_sc_hd__nor3_1
X_10908_ _10909_/A _10909_/B vssd1 vssd1 vccd1 vccd1 _10908_/Y sky130_fd_sc_hd__nand2_1
X_11888_ _12710_/B2 _11364_/X _11377_/Y _09860_/A vssd1 vssd1 vccd1 vccd1 _11889_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_104_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13627_ _13725_/CLK _13627_/D vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__dfxtp_1
X_10839_ _10838_/A _10838_/B _10840_/A vssd1 vssd1 vccd1 vccd1 _10839_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_27_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10149__A _10631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10036__A2 _11587_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13558_ hold282/A _13557_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13558_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_82_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12509_ _12364_/X _12508_/X _12507_/Y vssd1 vssd1 vccd1 vccd1 _12509_/X sky130_fd_sc_hd__o21a_1
X_13489_ _13489_/A _13489_/B vssd1 vssd1 vccd1 vccd1 _13489_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__09729__A2 _07643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07458__A _10263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13179__B _13191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07177__B _07398_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout108 _11072_/A vssd1 vssd1 vccd1 vccd1 _10507_/A sky130_fd_sc_hd__buf_12
Xfanout119 _07456_/Y vssd1 vssd1 vccd1 vccd1 _09173_/B2 sky130_fd_sc_hd__buf_6
X_07981_ _08933_/B _11922_/A wire101/A _07175_/X vssd1 vssd1 vccd1 vccd1 _07982_/B
+ sky130_fd_sc_hd__a22o_1
X_09720_ curr_PC[0] curr_PC[1] vssd1 vssd1 vccd1 vccd1 _09720_/X sky130_fd_sc_hd__or2_1
X_06932_ reg1_val[13] _07522_/A vssd1 vssd1 vccd1 vccd1 _11373_/A sky130_fd_sc_hd__or2_1
XANTENNA__11708__A _11708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09362__B1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ _09001_/A _09001_/B _09986_/A _09316_/X _10150_/A vssd1 vssd1 vccd1 vccd1
+ _09654_/A sky130_fd_sc_hd__a2111o_1
X_06863_ _06863_/A _06863_/B vssd1 vssd1 vccd1 vccd1 _12218_/A sky130_fd_sc_hd__and2_2
X_08602_ _08642_/A vssd1 vssd1 vccd1 vccd1 _08602_/Y sky130_fd_sc_hd__inv_2
X_09582_ _09582_/A _10787_/B _10787_/C vssd1 vssd1 vccd1 vccd1 _09585_/B sky130_fd_sc_hd__or3_1
X_06794_ _06794_/A _06794_/B vssd1 vssd1 vccd1 vccd1 _12778_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_54_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08533_ _08866_/B2 fanout85/X fanout82/X _08950_/B vssd1 vssd1 vccd1 vccd1 _08534_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout160_A _13445_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_A _07535_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08464_ _08514_/B _08514_/A vssd1 vssd1 vccd1 vccd1 _08464_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_77_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07132__S _07135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07415_ _12421_/A _07422_/B vssd1 vssd1 vccd1 vccd1 _07415_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_108_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08395_ _09671_/S _08395_/B vssd1 vssd1 vccd1 vccd1 _08457_/B sky130_fd_sc_hd__nor2_1
X_07346_ _08907_/B _08907_/C vssd1 vssd1 vccd1 vccd1 _10104_/A sky130_fd_sc_hd__nor2_8
XFILLER_0_115_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07277_ _10542_/A _10366_/A _07275_/Y vssd1 vssd1 vccd1 vccd1 _09928_/A sky130_fd_sc_hd__o21bai_1
XFILLER_0_103_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09016_ _09016_/A _09016_/B _09016_/C vssd1 vssd1 vccd1 vccd1 _09017_/B sky130_fd_sc_hd__and3_1
XFILLER_0_60_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold140 hold140/A vssd1 vssd1 vccd1 vccd1 hold140/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 hold151/A vssd1 vssd1 vccd1 vccd1 hold151/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 hold162/A vssd1 vssd1 vccd1 vccd1 hold162/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 hold173/A vssd1 vssd1 vccd1 vccd1 hold173/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 hold184/A vssd1 vssd1 vccd1 vccd1 hold184/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 hold195/A vssd1 vssd1 vccd1 vccd1 hold195/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06954__A2 _06936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09918_ _09919_/A _09919_/B vssd1 vssd1 vccd1 vccd1 _10060_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08199__A _09949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10522__A _10522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09849_ _09847_/X _09848_/X _10176_/A vssd1 vssd1 vccd1 vccd1 _09849_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07903__A1 _10814_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07903__B2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12860_ reg1_val[9] curr_PC[9] _12867_/S vssd1 vssd1 vccd1 vccd1 _12862_/B sky130_fd_sc_hd__mux2_1
X_11811_ fanout20/X _07891_/X fanout10/X fanout18/X vssd1 vssd1 vccd1 vccd1 _11812_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ reg1_val[31] _07398_/B _09519_/Y vssd1 vssd1 vccd1 vccd1 _12791_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_96_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _11619_/A _11619_/B _11611_/A vssd1 vssd1 vccd1 vccd1 _11745_/A sky130_fd_sc_hd__o21bai_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _07094_/A _11566_/B _06919_/B vssd1 vssd1 vccd1 vccd1 _11674_/B sky130_fd_sc_hd__o21ai_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13204__A2 _13598_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10018__A2 _10010_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13412_ hold132/X _13416_/A2 _13420_/B1 hold107/X _13430_/C1 vssd1 vssd1 vccd1 vccd1
+ hold137/A sky130_fd_sc_hd__o221a_1
X_10624_ _10585_/Y _10623_/X _12867_/S vssd1 vssd1 vccd1 vccd1 _10624_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_107_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13343_ _13359_/A hold215/X vssd1 vssd1 vccd1 vccd1 _13653_/D sky130_fd_sc_hd__and2_1
XANTENNA__11800__B fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10555_ _10554_/B _10554_/C _10554_/A vssd1 vssd1 vccd1 vccd1 _10556_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13274_ hold83/X hold264/X vssd1 vssd1 vccd1 vccd1 _13274_/X sky130_fd_sc_hd__and2b_1
X_10486_ _10371_/A _10371_/B _10362_/X vssd1 vssd1 vccd1 vccd1 _10500_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__12715__A1 _09254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12225_ _12225_/A _12225_/B vssd1 vssd1 vccd1 vccd1 _12225_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09526__A2_N _11688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12156_ _12146_/Y _12147_/X _12151_/X _12155_/Y vssd1 vssd1 vccd1 vccd1 _12156_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__06945__A2 _06936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11107_ _11107_/A _11343_/A vssd1 vssd1 vccd1 vccd1 _11107_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12479__B1 _12971_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13446__C fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12087_ _12087_/A _12666_/A _12087_/C vssd1 vssd1 vccd1 vccd1 _12088_/B sky130_fd_sc_hd__nor3_1
X_11038_ _11038_/A _11038_/B vssd1 vssd1 vccd1 vccd1 _11039_/B sky130_fd_sc_hd__or2_1
XFILLER_0_91_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12989_ reg1_val[2] _12990_/B vssd1 vssd1 vccd1 vccd1 _12989_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_59_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13443__A2 _13445_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08870__A2 _09910_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07200_ _07200_/A _07200_/B vssd1 vssd1 vccd1 vccd1 _07200_/Y sky130_fd_sc_hd__nand2_2
X_08180_ _08866_/A2 fanout24/X _08486_/B _09216_/B2 vssd1 vssd1 vccd1 vccd1 _08181_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07131_ instruction[26] instruction[19] _07135_/S vssd1 vssd1 vccd1 vccd1 reg2_idx[1]
+ sky130_fd_sc_hd__mux2_8
XANTENNA__08083__B1 _08246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12094__A _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06804__B _13059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07062_ reg1_val[28] _07062_/B vssd1 vssd1 vccd1 vccd1 _07062_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_42_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07964_ _07964_/A _07964_/B vssd1 vssd1 vccd1 vccd1 _07965_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10342__A _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08138__A1 _08806_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08138__B2 _08806_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09703_ _12515_/S _09703_/B _09703_/C _09703_/D vssd1 vssd1 vccd1 vccd1 _09703_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__11157__B fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06915_ _07544_/A reg1_val[15] vssd1 vssd1 vccd1 vccd1 _11675_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07895_ _09659_/B _07895_/B _07895_/C vssd1 vssd1 vccd1 vccd1 _07897_/B sky130_fd_sc_hd__nand3_1
X_09634_ _09634_/A _09634_/B vssd1 vssd1 vccd1 vccd1 _09635_/B sky130_fd_sc_hd__nor2_2
X_06846_ _07410_/A _07221_/A vssd1 vssd1 vccd1 vccd1 _06847_/B sky130_fd_sc_hd__nor2_1
X_09565_ _09359_/A _09359_/B _09358_/A vssd1 vssd1 vccd1 vccd1 _09567_/B sky130_fd_sc_hd__o21a_1
X_06777_ instruction[0] instruction[2] instruction[1] pred_val vssd1 vssd1 vccd1 vccd1
+ _06920_/B sky130_fd_sc_hd__or4bb_4
XANTENNA__13434__A2 _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08516_ _08458_/B _08516_/B vssd1 vssd1 vccd1 vccd1 _08517_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_77_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09496_ _09488_/X _10176_/B _09496_/S vssd1 vssd1 vccd1 vccd1 _09496_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11996__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08447_ _08447_/A vssd1 vssd1 vccd1 vccd1 _08506_/A sky130_fd_sc_hd__inv_2
XFILLER_0_93_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13198__A1 _12496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11901__A _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08482__A _10542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08378_ _08379_/A _08379_/B vssd1 vssd1 vccd1 vccd1 _08378_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08074__B1 _08704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07329_ reg1_val[16] reg1_val[17] vssd1 vssd1 vccd1 vccd1 _07435_/B sky130_fd_sc_hd__or2_4
XFILLER_0_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10340_ curr_PC[4] curr_PC[5] _10340_/C vssd1 vssd1 vccd1 vccd1 _10480_/B sky130_fd_sc_hd__and3_1
XFILLER_0_116_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07821__B1 _09885_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10271_ _10271_/A _10271_/B vssd1 vssd1 vccd1 vccd1 _10274_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09574__B1 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12010_ _12010_/A _12010_/B vssd1 vssd1 vccd1 vccd1 _12011_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13122__B2 _07634_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12912_ _12912_/A _12912_/B _12912_/C vssd1 vssd1 vccd1 vccd1 _12913_/B sky130_fd_sc_hd__nand3_1
X_12843_ _12844_/A _12844_/B _12844_/C vssd1 vssd1 vccd1 vccd1 _12851_/B sky130_fd_sc_hd__a21o_1
XANTENNA__13425__A2 _13445_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _12732_/Y _12733_/X _12770_/X _12772_/Y _12374_/A vssd1 vssd1 vccd1 vccd1
+ _12774_/X sky130_fd_sc_hd__o221a_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _11725_/A _11725_/B vssd1 vssd1 vccd1 vccd1 _11727_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_84_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08852__A2 _10104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11656_ _11657_/A _11657_/B vssd1 vssd1 vccd1 vccd1 _11758_/B sky130_fd_sc_hd__or2_1
XFILLER_0_36_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06905__A _06928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout90 _07433_/X vssd1 vssd1 vccd1 vccd1 _11507_/A sky130_fd_sc_hd__buf_6
XANTENNA__08065__B1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10607_ _06979_/B _12793_/A2 _11586_/B vssd1 vssd1 vccd1 vccd1 _10607_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09801__A1 _09604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11587_ _06919_/B _11587_/A2 _12657_/B1 reg1_val[15] _11586_/Y vssd1 vssd1 vccd1
+ vccd1 _11587_/X sky130_fd_sc_hd__o221a_1
XANTENNA__10947__B1 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13326_ hold226/X _13463_/B2 _13450_/B hold238/X vssd1 vssd1 vccd1 vccd1 hold239/A
+ sky130_fd_sc_hd__a22o_1
X_10538_ _10538_/A _10787_/B _10787_/C vssd1 vssd1 vccd1 vccd1 _10541_/B sky130_fd_sc_hd__or3_1
XFILLER_0_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13257_ hold51/X hold291/A vssd1 vssd1 vccd1 vccd1 _13257_/X sky130_fd_sc_hd__and2b_1
X_10469_ _10335_/A _10332_/Y _10334_/B vssd1 vssd1 vccd1 vccd1 _10473_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_86_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07736__A _10078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12208_ _12208_/A _12208_/B vssd1 vssd1 vccd1 vccd1 _12208_/X sky130_fd_sc_hd__and2_1
X_13188_ _07198_/Y _13196_/A2 hold86/X _13591_/A vssd1 vssd1 vccd1 vccd1 hold87/A
+ sky130_fd_sc_hd__o211a_1
X_12139_ reg1_val[21] curr_PC[21] vssd1 vssd1 vccd1 vccd1 _12140_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07591__A2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09951__A _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07879__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07680_ _07680_/A _07680_/B vssd1 vssd1 vccd1 vccd1 _07714_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09350_ _07230_/Y _10536_/A1 _10536_/B2 _12331_/A vssd1 vssd1 vccd1 vccd1 _09351_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08301_ _08301_/A _08301_/B vssd1 vssd1 vccd1 vccd1 _08358_/A sky130_fd_sc_hd__nand2_2
XANTENNA__10613__B1_N _10609_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09281_ _10915_/A fanout21/X _08246_/B _11047_/A vssd1 vssd1 vccd1 vccd1 _09282_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08232_ _08232_/A _08232_/B vssd1 vssd1 vccd1 vccd1 _08297_/B sky130_fd_sc_hd__xor2_1
XANTENNA__11721__A _12253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10650__A2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08163_ _08169_/B _08169_/A vssd1 vssd1 vccd1 vccd1 _08234_/B sky130_fd_sc_hd__and2b_1
XANTENNA__08056__B1 _08118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout123_A _07451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07114_ _13748_/A _07123_/B _09514_/B vssd1 vssd1 vccd1 vccd1 _13142_/B sky130_fd_sc_hd__and3_1
XFILLER_0_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10402__A2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08094_ _08096_/A _08096_/B vssd1 vssd1 vccd1 vccd1 _08094_/X sky130_fd_sc_hd__and2b_1
XANTENNA__07349__C _13082_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07045_ _06923_/X _07044_/X _06918_/X vssd1 vssd1 vccd1 vccd1 _11675_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_113_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12155__A2 _12754_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07031__B2 _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08996_ _08997_/A _08997_/B vssd1 vssd1 vccd1 vccd1 _08996_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_76_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07947_ _07506_/A _07506_/B _07505_/A vssd1 vssd1 vccd1 vccd1 _07952_/A sky130_fd_sc_hd__a21o_2
XANTENNA__09859__A1 _12525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10800__A _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07878_ _12617_/A _11823_/A _07876_/Y vssd1 vssd1 vccd1 vccd1 _07878_/X sky130_fd_sc_hd__a21o_1
XANTENNA__08477__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09617_ _09631_/A vssd1 vssd1 vccd1 vccd1 _09617_/Y sky130_fd_sc_hd__inv_2
X_06829_ reg1_val[25] _07252_/B vssd1 vssd1 vccd1 vccd1 _06831_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09548_ _07699_/B _10522_/A _07557_/Y fanout35/X vssd1 vssd1 vccd1 vccd1 _09549_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout36_A _08118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12091__A1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09479_ _09477_/X _09478_/X _09688_/S vssd1 vssd1 vccd1 vccd1 _09479_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12091__B2 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11510_ _11510_/A _11510_/B vssd1 vssd1 vccd1 vccd1 _11524_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_108_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12490_ _12491_/A _12491_/B _12491_/C vssd1 vssd1 vccd1 vccd1 _12565_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11441_ _11441_/A _11441_/B vssd1 vssd1 vccd1 vccd1 _11443_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08598__A1 _08806_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08598__B2 _08806_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09795__B1 _07478_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11372_ _11372_/A _11372_/B _12598_/C vssd1 vssd1 vccd1 vccd1 _11372_/X sky130_fd_sc_hd__or3_2
XANTENNA__08940__A _09371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13111_ _13111_/A _13111_/B vssd1 vssd1 vccd1 vccd1 _13121_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10323_ hold182/A _10323_/B vssd1 vssd1 vccd1 vccd1 _10323_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__12462__A _12782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13042_ reg1_val[12] _13042_/B vssd1 vssd1 vccd1 vccd1 _13051_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07556__A _07556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10254_ _10255_/A _10255_/B vssd1 vssd1 vccd1 vccd1 _10254_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10185_ _07003_/B _12793_/A2 _11586_/B vssd1 vssd1 vccd1 vccd1 _10185_/Y sky130_fd_sc_hd__a21oi_1
Xfanout280 _13568_/A vssd1 vssd1 vccd1 vccd1 _13605_/A sky130_fd_sc_hd__buf_4
Xfanout291 reg1_val[0] vssd1 vssd1 vccd1 vccd1 _09501_/A sky130_fd_sc_hd__buf_8
XANTENNA__08522__A1 _09910_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07291__A _10542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08522__B2 _07420_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12826_ _13000_/B _12827_/B vssd1 vssd1 vccd1 vccd1 _12837_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_57_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ _13129_/A _09254_/A _09515_/Y _12755_/X _12756_/Y vssd1 vssd1 vccd1 vccd1
+ _12757_/X sky130_fd_sc_hd__a311o_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11708_ _11708_/A _11709_/B vssd1 vssd1 vccd1 vccd1 _11708_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12688_ _12733_/A _12635_/A _12733_/B _12634_/X _12735_/A1 vssd1 vssd1 vccd1 vccd1
+ _12688_/X sky130_fd_sc_hd__o41a_1
XFILLER_0_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11639_ _07547_/X _11802_/B _11638_/C vssd1 vssd1 vccd1 vccd1 _11640_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08589__A1 _07238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08589__B2 _07239_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09250__A2 _12614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13309_ _13222_/B _13565_/B _13222_/A vssd1 vssd1 vccd1 vccd1 _13570_/A sky130_fd_sc_hd__o21bai_2
XANTENNA__12372__A _12372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07466__A _11508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13187__B _13191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08850_ _08850_/A _08850_/B vssd1 vssd1 vccd1 vccd1 _08857_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07801_ _08806_/A2 _07544_/Y _11638_/A _08806_/B1 vssd1 vssd1 vccd1 vccd1 _07802_/B
+ sky130_fd_sc_hd__a22o_1
X_08781_ _08791_/A _08818_/A _08781_/C vssd1 vssd1 vccd1 vccd1 _08781_/X sky130_fd_sc_hd__and3_1
X_07732_ _07744_/B _07732_/B vssd1 vssd1 vccd1 vccd1 _07811_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11716__A _12092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07663_ _09591_/A _07663_/B vssd1 vssd1 vccd1 vccd1 _07667_/B sky130_fd_sc_hd__xnor2_1
X_09402_ _09402_/A _09402_/B vssd1 vssd1 vccd1 vccd1 _09405_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07594_ _09254_/C _07594_/B vssd1 vssd1 vccd1 vccd1 _07595_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_87_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09333_ _11731_/A _09333_/B vssd1 vssd1 vccd1 vccd1 _09337_/A sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout240_A _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09264_ _09264_/A _09264_/B vssd1 vssd1 vccd1 vccd1 _09278_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_62_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08215_ _08258_/B vssd1 vssd1 vccd1 vccd1 _08216_/B sky130_fd_sc_hd__inv_2
X_09195_ _09195_/A _09195_/B vssd1 vssd1 vccd1 vccd1 _09197_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09777__B1 _10536_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08146_ _10522_/A _08580_/B _08868_/B1 fanout84/X vssd1 vssd1 vccd1 vccd1 _08147_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_71_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10387__A1 _07282_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10387__B2 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11584__B1 _12533_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08077_ _10522_/A fanout84/X _08580_/B _09885_/B1 vssd1 vssd1 vccd1 vccd1 _08078_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_3_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07028_ _06928_/A _06928_/B _12806_/A _07027_/X vssd1 vssd1 vccd1 vccd1 _07028_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_0_30_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13097__B _13129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__09591__A _09591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ _08724_/X _09044_/A _09041_/B _08723_/X _08725_/A vssd1 vssd1 vccd1 vccd1
+ _09049_/A sky130_fd_sc_hd__a32o_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11626__A _12092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__A1 _07547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11990_ _12253_/A _11990_/B vssd1 vssd1 vccd1 vccd1 _11994_/A sky130_fd_sc_hd__xnor2_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
X_10941_ _10941_/A _10941_/B vssd1 vssd1 vccd1 vccd1 _10959_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08000__A _11708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13660_ _13717_/CLK hold187/X vssd1 vssd1 vccd1 vccd1 _13660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10872_ _10742_/A _10739_/Y _10741_/B vssd1 vssd1 vccd1 vccd1 _10876_/A sky130_fd_sc_hd__o21a_1
XANTENNA__09530__S _09703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12611_ _12612_/A _12612_/B vssd1 vssd1 vccd1 vccd1 _12675_/A sky130_fd_sc_hd__and2_1
XANTENNA__08268__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13591_ _13591_/A hold141/X vssd1 vssd1 vccd1 vccd1 hold142/A sky130_fd_sc_hd__and2_1
XFILLER_0_54_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10075__B1 _08704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12542_ curr_PC[26] _12543_/B vssd1 vssd1 vccd1 vccd1 _12544_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10614__A2 _11587_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11811__A1 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11811__B2 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12473_ _09504_/Y _12462_/B _10458_/X _12710_/B2 _12472_/X vssd1 vssd1 vccd1 vccd1
+ _12473_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_34_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11424_ _11424_/A _11424_/B vssd1 vssd1 vccd1 vccd1 _11426_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_8 instruction[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07243__A1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07243__B2 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08440__B1 _08778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11355_ _11463_/A _06939_/Y _07042_/X _11354_/Y vssd1 vssd1 vccd1 vccd1 _11356_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07794__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10306_ _11864_/A _10306_/B _10306_/C vssd1 vssd1 vccd1 vccd1 _10306_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_21_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11286_ _11286_/A _11286_/B _11286_/C vssd1 vssd1 vccd1 vccd1 _11288_/B sky130_fd_sc_hd__nand3_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13025_ reg1_val[9] _13025_/B vssd1 vssd1 vccd1 vccd1 _13033_/A sky130_fd_sc_hd__nand2_1
X_10237_ _10536_/A1 _12614_/A _12667_/A _10536_/B2 vssd1 vssd1 vccd1 vccd1 _10238_/B
+ sky130_fd_sc_hd__a22o_1
X_10168_ reg1_val[4] curr_PC[4] vssd1 vssd1 vccd1 vccd1 _10169_/B sky130_fd_sc_hd__nand2_1
X_10099_ _10099_/A _10099_/B vssd1 vssd1 vccd1 vccd1 _10100_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_88_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12809_ _12809_/A _12809_/B vssd1 vssd1 vccd1 vccd1 _12810_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12055__A1 _12056_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08000_ _11708_/A _08000_/B vssd1 vssd1 vccd1 vccd1 _08006_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08580__A _09674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08431__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06812__B _09254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09951_ _09951_/A _09951_/B vssd1 vssd1 vccd1 vccd1 _09953_/B sky130_fd_sc_hd__xnor2_2
X_08902_ _08902_/A _08902_/B vssd1 vssd1 vccd1 vccd1 _08911_/B sky130_fd_sc_hd__xnor2_1
X_09882_ _09822_/A _09822_/B _09820_/X vssd1 vssd1 vccd1 vccd1 _09985_/A sky130_fd_sc_hd__a21oi_4
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08734__A1 _08821_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ _09381_/A _08833_/B vssd1 vssd1 vccd1 vccd1 _08834_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08734__B2 _08821_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07643__B _07643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08764_ _08764_/A _08764_/B vssd1 vssd1 vccd1 vccd1 _08789_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_79_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07135__S _07135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07715_ _07715_/A _07715_/B vssd1 vssd1 vccd1 vccd1 _07719_/B sky130_fd_sc_hd__nand2_1
X_08695_ _08724_/A _08724_/B vssd1 vssd1 vccd1 vccd1 _08725_/A sky130_fd_sc_hd__or2_1
X_07646_ _07870_/A _07646_/B vssd1 vssd1 vccd1 vccd1 _07647_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_95_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07577_ _10934_/A _07577_/B vssd1 vssd1 vccd1 vccd1 _07577_/X sky130_fd_sc_hd__or2_2
XFILLER_0_75_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09316_ _09318_/A _09825_/A vssd1 vssd1 vccd1 vccd1 _09316_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09247_ _09248_/A _09248_/B vssd1 vssd1 vccd1 vccd1 _09249_/A sky130_fd_sc_hd__or2_1
XFILLER_0_90_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11006__C1 _12533_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09178_ _09179_/A _09179_/B _09179_/C vssd1 vssd1 vccd1 vccd1 _09301_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09214__A2 _07451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07225__A1 _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08129_ _08130_/A _08129_/B _08129_/C vssd1 vssd1 vccd1 vccd1 _08174_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_121_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07225__B2 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08422__B1 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10525__A _12551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11140_ _07093_/A _09509_/X _11587_/A2 _06950_/B _11139_/X vssd1 vssd1 vccd1 vccd1
+ _11140_/X sky130_fd_sc_hd__o221a_1
X_11071_ _10787_/A fanout10/X fanout5/X _07546_/X vssd1 vssd1 vccd1 vccd1 _11072_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07528__A2 _07522_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10022_ _10022_/A vssd1 vssd1 vccd1 vccd1 _10022_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06883__A_N _07281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11973_ _12311_/B1 _12148_/C _13660_/Q vssd1 vssd1 vccd1 vccd1 _11975_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10924_ _10925_/A _10925_/B vssd1 vssd1 vccd1 vccd1 _10924_/X sky130_fd_sc_hd__and2_1
X_13712_ _13736_/CLK _13712_/D vssd1 vssd1 vccd1 vccd1 hold301/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10855_ _10981_/B _10981_/C vssd1 vssd1 vccd1 vccd1 _11107_/A sky130_fd_sc_hd__nor2_1
X_13643_ _13649_/CLK _13643_/D vssd1 vssd1 vccd1 vccd1 hold243/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13574_ _13311_/B _13574_/B vssd1 vssd1 vccd1 vccd1 _13575_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_26_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10786_ _11076_/A _10786_/B vssd1 vssd1 vccd1 vccd1 _10794_/A sky130_fd_sc_hd__xnor2_2
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11796__B1 _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12525_ _12525_/A _12525_/B vssd1 vssd1 vccd1 vccd1 _12525_/Y sky130_fd_sc_hd__nor2_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13510__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12456_ _09082_/A _12454_/X _12455_/Y vssd1 vssd1 vccd1 vccd1 _12476_/C sky130_fd_sc_hd__a21oi_4
XFILLER_0_124_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11407_ _11521_/A _11521_/B vssd1 vssd1 vccd1 vccd1 _11415_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11012__A2 _11587_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12387_ _12385_/Y _12387_/B vssd1 vssd1 vccd1 vccd1 _12388_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_22_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07767__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11338_ _11340_/A _11340_/B _11340_/C vssd1 vssd1 vccd1 vccd1 _11341_/A sky130_fd_sc_hd__a21oi_1
Xclkbuf_4_9_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13700_/CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA__10771__A1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10771__B2 _12557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11269_ _13180_/A1 fanout16/X _07877_/X _07548_/X vssd1 vssd1 vccd1 vccd1 _11270_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_13008_ _13007_/A _13004_/Y _13006_/B vssd1 vssd1 vccd1 vccd1 _13012_/A sky130_fd_sc_hd__o21a_2
XANTENNA__11976__A2_N _11688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11720__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08192__A2 _07541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11266__A _12867_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07500_ _07500_/A _07500_/B vssd1 vssd1 vccd1 vccd1 _07502_/B sky130_fd_sc_hd__nand2_1
X_08480_ _08480_/A _08480_/B vssd1 vssd1 vccd1 vccd1 _08551_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07152__B1 _10889_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07431_ reg1_val[18] _07634_/B _07435_/B reg1_val[19] vssd1 vssd1 vccd1 vccd1 _07431_/Y
+ sky130_fd_sc_hd__o31ai_4
XFILLER_0_76_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06807__B _09254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07362_ _12177_/A _07368_/B _12252_/A vssd1 vssd1 vccd1 vccd1 _07362_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09101_ _07912_/A _07912_/B _07910_/Y vssd1 vssd1 vccd1 vccd1 _09116_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_127_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07293_ reg1_val[8] reg1_val[9] vssd1 vssd1 vccd1 vccd1 _07320_/D sky130_fd_sc_hd__or2_2
XFILLER_0_72_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09032_ _09034_/A _11233_/A _11117_/B vssd1 vssd1 vccd1 vccd1 _09032_/X sky130_fd_sc_hd__or3b_1
XANTENNA__07919__A _10119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold300 hold300/A vssd1 vssd1 vccd1 vccd1 hold300/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout203_A _12799_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08955__B2 _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09934_ _09934_/A _09934_/B vssd1 vssd1 vccd1 vccd1 _09935_/B sky130_fd_sc_hd__or2_1
XFILLER_0_110_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08707__A1 _07239_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08707__B2 _07238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09904__B1 _07522_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06981__A3 _13015_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09865_ _12515_/S _09865_/B vssd1 vssd1 vccd1 vccd1 _09865_/Y sky130_fd_sc_hd__nand2_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11176__A _11913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08816_ _08846_/A _08816_/B vssd1 vssd1 vccd1 vccd1 _08838_/A sky130_fd_sc_hd__xnor2_1
X_09796_ _10119_/A _09796_/B vssd1 vssd1 vccd1 vccd1 _09798_/B sky130_fd_sc_hd__xnor2_1
X_08747_ _08753_/A _08753_/B vssd1 vssd1 vccd1 vccd1 _08747_/Y sky130_fd_sc_hd__nand2_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ _08701_/A _08701_/B _08674_/X vssd1 vssd1 vccd1 vccd1 _08690_/B sky130_fd_sc_hd__a21o_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07629_ _07630_/A _07630_/B vssd1 vssd1 vccd1 vccd1 _07940_/B sky130_fd_sc_hd__or2_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10640_ _10641_/A _10641_/B vssd1 vssd1 vccd1 vccd1 _10780_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_36_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10571_ _10571_/A _10571_/B vssd1 vssd1 vccd1 vccd1 _10572_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_91_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08932__B _08933_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12310_ _10758_/X _12309_/Y _12782_/B vssd1 vssd1 vccd1 vccd1 _12310_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13290_ _13478_/B _13479_/A _13267_/X vssd1 vssd1 vccd1 vccd1 _13484_/A sky130_fd_sc_hd__a21o_1
X_12241_ _12241_/A _12241_/B _12241_/C _12241_/D vssd1 vssd1 vccd1 vccd1 _12241_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_106_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12172_ _12173_/A _12173_/B _12173_/C vssd1 vssd1 vccd1 vccd1 _12174_/A sky130_fd_sc_hd__a21o_1
X_11123_ _11122_/A _11122_/B _11122_/Y _12047_/C1 vssd1 vssd1 vccd1 vccd1 _11123_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13152__C1 _13543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11054_ fanout53/X fanout20/X fanout18/X fanout47/X vssd1 vssd1 vccd1 vccd1 _11055_/B
+ sky130_fd_sc_hd__o22a_1
X_10005_ _09679_/X _09681_/X _10005_/S vssd1 vssd1 vccd1 vccd1 _10005_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13505__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11814__A _12092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11466__C1 _12047_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08395__A _09671_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11956_ _12742_/A _11957_/B _11957_/C vssd1 vssd1 vccd1 vccd1 _11956_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_98_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10907_ _12668_/A _10907_/B vssd1 vssd1 vccd1 vccd1 _10909_/B sky130_fd_sc_hd__xnor2_1
X_11887_ _07092_/B _12709_/A2 _11884_/X _11886_/X vssd1 vssd1 vccd1 vccd1 _11887_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10838_ _10838_/A _10838_/B vssd1 vssd1 vccd1 vccd1 _10840_/B sky130_fd_sc_hd__nor2_1
X_13626_ _13725_/CLK _13626_/D vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10769_ fanout46/X fanout25/X fanout23/X fanout50/X vssd1 vssd1 vccd1 vccd1 _10770_/B
+ sky130_fd_sc_hd__o22a_1
X_13557_ _13557_/A _13557_/B vssd1 vssd1 vccd1 vccd1 _13557_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12508_ _12508_/A _12570_/A vssd1 vssd1 vccd1 vccd1 _12508_/X sky130_fd_sc_hd__or2_1
XFILLER_0_125_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13488_ _13263_/X _13488_/B vssd1 vssd1 vccd1 vccd1 _13489_/B sky130_fd_sc_hd__nand2b_1
X_12439_ _12442_/A _12508_/A vssd1 vssd1 vccd1 vccd1 _12440_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_1_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07980_ _07991_/B _07991_/A vssd1 vssd1 vccd1 vccd1 _07980_/X sky130_fd_sc_hd__and2b_1
Xfanout109 _07510_/Y vssd1 vssd1 vccd1 vccd1 _11072_/A sky130_fd_sc_hd__buf_8
X_06931_ reg1_val[13] _07523_/A vssd1 vssd1 vccd1 vccd1 _06931_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13195__B _13207_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09362__A1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09362__B2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09650_ _09650_/A _09650_/B vssd1 vssd1 vccd1 vccd1 _10298_/A sky130_fd_sc_hd__xnor2_4
X_06862_ _07357_/A _07212_/B vssd1 vssd1 vccd1 vccd1 _06863_/B sky130_fd_sc_hd__nand2_1
X_08601_ _08647_/A _08647_/B _08597_/Y vssd1 vssd1 vccd1 vccd1 _08642_/A sky130_fd_sc_hd__o21ai_2
X_09581_ _09951_/A _09581_/B vssd1 vssd1 vccd1 vccd1 _09588_/A sky130_fd_sc_hd__xnor2_1
X_06793_ _13135_/A _07398_/B vssd1 vssd1 vccd1 vccd1 _06794_/B sky130_fd_sc_hd__nand2_1
X_08532_ _08532_/A _08532_/B vssd1 vssd1 vccd1 vccd1 _08606_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08463_ _08463_/A _08463_/B vssd1 vssd1 vccd1 vccd1 _08514_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08873__B1 _08891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07414_ _07414_/A _07414_/B _07414_/C _07414_/D vssd1 vssd1 vccd1 vccd1 _07422_/B
+ sky130_fd_sc_hd__nand4_4
X_08394_ _09940_/A _08394_/B vssd1 vssd1 vccd1 vccd1 _08457_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07345_ _07186_/B _07594_/B _10603_/S vssd1 vssd1 vccd1 vccd1 _08907_/C sky130_fd_sc_hd__and3b_2
X_07276_ _10542_/A _10366_/A _07275_/Y vssd1 vssd1 vccd1 vccd1 _07276_/X sky130_fd_sc_hd__o21ba_2
XFILLER_0_72_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09015_ _09016_/A _09016_/B _09016_/C vssd1 vssd1 vccd1 vccd1 _09017_/A sky130_fd_sc_hd__a21oi_1
Xhold130 hold130/A vssd1 vssd1 vccd1 vccd1 hold130/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 hold141/A vssd1 vssd1 vccd1 vccd1 hold141/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10735__A1 _10734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold152 hold152/A vssd1 vssd1 vccd1 vccd1 hold152/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 hold163/A vssd1 vssd1 vccd1 vccd1 hold163/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 hold174/A vssd1 vssd1 vccd1 vccd1 hold174/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 hold203/X vssd1 vssd1 vccd1 vccd1 hold185/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10803__A _11825_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold196 hold196/A vssd1 vssd1 vccd1 vccd1 hold196/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06954__A3 _13036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09917_ _09800_/A _09799_/B _09797_/X vssd1 vssd1 vccd1 vccd1 _09919_/B sky130_fd_sc_hd__a21o_1
XANTENNA__10522__B _10522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09848_ _09472_/X _09476_/X _10005_/S vssd1 vssd1 vccd1 vccd1 _09848_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07364__B1 _07476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout66_A _08778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07903__A2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09779_ _09779_/A _09780_/B vssd1 vssd1 vccd1 vccd1 _09779_/X sky130_fd_sc_hd__and2_1
XFILLER_0_68_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11810_ _11810_/A vssd1 vssd1 vccd1 vccd1 _11819_/A sky130_fd_sc_hd__inv_2
X_12790_ reg1_val[31] _11688_/B _12799_/A2 vssd1 vssd1 vccd1 vccd1 _12790_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _11637_/A _11637_/B _11640_/A vssd1 vssd1 vccd1 vccd1 _11746_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12660__A1 _12710_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10671__B1 _08580_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11672_ _11672_/A _11672_/B vssd1 vssd1 vccd1 vccd1 _11672_/Y sky130_fd_sc_hd__xnor2_2
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10623_ _10586_/Y _10587_/X _10593_/X _10622_/X vssd1 vssd1 vccd1 vccd1 _10623_/X
+ sky130_fd_sc_hd__a211o_1
X_13411_ _07516_/Y _13419_/A2 hold133/X vssd1 vssd1 vccd1 vccd1 _13687_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_119_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07559__A _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13342_ hold209/X _13506_/B2 _13506_/A2 hold214/X vssd1 vssd1 vccd1 vccd1 hold215/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10554_ _10554_/A _10554_/B _10554_/C vssd1 vssd1 vccd1 vccd1 _10556_/A sky130_fd_sc_hd__and3_1
XFILLER_0_24_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13273_ _13271_/X _13273_/B vssd1 vssd1 vccd1 vccd1 _13469_/A sky130_fd_sc_hd__nand2b_1
X_10485_ _10424_/A _10424_/B _10425_/X vssd1 vssd1 vccd1 vccd1 _10572_/A sky130_fd_sc_hd__o21bai_4
XFILLER_0_121_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12715__A2 _12799_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12224_ _12224_/A _12224_/B vssd1 vssd1 vccd1 vccd1 _12224_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_121_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12155_ _07351_/X _12754_/C _12154_/X vssd1 vssd1 vccd1 vccd1 _12155_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11809__A _12253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11106_ _11106_/A _11225_/A vssd1 vssd1 vccd1 vccd1 _11343_/A sky130_fd_sc_hd__nor2_1
XANTENNA__06945__A3 _13042_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12086_ _12173_/B _12086_/B vssd1 vssd1 vccd1 vccd1 _12088_/A sky130_fd_sc_hd__nand2_1
X_11037_ _11038_/A _11038_/B vssd1 vssd1 vccd1 vccd1 _11161_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13428__B1 _13444_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12988_ _12987_/A _12986_/B _12984_/Y vssd1 vssd1 vccd1 vccd1 _12992_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_47_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11939_ _11940_/A _11940_/B vssd1 vssd1 vccd1 vccd1 _12032_/A sky130_fd_sc_hd__and2_1
XFILLER_0_59_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09949__A _09949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08853__A _09371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12403__A1 _12760_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13609_ _13705_/CLK hold14/X vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07130_ instruction[25] instruction[18] _07135_/S vssd1 vssd1 vccd1 vccd1 reg2_idx[0]
+ sky130_fd_sc_hd__mux2_8
XFILLER_0_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08083__A1 _08873_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08083__B2 _07406_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07061_ reg1_val[29] _07061_/B vssd1 vssd1 vccd1 vccd1 _07061_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_112_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12167__B1 _07699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11719__A _11719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07963_ _07963_/A _07963_/B vssd1 vssd1 vccd1 vccd1 _08999_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08138__A2 _07477_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09702_ _12515_/S _09703_/B _09703_/C _09703_/D vssd1 vssd1 vccd1 vccd1 _09702_/Y
+ sky130_fd_sc_hd__a22oi_1
X_06914_ _06936_/A _13082_/A _06928_/B _06913_/X vssd1 vssd1 vccd1 vccd1 _07544_/A
+ sky130_fd_sc_hd__a31o_4
X_07894_ _08907_/A _10787_/B _10787_/C vssd1 vssd1 vccd1 vccd1 _07895_/C sky130_fd_sc_hd__or3_1
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09633_ _09633_/A _09633_/B vssd1 vssd1 vccd1 vccd1 _09634_/B sky130_fd_sc_hd__nor2_1
X_06845_ reg1_val[24] _07252_/D vssd1 vssd1 vccd1 vccd1 _06847_/A sky130_fd_sc_hd__nor2_1
XANTENNA_fanout270_A _06936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09564_ _09402_/A _09402_/B _09400_/Y vssd1 vssd1 vccd1 vccd1 _09567_/A sky130_fd_sc_hd__o21a_1
X_06776_ instruction[0] instruction[2] instruction[1] pred_val vssd1 vssd1 vccd1 vccd1
+ _06776_/X sky130_fd_sc_hd__and4bb_1
XFILLER_0_77_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08515_ _08569_/A _08569_/B vssd1 vssd1 vccd1 vccd1 _08515_/X sky130_fd_sc_hd__and2_1
XFILLER_0_78_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09495_ _09491_/X _09494_/X _10007_/S vssd1 vssd1 vccd1 vccd1 _10176_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_93_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08446_ _11072_/A _08446_/B vssd1 vssd1 vccd1 vccd1 _08447_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13198__A2 _13598_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08377_ _08377_/A _08377_/B vssd1 vssd1 vccd1 vccd1 _08379_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07328_ _11126_/A _07328_/B _07328_/C _07328_/D vssd1 vssd1 vccd1 vccd1 _07634_/B
+ sky130_fd_sc_hd__or4_4
XANTENNA__08074__A1 _10049_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08074__B2 _09173_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07259_ _09950_/A _07259_/B vssd1 vssd1 vccd1 vccd1 _07261_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_21_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07821__A1 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07821__B2 _08486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09594__A _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10270_ _10270_/A _10270_/B vssd1 vssd1 vccd1 vccd1 _10271_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09574__A1 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09574__B2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11381__A1 _10730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12911_ _12912_/A _12912_/B _12912_/C vssd1 vssd1 vccd1 vccd1 _12922_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_69_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10892__B1 _09520_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12842_ _12851_/A _12842_/B vssd1 vssd1 vccd1 vccd1 _12844_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_96_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _12773_/A _12773_/B vssd1 vssd1 vccd1 vccd1 _12773_/X sky130_fd_sc_hd__or2_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _11724_/A _11724_/B vssd1 vssd1 vccd1 vccd1 _11725_/B sky130_fd_sc_hd__and2_1
XANTENNA__08673__A _08746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ _11544_/A _11543_/B _11543_/A vssd1 vssd1 vccd1 vccd1 _11657_/B sky130_fd_sc_hd__o21ba_1
Xfanout80 _07524_/Y vssd1 vssd1 vccd1 vccd1 _08580_/B sky130_fd_sc_hd__buf_8
XFILLER_0_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06905__B _12806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout91 _12420_/A vssd1 vssd1 vccd1 vccd1 _12092_/A sky130_fd_sc_hd__buf_12
XFILLER_0_126_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08065__A1 _08866_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10606_ hold180/A _10606_/A2 _10882_/C _12533_/B1 vssd1 vssd1 vccd1 vccd1 _10606_/X
+ sky130_fd_sc_hd__a31o_1
X_11586_ _11586_/A _11586_/B vssd1 vssd1 vccd1 vccd1 _11586_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10947__A1 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09801__A2 _10518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10947__B2 _12557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10537_ _10537_/A _10537_/B vssd1 vssd1 vccd1 vccd1 _10544_/A sky130_fd_sc_hd__xor2_2
X_13325_ _13459_/A hold227/X vssd1 vssd1 vccd1 vccd1 hold228/A sky130_fd_sc_hd__and2_1
XFILLER_0_101_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10468_ _06986_/Y _11587_/A2 _10462_/Y _10590_/A _10467_/X vssd1 vssd1 vccd1 vccd1
+ _10468_/X sky130_fd_sc_hd__o221a_1
X_13256_ hold271/X hold57/X vssd1 vssd1 vccd1 vccd1 _13508_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_86_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12207_ _12207_/A _12207_/B _12440_/A vssd1 vssd1 vccd1 vccd1 _12208_/B sky130_fd_sc_hd__nand3_1
X_13187_ hold85/X _13191_/B vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__or2_1
X_10399_ _10253_/A _10253_/B _10254_/Y vssd1 vssd1 vccd1 vccd1 _10414_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_20_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12138_ reg1_val[21] curr_PC[21] vssd1 vssd1 vccd1 vccd1 _12140_/A sky130_fd_sc_hd__or2_1
XANTENNA__13113__A2 _07378_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12069_ curr_PC[19] _12070_/C curr_PC[20] vssd1 vssd1 vccd1 vccd1 _12071_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__09868__A2 _12793_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07879__A1 _09604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07879__B2 _09161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08300_ _08300_/A _08300_/B vssd1 vssd1 vccd1 vccd1 _08301_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10635__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09280_ _09108_/A _09108_/B _09111_/A vssd1 vssd1 vccd1 vccd1 _09293_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__11978__A3 _12754_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08231_ _08229_/A _08229_/B _08230_/X vssd1 vssd1 vccd1 vccd1 _08297_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_51_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10618__A _13015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08162_ _08162_/A _08162_/B vssd1 vssd1 vccd1 vccd1 _08169_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08056__A1 _09381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08056__B2 _08873_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07113_ _13748_/A _09514_/B vssd1 vssd1 vccd1 vccd1 _09523_/B sky130_fd_sc_hd__nand2_2
X_08093_ _08093_/A _08093_/B vssd1 vssd1 vccd1 vccd1 _08096_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_113_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12833__A _13005_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout116_A _11508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07044_ _06931_/Y _07043_/X _11465_/A vssd1 vssd1 vccd1 vccd1 _07044_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_11_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13352__A2 _13506_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10353__A _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08995_ _08991_/X _08993_/X _08167_/X vssd1 vssd1 vccd1 vccd1 _09089_/A sky130_fd_sc_hd__a21oi_4
X_07946_ _07651_/A _07650_/B _07648_/Y vssd1 vssd1 vccd1 vccd1 _07956_/A sky130_fd_sc_hd__a21o_2
XANTENNA__09859__A2 _09858_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07877_ _07642_/A _07876_/A _12668_/A vssd1 vssd1 vccd1 vccd1 _07877_/X sky130_fd_sc_hd__mux2_2
X_09616_ _09338_/A _09338_/B _09336_/Y vssd1 vssd1 vccd1 vccd1 _09631_/A sky130_fd_sc_hd__o21ai_2
X_06828_ _07252_/B vssd1 vssd1 vccd1 vccd1 _07223_/A sky130_fd_sc_hd__inv_2
X_09547_ _09380_/A _09380_/B _09378_/X vssd1 vssd1 vccd1 vccd1 _09562_/A sky130_fd_sc_hd__o21ba_2
X_06759_ reg1_val[26] vssd1 vssd1 vccd1 vccd1 _07392_/A sky130_fd_sc_hd__inv_2
XANTENNA__12615__A1 _12614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08493__A _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09478_ reg1_val[15] reg1_val[16] _09493_/S vssd1 vssd1 vccd1 vccd1 _09478_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12091__A2 _12614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout29_A _07447_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08429_ _08806_/B1 wire122/A _10637_/A _08806_/A2 vssd1 vssd1 vccd1 vccd1 _08430_/B
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_11_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13701_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11440_ _11440_/A _11440_/B vssd1 vssd1 vccd1 vccd1 _11441_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_80_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09244__B1 _08704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08598__A2 _10225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09795__A1 fanout39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09795__B2 _08118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11371_ hold289/A _12058_/A _11579_/C _12748_/B1 vssd1 vssd1 vccd1 vccd1 _11371_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_116_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13110_ reg1_val[26] _13136_/A vssd1 vssd1 vccd1 vccd1 _13111_/B sky130_fd_sc_hd__nand2_1
X_10322_ hold238/A _10459_/C _10606_/A2 vssd1 vssd1 vccd1 vccd1 _10323_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13041_ reg1_val[12] _13042_/B vssd1 vssd1 vccd1 vccd1 _13043_/A sky130_fd_sc_hd__or2_1
X_10253_ _10253_/A _10253_/B vssd1 vssd1 vccd1 vccd1 _10255_/B sky130_fd_sc_hd__xor2_1
XANTENNA__10263__A _10263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07558__B1 _08868_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ hold238/A _10606_/A2 _10459_/C _10183_/Y _12533_/B1 vssd1 vssd1 vccd1 vccd1
+ _10184_/X sky130_fd_sc_hd__a311o_1
Xfanout270 _06936_/A vssd1 vssd1 vccd1 vccd1 _06928_/A sky130_fd_sc_hd__buf_8
Xfanout281 _13444_/C1 vssd1 vssd1 vccd1 vccd1 _13568_/A sky130_fd_sc_hd__clkbuf_4
Xfanout292 reg1_val[0] vssd1 vssd1 vccd1 vccd1 _12982_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__08522__A2 _07541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12825_ reg1_val[4] curr_PC[4] _12825_/S vssd1 vssd1 vccd1 vccd1 _12827_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_29_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09483__A0 _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _13129_/A _11688_/B _12799_/A2 vssd1 vssd1 vccd1 vccd1 _12756_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _12094_/A _11707_/B vssd1 vssd1 vccd1 vccd1 _11709_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12687_ _12765_/A _12687_/B vssd1 vssd1 vccd1 vccd1 _12733_/C sky130_fd_sc_hd__xor2_2
XANTENNA__09235__B1 _10235_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11638_ _11638_/A _11802_/B _11638_/C vssd1 vssd1 vccd1 vccd1 _11640_/A sky130_fd_sc_hd__and3_1
XFILLER_0_24_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08589__A2 _13168_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11968__S _12525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13582__A2 _13584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11569_ _06918_/X _11567_/X _11568_/X vssd1 vssd1 vccd1 vccd1 _11569_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__12790__B1 _12799_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11593__B2 _09493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13308_ _13561_/A _13561_/B _13225_/A vssd1 vssd1 vccd1 vccd1 _13565_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_122_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09538__B2 _09839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13334__A2 _13506_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13239_ _13237_/X _13239_/B vssd1 vssd1 vccd1 vccd1 _13540_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__07549__B1 _07545_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11345__A1 _11109_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07013__A2 _06936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07800_ _10239_/A _07800_/B vssd1 vssd1 vccd1 vccd1 _07807_/A sky130_fd_sc_hd__xnor2_1
X_08780_ _08818_/A _08781_/C vssd1 vssd1 vccd1 vccd1 _08791_/B sky130_fd_sc_hd__nand2_1
X_07731_ _07731_/A _07731_/B vssd1 vssd1 vccd1 vccd1 _07732_/B sky130_fd_sc_hd__or2_1
XFILLER_0_79_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07662_ _11047_/A fanout83/X fanout79/X fanout85/X vssd1 vssd1 vccd1 vccd1 _07663_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10856__B1 _10854_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09401_ _09401_/A _09401_/B vssd1 vssd1 vccd1 vccd1 _09402_/B sky130_fd_sc_hd__xnor2_1
X_07593_ _07594_/B _09254_/D _09254_/C vssd1 vssd1 vccd1 vccd1 _10787_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_62_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11732__A _11732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09332_ _10104_/A _07643_/B fanout13/X _09955_/A vssd1 vssd1 vccd1 vccd1 _09333_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12073__A2 _12164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06826__A _06928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09263_ _09264_/A _09264_/B vssd1 vssd1 vccd1 vccd1 _09263_/X sky130_fd_sc_hd__and2b_1
XANTENNA_fanout233_A _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08214_ _08214_/A _08214_/B vssd1 vssd1 vccd1 vccd1 _08258_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_62_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09194_ _07952_/A _07952_/B _07950_/X vssd1 vssd1 vccd1 vccd1 _09195_/B sky130_fd_sc_hd__a21oi_2
X_08145_ _11286_/A _08145_/B vssd1 vssd1 vccd1 vccd1 _08172_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09777__A1 _07175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11033__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09777__B2 _08933_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10387__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08076_ _08080_/A _08080_/B vssd1 vssd1 vccd1 vccd1 _08076_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07027_ reg2_val[0] _07110_/A vssd1 vssd1 vccd1 vccd1 _07027_/X sky130_fd_sc_hd__and2_1
XFILLER_0_101_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12533__B1 _12533_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ _09044_/B _09033_/A _09033_/B _08785_/X _08760_/Y vssd1 vssd1 vccd1 vccd1
+ _09041_/B sky130_fd_sc_hd__a32o_2
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ _07929_/A _07929_/B vssd1 vssd1 vccd1 vccd1 _07930_/B sky130_fd_sc_hd__or2_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__A2 _11802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10940_ _10941_/A _10941_/B vssd1 vssd1 vccd1 vccd1 _10940_/Y sky130_fd_sc_hd__nand2_1
X_10871_ _10870_/A _10870_/B _10870_/Y _09507_/X vssd1 vssd1 vccd1 vccd1 _10897_/A
+ sky130_fd_sc_hd__a211o_1
X_12610_ _12666_/A _12610_/B vssd1 vssd1 vccd1 vccd1 _12612_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08268__A1 _08821_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08268__B2 _08821_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13590_ hold233/A _13599_/D _13589_/X _13584_/B hold140/X vssd1 vssd1 vccd1 vccd1
+ hold141/A sky130_fd_sc_hd__a32o_1
XFILLER_0_66_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10075__A1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10075__B2 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12541_ _09429_/X _12512_/X _12513_/Y _12517_/X _12540_/X vssd1 vssd1 vccd1 vccd1
+ _12541_/X sky130_fd_sc_hd__o311a_1
XANTENNA__11811__A2 _07891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12472_ _12452_/A _12709_/A2 _09515_/Y _06831_/B _12471_/Y vssd1 vssd1 vccd1 vccd1
+ _12472_/X sky130_fd_sc_hd__a221o_1
XANTENNA__08951__A _08951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11423_ _11423_/A _11825_/A vssd1 vssd1 vccd1 vccd1 _11424_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_21_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_9 instruction[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11354_ _11958_/A _11354_/B vssd1 vssd1 vccd1 vccd1 _11354_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07243__A2 _08866_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08440__A1 _08868_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08440__B2 _10522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10305_ _10201_/X _10727_/A _10304_/Y vssd1 vssd1 vccd1 vccd1 _10305_/Y sky130_fd_sc_hd__a21oi_1
X_11285_ _11708_/A _11285_/B _11285_/C vssd1 vssd1 vccd1 vccd1 _11286_/C sky130_fd_sc_hd__nand3_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13024_ reg1_val[9] _13025_/B vssd1 vssd1 vccd1 vccd1 _13031_/B sky130_fd_sc_hd__or2_1
X_10236_ _10236_/A _10236_/B vssd1 vssd1 vccd1 vccd1 _10241_/A sky130_fd_sc_hd__xnor2_1
X_10167_ reg1_val[4] curr_PC[4] vssd1 vssd1 vccd1 vccd1 _10167_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_max_cap78_A _07526_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10098_ _10099_/A _10099_/B vssd1 vssd1 vccd1 vccd1 _10098_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_89_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12648__A _12648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12808_ _12809_/A _12809_/B vssd1 vssd1 vccd1 vccd1 _12816_/B sky130_fd_sc_hd__or2_1
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12739_ _12740_/A _12739_/B vssd1 vssd1 vccd1 vccd1 _12739_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13555__A2 _13555_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08580__B _08580_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08431__A1 _08821_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08431__B2 _08821_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09950_ _09950_/A _09950_/B vssd1 vssd1 vccd1 vccd1 _09951_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_110_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08901_ _08901_/A _08901_/B vssd1 vssd1 vccd1 vccd1 _08911_/A sky130_fd_sc_hd__xor2_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _09881_/A _10726_/A _10726_/B _09656_/C vssd1 vssd1 vccd1 vccd1 _10044_/A
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08195__B1 _11638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08734__A2 _10522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ _10542_/A _08832_/B vssd1 vssd1 vccd1 vccd1 _08862_/A sky130_fd_sc_hd__xnor2_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10631__A _10631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07416__S _12420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08763_ _08764_/A _08764_/B vssd1 vssd1 vccd1 vccd1 _08763_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07714_ _07714_/A _07714_/B vssd1 vssd1 vccd1 vccd1 _07715_/B sky130_fd_sc_hd__nand2_1
X_08694_ _08694_/A _08694_/B vssd1 vssd1 vccd1 vccd1 _08724_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__13491__B2 _13542_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07645_ _07644_/C _07644_/B _07869_/A vssd1 vssd1 vccd1 vccd1 _07646_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07576_ _11076_/A _10934_/A _07575_/X vssd1 vssd1 vccd1 vccd1 _07576_/Y sky130_fd_sc_hd__a21oi_1
X_09315_ _07961_/X _09201_/X _09202_/X vssd1 vssd1 vccd1 vccd1 _09315_/X sky130_fd_sc_hd__a21o_1
XANTENNA__11254__B1 _12657_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10078__A _10078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09246_ _09246_/A _09246_/B vssd1 vssd1 vccd1 vccd1 _09248_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09177_ _09228_/A _09177_/B vssd1 vssd1 vccd1 vccd1 _09179_/C sky130_fd_sc_hd__nand2_1
XANTENNA__13546__A2 _13555_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08128_ _09951_/A _08128_/B vssd1 vssd1 vccd1 vccd1 _08129_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__07225__A2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08422__A1 _08866_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08422__B2 _08950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08059_ _08821_/B2 _11732_/A _10814_/A1 _08821_/A1 vssd1 vssd1 vccd1 vccd1 _08060_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout96_A _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11070_ _10914_/A _10914_/B _10916_/X vssd1 vssd1 vccd1 vccd1 _11084_/A sky130_fd_sc_hd__a21oi_1
X_10021_ _10458_/S _10020_/X _09537_/B vssd1 vssd1 vccd1 vccd1 _10022_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_101_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09107__A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08011__A _10263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11972_ hold203/A _11972_/B vssd1 vssd1 vccd1 vccd1 _12148_/C sky130_fd_sc_hd__or2_1
X_13711_ _13736_/CLK _13711_/D vssd1 vssd1 vccd1 vccd1 hold287/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10923_ _11913_/A _10923_/B vssd1 vssd1 vccd1 vccd1 _10925_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11493__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13642_ _13649_/CLK hold190/X vssd1 vssd1 vccd1 vccd1 _13642_/Q sky130_fd_sc_hd__dfxtp_1
X_10854_ _10573_/X _10721_/Y _10722_/Y vssd1 vssd1 vccd1 vccd1 _10854_/Y sky130_fd_sc_hd__a21oi_2
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13573_ _13605_/A hold250/X vssd1 vssd1 vccd1 vccd1 _13732_/D sky130_fd_sc_hd__and2_1
X_10785_ _10538_/A fanout10/X fanout5/X _08778_/B vssd1 vssd1 vccd1 vccd1 _10786_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12524_ _12524_/A _12524_/B vssd1 vssd1 vccd1 vccd1 _12524_/Y sky130_fd_sc_hd__xnor2_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08681__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12455_ _09082_/A _12454_/X _12781_/A vssd1 vssd1 vccd1 vccd1 _12455_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__06913__B _07110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11406_ _11521_/A _11521_/B vssd1 vssd1 vccd1 vccd1 _11522_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12386_ reg1_val[24] curr_PC[24] vssd1 vssd1 vccd1 vccd1 _12387_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11337_ _11337_/A _11337_/B vssd1 vssd1 vccd1 vccd1 _11340_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__10771__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11268_ _12372_/A _11600_/A vssd1 vssd1 vccd1 vccd1 _11348_/B sky130_fd_sc_hd__or2_1
X_13007_ _13007_/A _13007_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[5] sky130_fd_sc_hd__xor2_4
X_10219_ _10219_/A _10219_/B vssd1 vssd1 vccd1 vccd1 _10279_/A sky130_fd_sc_hd__xor2_4
X_11199_ _11326_/C _11197_/Y _11075_/Y _11079_/A vssd1 vssd1 vccd1 vccd1 _11200_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11720__A1 _12557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11720__B2 _12557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07152__A1 _13748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07430_ reg1_val[18] _07634_/B _07435_/B vssd1 vssd1 vccd1 vccd1 _11884_/A sky130_fd_sc_hd__or3_1
XFILLER_0_9_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10039__A1 _11866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07361_ _12253_/A _07368_/B vssd1 vssd1 vccd1 vccd1 _07361_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_128_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09100_ _07954_/A _07954_/B _07955_/Y vssd1 vssd1 vccd1 vccd1 _09200_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_128_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07292_ _13015_/A reg1_val[8] _07320_/C vssd1 vssd1 vccd1 vccd1 _10750_/A sky130_fd_sc_hd__or3_2
XFILLER_0_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09031_ _09031_/A _09031_/B vssd1 vssd1 vccd1 vccd1 _11233_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_60_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold301 hold301/A vssd1 vssd1 vccd1 vccd1 hold301/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12841__A _13010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07935__A _09591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09933_ _09932_/B _09932_/C _09932_/A vssd1 vssd1 vccd1 vccd1 _09934_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__08707__A2 wire122/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11457__A _11458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09904__A1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09904__B2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09864_ _07022_/Y _09703_/C _12515_/S vssd1 vssd1 vccd1 vccd1 _09864_/X sky130_fd_sc_hd__a21o_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08815_ _08815_/A _08815_/B vssd1 vssd1 vccd1 vccd1 _08843_/A sky130_fd_sc_hd__xnor2_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ fanout39/X _07471_/Y _07478_/Y _08118_/B vssd1 vssd1 vccd1 vccd1 _09796_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_84_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08746_ _08746_/A _08746_/B vssd1 vssd1 vccd1 vccd1 _08753_/B sky130_fd_sc_hd__xnor2_1
X_08677_ _08677_/A _08677_/B vssd1 vssd1 vccd1 vccd1 _08701_/B sky130_fd_sc_hd__xor2_2
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07628_ _07628_/A _07628_/B vssd1 vssd1 vccd1 vccd1 _07630_/B sky130_fd_sc_hd__xnor2_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07559_ _12094_/A _07559_/B vssd1 vssd1 vccd1 vccd1 _07563_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11920__A _11920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10570_ _10571_/A _10571_/B vssd1 vssd1 vccd1 vccd1 _10570_/X sky130_fd_sc_hd__and2_1
XFILLER_0_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09229_ _09230_/B _09230_/A vssd1 vssd1 vccd1 vccd1 _09229_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_16_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12240_ _12710_/B2 _10879_/A _12235_/X _12239_/X vssd1 vssd1 vccd1 vccd1 _12241_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_252 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12171_ _12260_/A _12260_/B vssd1 vssd1 vccd1 vccd1 _12173_/C sky130_fd_sc_hd__xnor2_1
X_11122_ _11122_/A _11122_/B vssd1 vssd1 vccd1 vccd1 _11122_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_102_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11053_ _11913_/A _11053_/B vssd1 vssd1 vccd1 vccd1 _11061_/A sky130_fd_sc_hd__xor2_1
X_10004_ _09678_/X _09688_/X _10004_/S vssd1 vssd1 vccd1 vccd1 _10004_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08676__A _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11955_ _11955_/A _11955_/B _11955_/C vssd1 vssd1 vccd1 vccd1 _11955_/X sky130_fd_sc_hd__or3_1
XANTENNA__08331__B1 _11638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08395__B _08395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10906_ _07526_/Y fanout16/X fanout12/X _11309_/A vssd1 vssd1 vccd1 vccd1 _10907_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11886_ _06893_/B _09515_/Y _11586_/B _06891_/Y _11885_/X vssd1 vssd1 vccd1 vccd1
+ _11886_/X sky130_fd_sc_hd__a221o_1
X_13625_ _13725_/CLK _13625_/D vssd1 vssd1 vccd1 vccd1 hold126/A sky130_fd_sc_hd__dfxtp_1
X_10837_ _10669_/A _10669_/B _10667_/X vssd1 vssd1 vccd1 vccd1 _10840_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13556_ _13591_/A _13556_/B vssd1 vssd1 vccd1 vccd1 _13728_/D sky130_fd_sc_hd__and2_1
XANTENNA__09831__B1 _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10768_ _10713_/A _10713_/B _10714_/Y vssd1 vssd1 vccd1 vccd1 _10849_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12507_ _12363_/A _12436_/Y _12438_/B vssd1 vssd1 vccd1 vccd1 _12507_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_42_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13487_ _13539_/A _13487_/B vssd1 vssd1 vccd1 vccd1 _13713_/D sky130_fd_sc_hd__and2_1
XFILLER_0_125_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10699_ _10699_/A _10699_/B vssd1 vssd1 vccd1 vccd1 _10701_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_23_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12438_ _12436_/Y _12438_/B vssd1 vssd1 vccd1 vccd1 _12570_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_2_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12369_ _12369_/A _12369_/B vssd1 vssd1 vccd1 vccd1 _12369_/X sky130_fd_sc_hd__and2_1
XFILLER_0_10_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11277__A _12417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06930_ reg2_val[13] _06980_/B _06928_/X vssd1 vssd1 vccd1 vccd1 _07523_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__09362__A2 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06861_ reg1_val[22] _07203_/A vssd1 vssd1 vccd1 vccd1 _06863_/A sky130_fd_sc_hd__nand2_1
X_08600_ _08600_/A _08600_/B vssd1 vssd1 vccd1 vccd1 _08647_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13492__A _13543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09580_ _07238_/X _10536_/A2 fanout6/X _07239_/Y vssd1 vssd1 vccd1 vccd1 _09581_/B
+ sky130_fd_sc_hd__a22o_1
X_06792_ _13135_/A _07398_/B vssd1 vssd1 vccd1 vccd1 _06794_/A sky130_fd_sc_hd__or2_2
XANTENNA__08586__A _09659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08531_ _08532_/A _08532_/B vssd1 vssd1 vccd1 vccd1 _08531_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08462_ _08460_/A _08460_/B _08461_/Y vssd1 vssd1 vccd1 vccd1 _08514_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__08873__A1 _09674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08873__B2 _08873_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07413_ _07414_/A _07414_/B _07414_/C _07414_/D vssd1 vssd1 vccd1 vccd1 _07422_/A
+ sky130_fd_sc_hd__a22o_1
X_08393_ _08873_/B2 fanout24/X _08486_/B _13149_/A vssd1 vssd1 vccd1 vccd1 _08394_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_57_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout146_A _08746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07344_ _07476_/B _07186_/B _07363_/B vssd1 vssd1 vccd1 vccd1 _08907_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07275_ _10095_/A _07285_/B vssd1 vssd1 vccd1 vccd1 _07275_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_72_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09014_ _10306_/C _10160_/B _10160_/C _10445_/A vssd1 vssd1 vccd1 vccd1 _09018_/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_115_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13382__B1 _13207_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold120 hold120/A vssd1 vssd1 vccd1 vccd1 hold120/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 hold131/A vssd1 vssd1 vccd1 vccd1 hold131/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 hold142/A vssd1 vssd1 vccd1 vccd1 hold142/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 hold153/A vssd1 vssd1 vccd1 vccd1 hold153/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 hold164/A vssd1 vssd1 vccd1 vccd1 hold164/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 hold175/A vssd1 vssd1 vccd1 vccd1 hold175/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold186 hold186/A vssd1 vssd1 vccd1 vccd1 hold186/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold197 hold197/A vssd1 vssd1 vccd1 vccd1 hold197/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11187__A _11731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09916_ _09765_/A _09765_/B _09762_/Y vssd1 vssd1 vccd1 vccd1 _09919_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__11145__C1 _11123_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09847_ _09469_/X _09494_/X _10004_/S vssd1 vssd1 vccd1 vccd1 _09847_/X sky130_fd_sc_hd__mux2_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07364__A1 _07363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09778_ _09948_/A _09778_/B vssd1 vssd1 vccd1 vccd1 _09780_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__13437__A1 _12417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout59_A _10522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08729_ _08729_/A _08729_/B vssd1 vssd1 vccd1 vccd1 _08758_/A sky130_fd_sc_hd__nor2_2
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _11633_/A _11633_/B _11641_/X vssd1 vssd1 vccd1 vccd1 _11751_/A sky130_fd_sc_hd__o21ba_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12660__A2 _10010_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10671__A1 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _11562_/B _09048_/B _11562_/A vssd1 vssd1 vccd1 vccd1 _11672_/B sky130_fd_sc_hd__a21o_1
XANTENNA__10671__B2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13410_ hold92/X _13416_/A2 _13420_/B1 hold132/X _13383_/A vssd1 vssd1 vccd1 vccd1
+ hold133/A sky130_fd_sc_hd__o221a_1
XFILLER_0_36_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10622_ _12759_/A1 _10596_/Y _10603_/X _10321_/X _10621_/X vssd1 vssd1 vccd1 vccd1
+ _10622_/X sky130_fd_sc_hd__a221o_1
XANTENNA__06744__A _13141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13341_ _13359_/A hold210/X vssd1 vssd1 vccd1 vccd1 hold211/A sky130_fd_sc_hd__and2_1
XANTENNA__11620__B1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10553_ _10552_/B _10552_/C _10552_/A vssd1 vssd1 vccd1 vccd1 _10554_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__10266__A _10266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13272_ hold283/X hold78/X vssd1 vssd1 vccd1 vccd1 _13273_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_122_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10484_ _10429_/A _10429_/B _10427_/X vssd1 vssd1 vccd1 vccd1 _10575_/A sky130_fd_sc_hd__a21oi_4
X_12223_ _12142_/A _12142_/B _12140_/B vssd1 vssd1 vccd1 vccd1 _12224_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_122_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12154_ _12759_/A1 _11001_/X _12143_/B _12537_/B2 _12153_/X vssd1 vssd1 vccd1 vccd1
+ _12154_/X sky130_fd_sc_hd__a221o_1
X_11105_ _11105_/A _11105_/B vssd1 vssd1 vccd1 vccd1 _11342_/A sky130_fd_sc_hd__or2_2
X_12085_ _12085_/A _12085_/B vssd1 vssd1 vccd1 vccd1 _12086_/B sky130_fd_sc_hd__or2_1
X_11036_ _11719_/A _11036_/B vssd1 vssd1 vccd1 vccd1 _11038_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11825__A _11825_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12987_ _12987_/A _12987_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[1] sky130_fd_sc_hd__xnor2_4
XANTENNA__07107__A1 _07135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08304__B1 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11938_ _11938_/A _11938_/B vssd1 vssd1 vccd1 vccd1 _11940_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11869_ _12738_/S _11868_/X _11867_/X vssd1 vssd1 vccd1 vccd1 _11869_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_27_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13608_ _13739_/CLK _13608_/D vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13539_ _13539_/A _13539_/B vssd1 vssd1 vccd1 vccd1 _13724_/D sky130_fd_sc_hd__and2_1
XANTENNA__08083__A2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07060_ _13129_/A _09146_/A vssd1 vssd1 vccd1 vccd1 _07060_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_70_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12167__A1 _12557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13364__B1 _13555_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12167__B2 _07597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07962_ _07962_/A _07962_/B vssd1 vssd1 vccd1 vccd1 _09318_/A sky130_fd_sc_hd__xnor2_4
X_09701_ _09701_/A _09701_/B vssd1 vssd1 vccd1 vccd1 _09703_/D sky130_fd_sc_hd__nand2_1
X_06913_ reg2_val[15] _07110_/A vssd1 vssd1 vccd1 vccd1 _06913_/X sky130_fd_sc_hd__and2_1
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07893_ _07892_/A _07892_/B _08328_/B2 vssd1 vssd1 vccd1 vccd1 _07895_/B sky130_fd_sc_hd__a21o_1
X_09632_ _09633_/A _09633_/B vssd1 vssd1 vccd1 vccd1 _09634_/A sky130_fd_sc_hd__and2_1
X_06844_ _06842_/Y _06872_/B1 _06873_/B1 reg2_val[24] vssd1 vssd1 vccd1 vccd1 _07252_/D
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09563_ _09369_/A _09369_/B _09368_/A vssd1 vssd1 vccd1 vccd1 _09568_/A sky130_fd_sc_hd__a21o_1
X_06775_ instruction[3] _06775_/B _07123_/A vssd1 vssd1 vccd1 vccd1 is_store sky130_fd_sc_hd__and3_4
XFILLER_0_78_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout263_A _13082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08514_ _08514_/A _08514_/B vssd1 vssd1 vccd1 vccd1 _08569_/B sky130_fd_sc_hd__xor2_2
X_09494_ _09492_/X _09493_/X _09688_/S vssd1 vssd1 vccd1 vccd1 _09494_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08445_ _08866_/A2 fanout75/X _08704_/B _09216_/B2 vssd1 vssd1 vccd1 vccd1 _08446_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08376_ _08418_/A _08418_/B vssd1 vssd1 vccd1 vccd1 _08379_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_46_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07327_ _11126_/A _07328_/B _07328_/C _07328_/D vssd1 vssd1 vccd1 vccd1 _07462_/B
+ sky130_fd_sc_hd__nor4_2
XANTENNA__11602__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08074__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07258_ fanout51/X _08907_/A fanout44/X _08328_/B2 vssd1 vssd1 vccd1 vccd1 _07259_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07821__A2 _10522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12158__A1 _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07189_ _07192_/A _07192_/B vssd1 vssd1 vccd1 vccd1 _07189_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09574__A2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11348__C _11600_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11669__B1 _12163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12910_ _12956_/A _12910_/B vssd1 vssd1 vccd1 vccd1 _12912_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__12330__B2 _12421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12841_ _13010_/B _12841_/B vssd1 vssd1 vccd1 vccd1 _12842_/B sky130_fd_sc_hd__or2_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _12773_/A _12773_/B vssd1 vssd1 vccd1 vccd1 _12772_/Y sky130_fd_sc_hd__nor2_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11723_ _11724_/A _11724_/B vssd1 vssd1 vccd1 vccd1 _11725_/A sky130_fd_sc_hd__nor2_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11654_ _11654_/A _11654_/B vssd1 vssd1 vccd1 vccd1 _11657_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout70 _07548_/X vssd1 vssd1 vccd1 vccd1 fanout70/X sky130_fd_sc_hd__buf_8
X_10605_ _10606_/A2 _10882_/C hold180/A vssd1 vssd1 vccd1 vccd1 _10605_/Y sky130_fd_sc_hd__a21oi_1
Xfanout92 _11514_/A vssd1 vssd1 vccd1 vccd1 _12421_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_107_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08065__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11585_ _11585_/A _12235_/C vssd1 vssd1 vccd1 vccd1 _11585_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_51_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10947__A2 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13324_ hold243/A _13463_/B2 _13450_/B hold226/X vssd1 vssd1 vccd1 vccd1 hold227/A
+ sky130_fd_sc_hd__a22o_1
X_10536_ _10536_/A1 _10536_/A2 fanout6/X _10536_/B2 vssd1 vssd1 vccd1 vccd1 _10537_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09708__A2_N _12235_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13346__B1 _13506_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13255_ hold57/X hold271/X vssd1 vssd1 vccd1 vccd1 _13255_/X sky130_fd_sc_hd__and2b_1
X_10467_ _07557_/A _11793_/B _10464_/Y _10465_/X _10466_/X vssd1 vssd1 vccd1 vccd1
+ _10467_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_110_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12206_ _12207_/A _12440_/A vssd1 vssd1 vccd1 vccd1 _12368_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_103_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13186_ _11997_/A _13194_/A2 hold135/X _13539_/A vssd1 vssd1 vccd1 vccd1 _13629_/D
+ sky130_fd_sc_hd__o211a_1
X_10398_ _10398_/A _10398_/B vssd1 vssd1 vccd1 vccd1 _10415_/A sky130_fd_sc_hd__nor2_2
XANTENNA__07576__A1 _11076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12137_ _12136_/A _12136_/B _09507_/X vssd1 vssd1 vccd1 vccd1 _12137_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_20_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12068_ _12040_/Y _12041_/X _12043_/Y _10866_/B _12067_/Y vssd1 vssd1 vccd1 vccd1
+ _12068_/X sky130_fd_sc_hd__o221a_1
X_11019_ curr_PC[9] _11020_/C curr_PC[10] vssd1 vssd1 vccd1 vccd1 _11019_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07879__A2 _07643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10635__A1 _07455_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10635__B2 wire122/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08230_ _08240_/B _08240_/A vssd1 vssd1 vccd1 vccd1 _08230_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_7_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08161_ _08159_/B _08239_/B _08157_/Y vssd1 vssd1 vccd1 vccd1 _08169_/A sky130_fd_sc_hd__a21o_1
XANTENNA__08056__A2 fanout39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07112_ _13748_/A _13744_/A _09516_/A vssd1 vssd1 vccd1 vccd1 _09524_/B sky130_fd_sc_hd__and3_1
X_08092_ _08092_/A _08092_/B vssd1 vssd1 vccd1 vccd1 _08096_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07043_ _06939_/Y _07042_/X _11356_/A vssd1 vssd1 vccd1 vccd1 _07043_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_113_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08994_ _08167_/X _08994_/B vssd1 vssd1 vccd1 vccd1 _09092_/A sky130_fd_sc_hd__nand2b_1
X_07945_ _07945_/A _07945_/B vssd1 vssd1 vccd1 vccd1 _07958_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06790__A2 _06906_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07876_ _07876_/A _11823_/A vssd1 vssd1 vccd1 vccd1 _07876_/Y sky130_fd_sc_hd__nor2_1
X_09615_ _09812_/B _09615_/B vssd1 vssd1 vccd1 vccd1 _09633_/A sky130_fd_sc_hd__nor2_1
X_06827_ _06826_/Y _06872_/B1 _07110_/A reg2_val[25] vssd1 vssd1 vccd1 vccd1 _07252_/B
+ sky130_fd_sc_hd__a2bb2o_4
X_09546_ _09419_/A _09419_/B _09420_/Y vssd1 vssd1 vccd1 vccd1 _09649_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_92_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06758_ reg1_val[24] vssd1 vssd1 vccd1 vccd1 _07410_/A sky130_fd_sc_hd__inv_2
XANTENNA__12615__A2 _12764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09477_ reg1_val[14] reg1_val[17] _09493_/S vssd1 vssd1 vccd1 vccd1 _09477_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08428_ _08503_/A _08503_/B _08421_/Y vssd1 vssd1 vccd1 vccd1 _08451_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_19_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09244__A1 _10814_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08359_ _08411_/A _08411_/B _08303_/Y vssd1 vssd1 vccd1 vccd1 _08364_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09244__B2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09795__A2 _07471_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11370_ _11252_/B _11579_/C hold289/A vssd1 vssd1 vccd1 vccd1 _11370_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13328__B1 _13506_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10321_ _12648_/A _12760_/A1 _12537_/B2 vssd1 vssd1 vccd1 vccd1 _10321_/X sky130_fd_sc_hd__a21o_1
X_13040_ _13045_/B _13040_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[11] sky130_fd_sc_hd__and2_4
X_10252_ _10252_/A _10252_/B vssd1 vssd1 vccd1 vccd1 _10253_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07558__A1 _07491_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07558__B2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10183_ _10606_/A2 _10459_/C hold238/A vssd1 vssd1 vccd1 vccd1 _10183_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__08949__A _09659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout260 _07155_/X vssd1 vssd1 vccd1 vccd1 _07572_/S sky130_fd_sc_hd__clkbuf_8
Xfanout271 _06776_/X vssd1 vssd1 vccd1 vccd1 _06936_/A sky130_fd_sc_hd__buf_4
Xfanout282 _06764_/Y vssd1 vssd1 vccd1 vccd1 _13444_/C1 sky130_fd_sc_hd__buf_4
Xfanout293 _11958_/A vssd1 vssd1 vccd1 vccd1 _11463_/A sky130_fd_sc_hd__buf_4
XFILLER_0_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12824_ _12830_/B _12824_/B vssd1 vssd1 vccd1 vccd1 new_PC[3] sky130_fd_sc_hd__and2_4
XFILLER_0_29_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12755_ _13129_/A _09254_/A _09519_/Y vssd1 vssd1 vccd1 vccd1 _12755_/X sky130_fd_sc_hd__o21a_1
XANTENNA__09483__A1 _13129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06916__B _07544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ fanout20/X _07597_/X _07891_/X fanout18/X vssd1 vssd1 vccd1 vccd1 _11707_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_56_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _12686_/A _12686_/B vssd1 vssd1 vccd1 vccd1 _12687_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09235__A1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11637_ _11637_/A _11637_/B vssd1 vssd1 vccd1 vccd1 _11638_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_24_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09235__B2 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13691__CLK _13701_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12535__A2_N _11688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11568_ _06918_/X _11567_/X _12047_/C1 vssd1 vssd1 vccd1 vccd1 _11568_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_80_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13307_ _13228_/B _13557_/B _13226_/X vssd1 vssd1 vccd1 vccd1 _13561_/B sky130_fd_sc_hd__a21o_1
X_10519_ _10520_/A _10520_/B vssd1 vssd1 vccd1 vccd1 _10521_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11499_ _11646_/A _11499_/B vssd1 vssd1 vccd1 vccd1 _11503_/A sky130_fd_sc_hd__or2_1
XANTENNA__12372__C _12372_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13238_ hold261/X hold134/X vssd1 vssd1 vccd1 vccd1 _13239_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07549__A1 _07541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07549__B2 _11638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07013__A3 _12995_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13169_ hold51/X _13193_/B vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__or2_1
XANTENNA__11285__A _11708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07730_ _07811_/A vssd1 vssd1 vccd1 vccd1 _07733_/A sky130_fd_sc_hd__inv_2
XANTENNA__09171__B1 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10856__A1 _10580_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07661_ _09575_/A _07661_/B vssd1 vssd1 vccd1 vccd1 _07667_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09710__A2 _11587_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09400_ _09401_/A _09401_/B vssd1 vssd1 vccd1 vccd1 _09400_/Y sky130_fd_sc_hd__nand2_1
X_07592_ _10239_/A _07592_/B vssd1 vssd1 vccd1 vccd1 _07601_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08594__A _08746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09331_ _09331_/A vssd1 vssd1 vccd1 vccd1 _09338_/A sky130_fd_sc_hd__inv_2
XANTENNA__11732__B _11825_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10629__A _10981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12073__A3 _12164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06826__B _13029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09262_ _09262_/A _09262_/B vssd1 vssd1 vccd1 vccd1 _09264_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08213_ _08857_/A _08213_/B vssd1 vssd1 vccd1 vccd1 _08258_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_7_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09193_ _09193_/A _09193_/B vssd1 vssd1 vccd1 vccd1 _09195_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_16_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11033__A1 _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08144_ _10637_/A _07541_/X _07545_/Y wire122/A vssd1 vssd1 vccd1 vccd1 _08145_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09777__A2 _12667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11033__B2 _12103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06842__A _06928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08075_ _11286_/A _08075_/B vssd1 vssd1 vccd1 vccd1 _08080_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07026_ _07026_/A _07026_/B vssd1 vssd1 vccd1 vccd1 _09701_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_113_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08737__B1 _09216_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__buf_1
X_08977_ _09028_/A _08974_/A _08974_/B _09031_/A _08975_/Y vssd1 vssd1 vccd1 vccd1
+ _09033_/B sky130_fd_sc_hd__a41o_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13089__A2 _13129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ _07929_/A _07929_/B vssd1 vssd1 vccd1 vccd1 _07930_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12297__B1 _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07392__B _07535_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09162__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07859_ fanout24/X fanout85/X _07522_/Y _08486_/B vssd1 vssd1 vccd1 vccd1 _07860_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10870_ _10870_/A _10870_/B vssd1 vssd1 vccd1 vccd1 _10870_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09529_ _13135_/A _09529_/B vssd1 vssd1 vccd1 vccd1 _09536_/B sky130_fd_sc_hd__nor2_2
XANTENNA__08268__A2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12064__A3 _12235_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10075__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12540_ _12518_/Y _12519_/X _12526_/X _12539_/X vssd1 vssd1 vccd1 vccd1 _12540_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12471_ _07223_/A _12799_/A2 _12657_/B1 reg1_val[25] _12470_/Y vssd1 vssd1 vccd1
+ vccd1 _12471_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_0_108_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07228__B1 _07521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11422_ _12668_/A _11422_/B vssd1 vssd1 vccd1 vccd1 _11424_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11353_ _07094_/D _11235_/B _06943_/B vssd1 vssd1 vccd1 vccd1 _11354_/B sky130_fd_sc_hd__o21a_1
XANTENNA__08440__A2 _10538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10304_ _10201_/X _10727_/A _10730_/B vssd1 vssd1 vccd1 vccd1 _10304_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11269__A1_N _13180_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11284_ _11285_/B _11285_/C _11708_/A vssd1 vssd1 vccd1 vccd1 _11286_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_104_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13023_ _13022_/A _13019_/Y _13021_/B vssd1 vssd1 vccd1 vccd1 _13027_/A sky130_fd_sc_hd__o21a_2
X_10235_ _10235_/A1 fanout10/X fanout5/X _10235_/B2 vssd1 vssd1 vccd1 vccd1 _10236_/B
+ sky130_fd_sc_hd__o22a_1
X_10166_ _10016_/A _10012_/Y _10016_/C vssd1 vssd1 vccd1 vccd1 _10170_/A sky130_fd_sc_hd__o21a_1
X_10097_ _07173_/Y fanout6/X _10096_/Y _10239_/A vssd1 vssd1 vccd1 vccd1 _10099_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13524__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12807_ _12816_/A _12807_/B vssd1 vssd1 vccd1 vccd1 _12809_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11552__B _11552_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10999_ _10999_/A _10999_/B _10999_/C vssd1 vssd1 vccd1 vccd1 _10999_/X sky130_fd_sc_hd__and3_1
XANTENNA__11263__A1 _10730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ _07084_/X _12740_/B _12738_/S vssd1 vssd1 vccd1 vccd1 _12739_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12669_ _12670_/A _12670_/B vssd1 vssd1 vccd1 vccd1 _12671_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11015__A1 _10603_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12212__B1 _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08431__A2 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08900_ _08970_/A _08970_/B vssd1 vssd1 vccd1 vccd1 _08900_/X sky130_fd_sc_hd__and2_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _10342_/A _10041_/B _09879_/X _09877_/X vssd1 vssd1 vccd1 vccd1 dest_val[2]
+ sky130_fd_sc_hd__a31o_4
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10526__B1 _07543_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08195__A1 _07175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08195__B2 _08933_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08831_ _08873_/A2 _08873_/B2 _13149_/A _08891_/B vssd1 vssd1 vccd1 vccd1 _08832_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10631__B _10857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _08762_/A _08762_/B vssd1 vssd1 vccd1 vccd1 _08764_/B sky130_fd_sc_hd__xor2_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09144__B1 _07521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07713_ _07713_/A _07713_/B vssd1 vssd1 vccd1 vccd1 _07719_/A sky130_fd_sc_hd__xnor2_2
X_08693_ _08722_/A _08722_/B _08661_/X vssd1 vssd1 vccd1 vccd1 _08724_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_73_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13491__A2 _13555_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07644_ _07869_/A _07644_/B _07644_/C vssd1 vssd1 vccd1 vccd1 _07870_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09213__A _12421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07575_ _11076_/A _07575_/B _10078_/A vssd1 vssd1 vccd1 vccd1 _07575_/X sky130_fd_sc_hd__and3b_1
X_09314_ _07961_/X _09201_/X _09202_/X vssd1 vssd1 vccd1 vccd1 _09314_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_118_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09245_ _10507_/A _09245_/B vssd1 vssd1 vccd1 vccd1 _09246_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09176_ _09176_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09177_/B sky130_fd_sc_hd__or2_1
X_08127_ _07239_/Y _11922_/A wire101/A _07238_/X vssd1 vssd1 vccd1 vccd1 _08128_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08422__A2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11962__C1 _12047_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08058_ _08068_/A _08068_/B vssd1 vssd1 vccd1 vccd1 _08058_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07009_ reg1_val[3] _07419_/A vssd1 vssd1 vccd1 vccd1 _07010_/B sky130_fd_sc_hd__nand2_2
XANTENNA__11918__A _12666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10517__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09383__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10020_ _11472_/S _10019_/X _09534_/C vssd1 vssd1 vccd1 vccd1 _10020_/X sky130_fd_sc_hd__o21a_1
XANTENNA_fanout89_A _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11971_ _12058_/A _12057_/B hold298/A vssd1 vssd1 vccd1 vccd1 _11971_/X sky130_fd_sc_hd__a21o_1
X_13710_ _13736_/CLK _13710_/D vssd1 vssd1 vccd1 vccd1 hold294/A sky130_fd_sc_hd__dfxtp_2
XFILLER_0_98_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10922_ _12268_/A fanout29/X fanout27/X fanout45/X vssd1 vssd1 vccd1 vccd1 _10923_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11493__A1 _13180_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07697__B1 _13151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11493__B2 _11638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09123__A _10078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13641_ _13708_/CLK _13641_/D vssd1 vssd1 vccd1 vccd1 hold188/A sky130_fd_sc_hd__dfxtp_1
X_10853_ _10853_/A _10853_/B vssd1 vssd1 vccd1 vccd1 _11106_/A sky130_fd_sc_hd__or2_4
XFILLER_0_79_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13572_ hold249/X _13584_/B _13571_/X _13599_/D vssd1 vssd1 vccd1 vccd1 hold250/A
+ sky130_fd_sc_hd__a22o_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10784_ _10962_/B _10784_/B vssd1 vssd1 vccd1 vccd1 _10832_/A sky130_fd_sc_hd__and2b_1
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12993__A1 _12992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12523_ _12521_/Y _12523_/B vssd1 vssd1 vccd1 vccd1 _12524_/B sky130_fd_sc_hd__nand2b_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12484__A _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12454_ _09082_/B _09082_/C _12130_/A vssd1 vssd1 vccd1 vccd1 _12454_/X sky130_fd_sc_hd__o21a_1
XANTENNA__09506__A_N _13744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11405_ _12417_/A _11405_/B vssd1 vssd1 vccd1 vccd1 _11521_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07297__B _07521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12385_ reg1_val[24] curr_PC[24] vssd1 vssd1 vccd1 vccd1 _12385_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07621__B1 _07833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11336_ _11337_/A _11337_/B vssd1 vssd1 vccd1 vccd1 _11449_/B sky130_fd_sc_hd__or2_1
XFILLER_0_120_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06975__A2 _06928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11267_ _12867_/S _11263_/X _11264_/X _11266_/Y vssd1 vssd1 vccd1 vccd1 dest_val[12]
+ sky130_fd_sc_hd__a22o_4
X_13006_ _13004_/Y _13006_/B vssd1 vssd1 vccd1 vccd1 _13007_/B sky130_fd_sc_hd__nand2b_2
XANTENNA__09374__B1 _09949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13170__A1 _07477_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10218_ _10218_/A _10218_/B vssd1 vssd1 vccd1 vccd1 _10219_/B sky130_fd_sc_hd__nor2_2
X_11198_ _11075_/Y _11079_/A _11326_/C _11197_/Y vssd1 vssd1 vccd1 vccd1 _11326_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__11720__A2 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10149_ _10631_/A vssd1 vssd1 vccd1 vccd1 _10155_/A sky130_fd_sc_hd__inv_2
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09126__B1 _10235_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07152__A2 _13744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11282__B _12614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07360_ _07360_/A _07360_/B _07360_/C _07360_/D vssd1 vssd1 vccd1 vccd1 _07368_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07291_ _10542_/A _07291_/B vssd1 vssd1 vccd1 vccd1 _07721_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10907__A _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09030_ _09028_/A _09023_/A _09023_/B _09023_/C _09029_/Y vssd1 vssd1 vccd1 vccd1
+ _09031_/B sky130_fd_sc_hd__a41o_1
XFILLER_0_115_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09932_ _09932_/A _09932_/B _09932_/C vssd1 vssd1 vccd1 vccd1 _09934_/A sky130_fd_sc_hd__and3_1
XFILLER_0_40_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09904__A2 _07478_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09863_ _07024_/Y _09659_/A _07026_/B vssd1 vssd1 vccd1 vccd1 _09865_/B sky130_fd_sc_hd__a21o_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08814_ _08814_/A _08814_/B _08814_/C vssd1 vssd1 vccd1 vccd1 _08976_/A sky130_fd_sc_hd__and3_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _10263_/A _09794_/B vssd1 vssd1 vccd1 vccd1 _09798_/A sky130_fd_sc_hd__xnor2_1
X_08745_ _09674_/S _10538_/A _08778_/B _08873_/B2 vssd1 vssd1 vccd1 vccd1 _08746_/B
+ sky130_fd_sc_hd__o22a_1
X_08676_ _11072_/A _08676_/B vssd1 vssd1 vccd1 vccd1 _08701_/A sky130_fd_sc_hd__xnor2_2
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07627_ _07628_/A _07628_/B vssd1 vssd1 vccd1 vccd1 _07940_/A sky130_fd_sc_hd__nand2_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10089__A _11281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07558_ _07491_/X _08246_/B _08868_/B1 fanout21/X vssd1 vssd1 vccd1 vccd1 _07559_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07489_ _07180_/C _07363_/B _07186_/B _07476_/B vssd1 vssd1 vccd1 vccd1 _07557_/B
+ sky130_fd_sc_hd__a31o_4
XANTENNA__10817__A _12421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10986__B1 _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09228_ _09228_/A _09228_/B vssd1 vssd1 vccd1 vccd1 _09230_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_91_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09159_ _13129_/A _07865_/B _11823_/A _09157_/X vssd1 vssd1 vccd1 vccd1 _12717_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12170_ _12668_/A _12170_/B vssd1 vssd1 vccd1 vccd1 _12260_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11121_ _11463_/A _06955_/Y _07040_/X _11120_/Y vssd1 vssd1 vccd1 vccd1 _11122_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11052_ fanout45/X fanout29/X fanout27/X fanout49/X vssd1 vssd1 vccd1 vccd1 _11053_/B
+ sky130_fd_sc_hd__o22a_1
X_10003_ _09999_/X _10002_/X _11575_/S vssd1 vssd1 vccd1 vccd1 _10003_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08957__A _09950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11954_ _12695_/A _11988_/A _12164_/A vssd1 vssd1 vccd1 vccd1 _11955_/C sky130_fd_sc_hd__and3_1
XANTENNA__12663__B1 _07108_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08331__A1 _07238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08331__B2 _07239_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10905_ _12420_/A _10905_/B vssd1 vssd1 vccd1 vccd1 _10909_/A sky130_fd_sc_hd__xnor2_1
X_11885_ reg1_val[18] _11688_/B _07310_/A _10889_/B vssd1 vssd1 vccd1 vccd1 _11885_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_104_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13624_ _13719_/CLK _13624_/D vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__dfxtp_1
X_10836_ _10703_/A _10703_/B _10701_/X vssd1 vssd1 vccd1 vccd1 _10841_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13555_ hold282/X _13555_/A2 _13554_/X _13563_/B2 vssd1 vssd1 vccd1 vccd1 _13556_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10767_ _11151_/A _11151_/B vssd1 vssd1 vccd1 vccd1 _10900_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10727__A _10727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12506_ _12506_/A _12506_/B vssd1 vssd1 vccd1 vccd1 _12627_/A sky130_fd_sc_hd__or2_2
XFILLER_0_89_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13486_ hold295/X _13555_/A2 _13485_/X _13542_/B2 vssd1 vssd1 vccd1 vccd1 _13487_/B
+ sky130_fd_sc_hd__a22o_1
X_10698_ _10699_/A _10699_/B vssd1 vssd1 vccd1 vccd1 _10798_/B sky130_fd_sc_hd__or2_1
XFILLER_0_35_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12437_ _12437_/A _12437_/B _12437_/C vssd1 vssd1 vccd1 vccd1 _12438_/B sky130_fd_sc_hd__nand3_1
XANTENNA__09595__B1 _08704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12368_ _12368_/A _12368_/B _12368_/C vssd1 vssd1 vccd1 vccd1 _12368_/X sky130_fd_sc_hd__or3_1
XFILLER_0_105_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11319_ _11319_/A _11319_/B _11319_/C vssd1 vssd1 vccd1 vccd1 _11321_/A sky130_fd_sc_hd__and3_1
X_12299_ _12299_/A _12299_/B vssd1 vssd1 vccd1 vccd1 _12299_/X sky130_fd_sc_hd__xor2_1
X_06860_ _06858_/Y _06872_/B1 _06873_/B1 reg2_val[22] vssd1 vssd1 vccd1 vccd1 _07203_/A
+ sky130_fd_sc_hd__a2bb2o_2
XANTENNA__08867__A _09371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06791_ instruction[41] _06936_/A _06789_/B _06778_/X vssd1 vssd1 vccd1 vccd1 _07398_/B
+ sky130_fd_sc_hd__a31o_4
XANTENNA__11293__A _12093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08530_ _09950_/A _08530_/B vssd1 vssd1 vccd1 vccd1 _08532_/B sky130_fd_sc_hd__xnor2_1
X_08461_ _08473_/A _08473_/B vssd1 vssd1 vccd1 vccd1 _08461_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_77_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08873__A2 _08873_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07412_ _12253_/A _07412_/B vssd1 vssd1 vccd1 vccd1 _12329_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08392_ _08391_/A _08455_/A _08397_/A vssd1 vssd1 vccd1 vccd1 _08392_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_45_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07343_ _07414_/A _07414_/B vssd1 vssd1 vccd1 vccd1 _12252_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_128_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10637__A _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07274_ _09948_/A _07274_/B vssd1 vssd1 vccd1 vccd1 _07285_/B sky130_fd_sc_hd__or2_1
XFILLER_0_73_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09013_ _09013_/A _09013_/B vssd1 vssd1 vccd1 vccd1 _10445_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold110 hold110/A vssd1 vssd1 vccd1 vccd1 hold110/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold121 hold121/A vssd1 vssd1 vccd1 vccd1 hold121/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13382__B2 _12982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10196__A1 _12047_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold132 hold132/A vssd1 vssd1 vccd1 vccd1 hold132/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11393__B1 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold143 hold143/A vssd1 vssd1 vccd1 vccd1 hold143/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 hold154/A vssd1 vssd1 vccd1 vccd1 hold154/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 hold165/A vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 hold176/A vssd1 vssd1 vccd1 vccd1 hold176/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold187 hold187/A vssd1 vssd1 vccd1 vccd1 hold187/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 hold198/A vssd1 vssd1 vccd1 vccd1 hold198/X sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ _09776_/A _09775_/B _09773_/X vssd1 vssd1 vccd1 vccd1 _09922_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07384__C _07634_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08010__B1 _08395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09846_ _09842_/X _09845_/X _11575_/S vssd1 vssd1 vccd1 vccd1 _09846_/X sky130_fd_sc_hd__mux2_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _07175_/X _12667_/A _10536_/A2 _08933_/B vssd1 vssd1 vccd1 vccd1 _09778_/B
+ sky130_fd_sc_hd__a22o_1
X_06989_ _07110_/A _06989_/B _13010_/B vssd1 vssd1 vccd1 vccd1 _06989_/X sky130_fd_sc_hd__or3b_2
XANTENNA__13437__A2 _13598_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08728_ _08728_/A _08728_/B vssd1 vssd1 vccd1 vccd1 _08729_/B sky130_fd_sc_hd__nor2_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _08659_/A _08659_/B vssd1 vssd1 vccd1 vccd1 _08692_/A sky130_fd_sc_hd__nor2_2
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _11231_/A _11601_/X _12163_/A _11955_/A vssd1 vssd1 vccd1 vccd1 _11670_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10671__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10621_ _12525_/A _12760_/A1 _10620_/Y _10615_/Y vssd1 vssd1 vccd1 vccd1 _10621_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08077__B1 _08580_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13340_ _13651_/Q _13506_/B2 _13506_/A2 hold209/X vssd1 vssd1 vccd1 vccd1 hold210/A
+ sky130_fd_sc_hd__a22o_1
X_10552_ _10552_/A _10552_/B _10552_/C vssd1 vssd1 vccd1 vccd1 _10554_/B sky130_fd_sc_hd__or3_1
XANTENNA__11620__A1 _12103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11620__B2 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13271_ hold78/X hold283/X vssd1 vssd1 vccd1 vccd1 _13271_/X sky130_fd_sc_hd__and2b_1
X_10483_ _10344_/X _10441_/X _12130_/A vssd1 vssd1 vccd1 vccd1 _10483_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_122_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12222_ _12222_/A _12222_/B vssd1 vssd1 vccd1 vccd1 _12224_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07856__A _10263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10187__A1 _12314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11384__B1 _12867_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12153_ _12136_/A _12709_/A2 _09515_/Y _06876_/A _12152_/Y vssd1 vssd1 vccd1 vccd1
+ _12153_/X sky130_fd_sc_hd__a221o_1
XANTENNA__09329__B1 _07699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11104_ _11104_/A _11104_/B _11104_/C vssd1 vssd1 vccd1 vccd1 _11105_/B sky130_fd_sc_hd__and3_1
X_12084_ _12085_/A _12085_/B vssd1 vssd1 vccd1 vccd1 _12173_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08001__B1 _08704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11035_ _07299_/Y fanout32/X fanout70/X fanout34/X vssd1 vssd1 vccd1 vccd1 _11036_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13428__A2 _06744_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12986_ _12984_/Y _12986_/B vssd1 vssd1 vccd1 vccd1 _12987_/B sky130_fd_sc_hd__nand2b_2
XANTENNA__12636__B1 _12056_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08304__A1 _08873_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08304__B2 _08891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11937_ _11938_/A _11938_/B vssd1 vssd1 vccd1 vccd1 _12029_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_115_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13532__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11868_ _06902_/A _11771_/X _06902_/B vssd1 vssd1 vccd1 vccd1 _11868_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_27_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11560__B _11561_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10819_ _11512_/A _10819_/B vssd1 vssd1 vccd1 vccd1 _10821_/B sky130_fd_sc_hd__xnor2_1
X_13607_ _13742_/CLK _13607_/D vssd1 vssd1 vccd1 vccd1 hold109/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11799_ _11601_/X _11896_/C _12695_/A vssd1 vssd1 vccd1 vccd1 _11862_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_54_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13538_ hold261/X _13555_/A2 _13537_/X _13542_/B2 vssd1 vssd1 vccd1 vccd1 _13539_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13469_ _13469_/A _13469_/B vssd1 vssd1 vccd1 vccd1 _13469_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09457__S _09674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12167__A2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11375__B1 _11587_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07961_ _07962_/A _07962_/B vssd1 vssd1 vccd1 vccd1 _07961_/X sky130_fd_sc_hd__or2_1
XFILLER_0_49_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09700_ _13642_/Q hold188/A _10606_/A2 _12795_/A1 vssd1 vssd1 vccd1 vccd1 _09700_/X
+ sky130_fd_sc_hd__a31o_1
X_06912_ _06912_/A _06912_/B vssd1 vssd1 vccd1 vccd1 _07092_/D sky130_fd_sc_hd__nor2_1
X_07892_ _07892_/A _07892_/B vssd1 vssd1 vccd1 vccd1 _12667_/A sky130_fd_sc_hd__nand2_8
X_09631_ _09631_/A _09631_/B vssd1 vssd1 vccd1 vccd1 _09633_/B sky130_fd_sc_hd__xnor2_1
X_06843_ reg2_val[24] _06873_/B1 _06872_/B1 _06842_/Y vssd1 vssd1 vccd1 vccd1 _07221_/A
+ sky130_fd_sc_hd__o2bb2a_2
X_09562_ _09562_/A _09562_/B vssd1 vssd1 vccd1 vccd1 _09635_/A sky130_fd_sc_hd__xnor2_4
X_06774_ _09524_/A _06775_/B _07123_/A vssd1 vssd1 vccd1 vccd1 is_load sky130_fd_sc_hd__and3_4
X_08513_ _08565_/A _08565_/B _08474_/X vssd1 vssd1 vccd1 vccd1 _08569_/A sky130_fd_sc_hd__a21oi_2
X_09493_ _13015_/A reg1_val[24] _09493_/S vssd1 vssd1 vccd1 vccd1 _09493_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12847__A _13015_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout256_A _12754_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08444_ _08448_/A _08448_/B vssd1 vssd1 vccd1 vccd1 _08449_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_92_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08059__B1 _10814_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08375_ _09659_/B _08375_/B vssd1 vssd1 vccd1 vccd1 _08418_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07326_ reg1_val[14] reg1_val[15] vssd1 vssd1 vccd1 vccd1 _07328_/D sky130_fd_sc_hd__or2_1
XANTENNA__11602__A1 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11602__B2 _12557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07257_ _07594_/B _09254_/D _07255_/X _07251_/Y vssd1 vssd1 vccd1 vccd1 _07257_/X
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_5_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07676__A _10266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07019__D1 _07110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07188_ _07522_/A _07188_/B _07188_/C _07187_/B vssd1 vssd1 vccd1 vccd1 _07193_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09891__A _12092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11669__A1 _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout71_A _07547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12330__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09731__B1 _07455_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09829_ _10435_/A _10435_/B _09827_/X _09828_/X vssd1 vssd1 vccd1 vccd1 _09830_/B
+ sky130_fd_sc_hd__o211a_2
X_12840_ _13010_/B _12841_/B vssd1 vssd1 vccd1 vccd1 _12851_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10892__A2 _11587_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _12773_/A _12773_/B vssd1 vssd1 vccd1 vccd1 _12771_/Y sky130_fd_sc_hd__nand2_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _11722_/A _11722_/B vssd1 vssd1 vccd1 vccd1 _11724_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _11654_/A _11654_/B vssd1 vssd1 vccd1 vccd1 _11758_/A sky130_fd_sc_hd__nand2_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout60 _09266_/X vssd1 vssd1 vccd1 vccd1 _10522_/B sky130_fd_sc_hd__buf_8
Xfanout71 _07547_/X vssd1 vssd1 vccd1 vccd1 _11638_/A sky130_fd_sc_hd__clkbuf_16
X_10604_ hold237/A _10604_/B vssd1 vssd1 vccd1 vccd1 _10882_/C sky130_fd_sc_hd__or2_1
XANTENNA__12397__A2 _09520_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout82 _07522_/Y vssd1 vssd1 vccd1 vccd1 fanout82/X sky130_fd_sc_hd__buf_8
X_11584_ hold195/A _11693_/A2 _11691_/B _12533_/B1 vssd1 vssd1 vccd1 vccd1 _11584_/X
+ sky130_fd_sc_hd__a31o_1
Xfanout93 _11719_/A vssd1 vssd1 vccd1 vccd1 _12417_/A sky130_fd_sc_hd__buf_8
XFILLER_0_24_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13323_ _13459_/A hold244/X vssd1 vssd1 vccd1 vccd1 _13643_/D sky130_fd_sc_hd__and2_1
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10535_ _10360_/A _10360_/B _10358_/X vssd1 vssd1 vccd1 vccd1 _10546_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_24_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13254_ hold289/X hold66/X vssd1 vssd1 vccd1 vccd1 _13513_/B sky130_fd_sc_hd__nand2b_1
X_10466_ _07270_/X _12235_/C _12657_/B1 reg1_val[6] vssd1 vssd1 vccd1 vccd1 _10466_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10724__B _10981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11357__B1 _09507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12205_ _12031_/X _12119_/Y _12121_/B vssd1 vssd1 vccd1 vccd1 _12208_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13185_ hold134/X _13191_/B vssd1 vssd1 vccd1 vccd1 hold135/A sky130_fd_sc_hd__or2_1
X_10397_ _10397_/A _10397_/B vssd1 vssd1 vccd1 vccd1 _10398_/B sky130_fd_sc_hd__nor2_1
X_12136_ _12136_/A _12136_/B vssd1 vssd1 vccd1 vccd1 _12136_/Y sky130_fd_sc_hd__nor2_1
X_12067_ _12760_/A1 _12053_/X _12066_/X _12047_/X vssd1 vssd1 vccd1 vccd1 _12067_/Y
+ sky130_fd_sc_hd__a211oi_4
X_11018_ _10985_/X _10986_/Y _10988_/Y _11866_/A _11017_/X vssd1 vssd1 vccd1 vccd1
+ _11018_/X sky130_fd_sc_hd__a221o_1
XANTENNA__08210__A _08746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12609__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12667__A _12667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12969_ _12979_/A _12960_/B _12964_/A _12964_/B vssd1 vssd1 vccd1 vccd1 _12970_/B
+ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__10635__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08160_ _08160_/A _08160_/B vssd1 vssd1 vccd1 vccd1 _08239_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_55_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11596__B1 _07544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07111_ _13744_/A _09516_/A vssd1 vssd1 vccd1 vccd1 _09514_/B sky130_fd_sc_hd__and2_2
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08091_ _08111_/A _08111_/B _08070_/Y vssd1 vssd1 vccd1 vccd1 _08098_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_43_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10915__A _10915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07042_ _06947_/Y _07041_/X _11237_/A vssd1 vssd1 vccd1 vccd1 _07042_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_30_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13010__B _13010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08993_ _08993_/A _08994_/B vssd1 vssd1 vccd1 vccd1 _08993_/X sky130_fd_sc_hd__and2_1
X_07944_ _07944_/A _07944_/B vssd1 vssd1 vccd1 vccd1 _07945_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07875_ _07617_/A _07617_/B _07615_/Y vssd1 vssd1 vccd1 vccd1 _07882_/A sky130_fd_sc_hd__o21a_1
XANTENNA__08120__A _10239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_2_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09614_ _09812_/A _09613_/C _09613_/A vssd1 vssd1 vccd1 vccd1 _09615_/B sky130_fd_sc_hd__o21a_1
X_06826_ _06928_/B _13029_/B vssd1 vssd1 vccd1 vccd1 _06826_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_97_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09545_ _09424_/A _09424_/B _09422_/X vssd1 vssd1 vccd1 vccd1 _09650_/A sky130_fd_sc_hd__a21oi_4
X_06757_ reg1_val[23] vssd1 vssd1 vccd1 vccd1 _07334_/B sky130_fd_sc_hd__inv_2
X_09476_ _09474_/X _09475_/X _09688_/S vssd1 vssd1 vccd1 vccd1 _09476_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12296__B _12372_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08427_ _08427_/A _08427_/B vssd1 vssd1 vccd1 vccd1 _08503_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09886__A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08358_ _08358_/A _08358_/B vssd1 vssd1 vccd1 vccd1 _08411_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_34_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09244__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11587__B1 _12657_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07309_ _07309_/A _07310_/B vssd1 vssd1 vccd1 vccd1 wire101/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_116_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08289_ _08288_/A _08288_/B _08288_/C vssd1 vssd1 vccd1 vccd1 _08292_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10320_ _10317_/X _10319_/X _10458_/S vssd1 vssd1 vccd1 vccd1 _10320_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_116_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10251_ _10252_/A _10252_/B vssd1 vssd1 vccd1 vccd1 _10251_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07558__A2 _08246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10182_ hold226/A hold243/A _13642_/Q hold188/A vssd1 vssd1 vccd1 vccd1 _10459_/C
+ sky130_fd_sc_hd__or4_2
Xfanout250 _13463_/B2 vssd1 vssd1 vccd1 vccd1 _13506_/B2 sky130_fd_sc_hd__buf_4
XANTENNA__09704__B1 _09520_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout261 _07155_/X vssd1 vssd1 vccd1 vccd1 _07865_/B sky130_fd_sc_hd__buf_4
Xfanout272 _13459_/A vssd1 vssd1 vccd1 vccd1 _13359_/A sky130_fd_sc_hd__clkbuf_4
Xfanout283 _06762_/Y vssd1 vssd1 vccd1 vccd1 _12515_/S sky130_fd_sc_hd__clkbuf_8
Xfanout294 _12578_/A vssd1 vssd1 vccd1 vccd1 _11958_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__11511__B1 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12823_ _12823_/A _12823_/B _12823_/C vssd1 vssd1 vccd1 vccd1 _12824_/B sky130_fd_sc_hd__nand3_1
XANTENNA__12067__A1 _12760_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12754_ _12754_/A _12754_/B _12754_/C vssd1 vssd1 vccd1 vccd1 _12754_/X sky130_fd_sc_hd__and3_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _11913_/A _11705_/B vssd1 vssd1 vccd1 vccd1 _11710_/A sky130_fd_sc_hd__xnor2_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12685_ _12443_/Y _12682_/C _12682_/D _12684_/X vssd1 vssd1 vccd1 vccd1 _12686_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09796__A _10119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11636_ _11825_/A _11636_/B vssd1 vssd1 vccd1 vccd1 _11637_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09235__A2 _10235_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12775__C1 _09429_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11567_ _11958_/A _06923_/X _07044_/X _11566_/Y vssd1 vssd1 vccd1 vccd1 _11567_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_24_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10518_ _10518_/A _10518_/B vssd1 vssd1 vccd1 vccd1 _10520_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12790__A2 _11688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13306_ _13552_/B _13553_/A _13229_/X vssd1 vssd1 vccd1 vccd1 _13557_/B sky130_fd_sc_hd__a21o_1
X_11498_ _11498_/A _11498_/B vssd1 vssd1 vccd1 vccd1 _11499_/B sky130_fd_sc_hd__nor2_1
XANTENNA__12372__D _12372_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13237_ hold134/X hold261/X vssd1 vssd1 vccd1 vccd1 _13237_/X sky130_fd_sc_hd__and2b_1
X_10449_ _10449_/A _10449_/B vssd1 vssd1 vccd1 vccd1 _10449_/X sky130_fd_sc_hd__xor2_1
XANTENNA__07549__A2 _07544_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13168_ _13168_/A1 _13194_/A2 hold63/X _13543_/A vssd1 vssd1 vccd1 vccd1 _13620_/D
+ sky130_fd_sc_hd__o211a_1
X_12119_ _12121_/A vssd1 vssd1 vccd1 vccd1 _12119_/Y sky130_fd_sc_hd__inv_2
X_13099_ reg1_val[24] _13136_/A vssd1 vssd1 vccd1 vccd1 _13101_/A sky130_fd_sc_hd__or2_1
XANTENNA__09171__A1 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09171__B2 _08395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07660_ fanout74/X fanout68/X fanout66/X fanout70/X vssd1 vssd1 vccd1 vccd1 _07661_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09470__S _09493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07591_ _08821_/B2 fanout47/X fanout45/X _08821_/A1 vssd1 vssd1 vccd1 vccd1 _07592_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_87_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09330_ _10050_/A _09330_/B vssd1 vssd1 vccd1 vccd1 _09331_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10629__B _10981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09261_ _09261_/A _09261_/B vssd1 vssd1 vccd1 vccd1 _09262_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_62_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13005__B _13005_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08682__B1 _08868_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08212_ _08806_/A2 _13168_/A1 _07477_/X _08806_/B1 vssd1 vssd1 vccd1 vccd1 _08213_/B
+ sky130_fd_sc_hd__a22o_1
X_09192_ _09192_/A _09192_/B vssd1 vssd1 vccd1 vccd1 _09193_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_28_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08143_ _08150_/A _08150_/B vssd1 vssd1 vccd1 vccd1 _08143_/X sky130_fd_sc_hd__and2b_1
XANTENNA__07237__A1 _09371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08434__B1 _11047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11033__A2 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06842__B _13025_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08074_ _10049_/A2 fanout75/X _08704_/B _09173_/B2 vssd1 vssd1 vccd1 vccd1 _08075_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_70_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07025_ _12985_/A _07025_/B _07025_/C vssd1 vssd1 vccd1 vccd1 _07026_/B sky130_fd_sc_hd__and3_1
XFILLER_0_30_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08737__A1 _08873_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08737__B2 _08891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ _08976_/A _08976_/B vssd1 vssd1 vccd1 vccd1 _09031_/A sky130_fd_sc_hd__nor2_2
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ _07927_/A _07927_/B vssd1 vssd1 vccd1 vccd1 _07929_/B sky130_fd_sc_hd__xor2_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09698__C1 _12760_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09162__A1 _09910_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09162__B2 _09604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07858_ _10266_/A _07858_/B vssd1 vssd1 vccd1 vccd1 _07862_/A sky130_fd_sc_hd__xnor2_1
X_06809_ _06928_/B _13054_/B vssd1 vssd1 vccd1 vccd1 _06809_/Y sky130_fd_sc_hd__nor2_1
X_07789_ _10049_/A2 fanout84/X _08580_/B _09173_/B2 vssd1 vssd1 vccd1 vccd1 _07790_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_39_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09528_ _09527_/X _09528_/B _09528_/C vssd1 vssd1 vccd1 vccd1 _09528_/X sky130_fd_sc_hd__and3b_1
XANTENNA_fanout34_A fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09459_ _11126_/A reg1_val[20] _09463_/S vssd1 vssd1 vccd1 vccd1 _09459_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_66_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11009__C1 _12748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12470_ reg1_val[25] _07252_/B _09519_/Y vssd1 vssd1 vccd1 vccd1 _12470_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11421_ wire101/X fanout16/X fanout12/X _13180_/A1 vssd1 vssd1 vccd1 vccd1 _11422_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11352_ _11352_/A _11352_/B vssd1 vssd1 vccd1 vccd1 _11352_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10303_ _10857_/A _10303_/B vssd1 vssd1 vccd1 vccd1 _10727_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_104_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11283_ _11283_/A _12667_/A vssd1 vssd1 vccd1 vccd1 _11285_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_104_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13022_ _13022_/A _13022_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[8] sky130_fd_sc_hd__xor2_4
X_10234_ _10392_/B _10234_/B vssd1 vssd1 vccd1 vccd1 _10257_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10165_ _10165_/A _10165_/B vssd1 vssd1 vccd1 vccd1 _10165_/X sky130_fd_sc_hd__or2_1
X_10096_ _10096_/A fanout6/X vssd1 vssd1 vccd1 vccd1 _10096_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_88_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12806_ _12806_/A _12806_/B vssd1 vssd1 vccd1 vccd1 _12807_/B sky130_fd_sc_hd__or2_1
XFILLER_0_97_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10998_ _10999_/A _10999_/B _10999_/C vssd1 vssd1 vccd1 vccd1 _10998_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11799__B1 _12695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _06813_/Y _12691_/Y _06815_/B vssd1 vssd1 vccd1 vccd1 _12740_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_45_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12668_ _12668_/A _12668_/B vssd1 vssd1 vccd1 vccd1 _12670_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12212__A1 _12695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11619_ _11619_/A _11619_/B vssd1 vssd1 vccd1 vccd1 _11633_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12599_ _06801_/Y _12709_/A2 _09519_/Y vssd1 vssd1 vccd1 vccd1 _12599_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08195__A2 _07544_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08830_ _08836_/B _08836_/A vssd1 vssd1 vccd1 vccd1 _08830_/Y sky130_fd_sc_hd__nand2b_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10631__C _10981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ _08761_/A _08761_/B vssd1 vssd1 vccd1 vccd1 _08764_/A sky130_fd_sc_hd__xnor2_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07712_ _07710_/A _07710_/B _07965_/A vssd1 vssd1 vccd1 vccd1 _07786_/A sky130_fd_sc_hd__a21bo_1
X_08692_ _08692_/A _08692_/B vssd1 vssd1 vccd1 vccd1 _08722_/B sky130_fd_sc_hd__xor2_4
X_07643_ _09161_/A _07643_/B vssd1 vssd1 vccd1 vccd1 _07869_/A sky130_fd_sc_hd__nand2_1
X_07574_ _10537_/A _07575_/B vssd1 vssd1 vccd1 vccd1 _07577_/B sky130_fd_sc_hd__and2_1
XFILLER_0_48_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09313_ _09313_/A _09313_/B vssd1 vssd1 vccd1 vccd1 _09986_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__11254__A2 _11793_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12855__A _13020_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09244_ _10814_/A1 fanout75/X _08704_/B fanout42/X vssd1 vssd1 vccd1 vccd1 _09245_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10462__B1 _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09175_ _09176_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09228_/A sky130_fd_sc_hd__nand2_2
XANTENNA__10375__A _10522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08126_ _08125_/B _08125_/C _08125_/A vssd1 vssd1 vccd1 vccd1 _08129_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10765__A1 _12825_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08057_ _10119_/A _08057_/B vssd1 vssd1 vccd1 vccd1 _08068_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07008_ reg1_val[3] _07419_/A vssd1 vssd1 vccd1 vccd1 _07008_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10517__A1 wire122/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10517__B2 _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09383__A1 _09910_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09383__B2 _09604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08959_ _08959_/A _08959_/B vssd1 vssd1 vccd1 vccd1 _08960_/B sky130_fd_sc_hd__xnor2_1
X_11970_ hold298/A _12058_/A _12057_/B vssd1 vssd1 vccd1 vccd1 _11970_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__07697__A1 _07347_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10921_ _12253_/A _10921_/B vssd1 vssd1 vccd1 vccd1 _10925_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07697__B2 fanout39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11493__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10852_ _10852_/A _10852_/B _10852_/C vssd1 vssd1 vccd1 vccd1 _10853_/B sky130_fd_sc_hd__and3_1
X_13640_ _13739_/CLK _13640_/D vssd1 vssd1 vccd1 vccd1 hold172/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11372__C _12598_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ _10783_/A _10783_/B _10781_/X vssd1 vssd1 vccd1 vccd1 _10784_/B sky130_fd_sc_hd__or3b_1
X_13571_ hold273/A _13570_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13571_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_39_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ reg1_val[26] curr_PC[26] vssd1 vssd1 vccd1 vccd1 _12523_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_54_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12453_ _12452_/A _12452_/B _12452_/Y _09506_/X vssd1 vssd1 vccd1 vccd1 _12476_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10205__B1 _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11404_ _07282_/X fanout34/X fanout32/X _12087_/A vssd1 vssd1 vccd1 vccd1 _11405_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_34_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12384_ _12305_/Y _12309_/B _12307_/B vssd1 vssd1 vccd1 vccd1 _12388_/A sky130_fd_sc_hd__o21a_1
XANTENNA__11953__B1 _12164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07621__A1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11335_ _11213_/A _11213_/B _11214_/Y vssd1 vssd1 vccd1 vccd1 _11337_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_105_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07621__B2 _10104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06975__A3 _13020_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11266_ _12867_/S _11266_/B vssd1 vssd1 vccd1 vccd1 _11266_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09374__A1 _08271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13005_ reg1_val[5] _13005_/B vssd1 vssd1 vccd1 vccd1 _13006_/B sky130_fd_sc_hd__nand2_1
X_10217_ _10217_/A _10217_/B _10217_/C vssd1 vssd1 vccd1 vccd1 _10218_/B sky130_fd_sc_hd__and3_1
XANTENNA__13170__A2 _13194_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11197_ _07477_/X _11802_/B _11058_/X _11062_/A vssd1 vssd1 vccd1 vccd1 _11197_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10148_ _10148_/A _10148_/B vssd1 vssd1 vccd1 vccd1 _10631_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__09126__A1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09126__B2 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10079_ _10080_/A _10080_/B vssd1 vssd1 vccd1 vccd1 _10081_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_43_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07290_ _10235_/A1 fanout42/X _10235_/B2 fanout40/X vssd1 vssd1 vccd1 vccd1 _07291_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_72_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10747__A1 _12056_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10923__A _11913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09931_ _10542_/A _09931_/B _09931_/C vssd1 vssd1 vccd1 vccd1 _09932_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09862_ hold243/A _09862_/B vssd1 vssd1 vccd1 vccd1 _09862_/Y sky130_fd_sc_hd__xnor2_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08813_ _08815_/A _08815_/B vssd1 vssd1 vccd1 vccd1 _08814_/C sky130_fd_sc_hd__nand2b_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ fanout28/X fanout74/X fanout70/X _08395_/B vssd1 vssd1 vccd1 vccd1 _09794_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08744_ _08744_/A _08744_/B vssd1 vssd1 vccd1 vccd1 _08753_/A sky130_fd_sc_hd__xnor2_1
X_08675_ _09674_/S fanout75/X _08704_/B _08873_/B2 vssd1 vssd1 vccd1 vccd1 _08676_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_95_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07626_ _10119_/A _07626_/B vssd1 vssd1 vccd1 vccd1 _07628_/B sky130_fd_sc_hd__xnor2_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11880__C1 _12533_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07557_ _07557_/A _07557_/B vssd1 vssd1 vccd1 vccd1 _07557_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__07679__A _10263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07488_ _11991_/A _07493_/B _12093_/A vssd1 vssd1 vccd1 vccd1 _07488_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_119_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09227_ _09130_/A _09130_/B _09128_/Y vssd1 vssd1 vccd1 vccd1 _09228_/B sky130_fd_sc_hd__o21a_1
XANTENNA__07398__B _07398_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09158_ _13129_/A _07865_/B _09157_/X vssd1 vssd1 vccd1 vccd1 _09160_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_44_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08109_ _08109_/A _08109_/B vssd1 vssd1 vccd1 vccd1 _08164_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08800__B1 _08868_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09089_ _09089_/A _09318_/B vssd1 vssd1 vccd1 vccd1 _12584_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11120_ _11463_/A _11120_/B vssd1 vssd1 vccd1 vccd1 _11120_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_102_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11051_ _11051_/A _11051_/B vssd1 vssd1 vccd1 vccd1 _11064_/A sky130_fd_sc_hd__or2_1
XANTENNA__13152__A2 _13193_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10002_ _10000_/X _10001_/X _10176_/A vssd1 vssd1 vccd1 vccd1 _10002_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_99_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09134__A _11286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11953_ _12695_/A _11988_/A _12164_/A vssd1 vssd1 vccd1 vccd1 _11955_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__08331__A2 _07544_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10904_ _13180_/A1 fanout15/X fanout31/X wire101/X vssd1 vssd1 vccd1 vccd1 _10905_/B
+ sky130_fd_sc_hd__a22o_1
X_11884_ _11884_/A _11884_/B _12235_/C vssd1 vssd1 vccd1 vccd1 _11884_/X sky130_fd_sc_hd__and3_1
XFILLER_0_86_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13623_ _13719_/CLK _13623_/D vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__dfxtp_1
X_10835_ _10704_/A _10704_/B _10685_/A vssd1 vssd1 vccd1 vccd1 _10845_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13554_ hold255/X _13553_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13554_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_27_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10766_ curr_PC[9] _11020_/C vssd1 vssd1 vccd1 vccd1 _10766_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__10727__B _10727_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12505_ _12505_/A _12505_/B _12505_/C vssd1 vssd1 vccd1 vccd1 _12506_/B sky130_fd_sc_hd__and3_1
X_10697_ _10798_/A _10697_/B vssd1 vssd1 vccd1 vccd1 _10699_/B sky130_fd_sc_hd__nand2_1
X_13485_ hold276/X _13484_/Y hold234/X vssd1 vssd1 vccd1 vccd1 _13485_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_82_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07101__B _13748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12436_ _12437_/A _12437_/B _12437_/C vssd1 vssd1 vccd1 vccd1 _12436_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09595__A1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09595__B2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12367_ _12368_/B _12368_/C vssd1 vssd1 vccd1 vccd1 _12369_/B sky130_fd_sc_hd__nor2_1
X_11318_ _11318_/A _11318_/B vssd1 vssd1 vccd1 vccd1 _11319_/C sky130_fd_sc_hd__xnor2_1
X_12298_ _09066_/Y _12214_/A _12742_/A vssd1 vssd1 vccd1 vccd1 _12299_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08213__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11249_ _11693_/A2 _11366_/B hold214/A vssd1 vssd1 vccd1 vccd1 _11249_/X sky130_fd_sc_hd__a21o_1
XANTENNA__11154__A1 _07472_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06790_ _06747_/Y _06906_/B1 _06778_/X vssd1 vssd1 vccd1 vccd1 _06790_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_54_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_7_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08460_ _08460_/A _08460_/B vssd1 vssd1 vccd1 vccd1 _08473_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_77_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07411_ _07414_/C _07414_/D vssd1 vssd1 vccd1 vccd1 _07412_/B sky130_fd_sc_hd__and2_1
X_08391_ _08391_/A _08455_/A vssd1 vssd1 vccd1 vccd1 _08397_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_92_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07342_ _07414_/A _07414_/B vssd1 vssd1 vccd1 vccd1 _11603_/A sky130_fd_sc_hd__and2_4
XANTENNA__09283__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10637__B _12764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07273_ _09948_/A _07274_/B vssd1 vssd1 vccd1 vccd1 _10366_/A sky130_fd_sc_hd__nand2_1
X_09012_ _09012_/A _09012_/B vssd1 vssd1 vccd1 vccd1 _10306_/C sky130_fd_sc_hd__xor2_2
XFILLER_0_73_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07011__B _07110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11917__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold100 hold100/A vssd1 vssd1 vccd1 vccd1 hold100/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13382__A2 _07118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold111 hold111/A vssd1 vssd1 vccd1 vccd1 hold111/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold122 hold122/A vssd1 vssd1 vccd1 vccd1 hold122/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 hold133/A vssd1 vssd1 vccd1 vccd1 hold133/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11393__A1 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11393__B2 _12557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold144 hold144/A vssd1 vssd1 vccd1 vccd1 hold144/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 hold155/A vssd1 vssd1 vccd1 vccd1 hold155/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08123__A _09949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold166 hold166/A vssd1 vssd1 vccd1 vccd1 hold166/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 hold212/X vssd1 vssd1 vccd1 vccd1 hold177/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold188 hold188/A vssd1 vssd1 vccd1 vccd1 hold188/X sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ _09914_/A _09914_/B vssd1 vssd1 vccd1 vccd1 _09966_/A sky130_fd_sc_hd__xnor2_1
Xhold199 hold199/A vssd1 vssd1 vccd1 vccd1 hold199/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11145__A1 _12760_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08010__A1 _07347_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08010__B2 _09216_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09845_ _09843_/X _09844_/X _10176_/A vssd1 vssd1 vccd1 vccd1 _09845_/X sky130_fd_sc_hd__mux2_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09776_ _09776_/A _09776_/B vssd1 vssd1 vccd1 vccd1 _09785_/A sky130_fd_sc_hd__xor2_4
X_06988_ _06747_/Y _07110_/B _06785_/Y _13010_/B _06936_/A vssd1 vssd1 vccd1 vccd1
+ _06988_/X sky130_fd_sc_hd__o2111a_1
X_08727_ _08727_/A _08727_/B vssd1 vssd1 vccd1 vccd1 _08786_/A sky130_fd_sc_hd__xor2_4
XANTENNA__12645__A1 _12695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09510__A1 _09507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09889__A _11731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _08658_/A _08658_/B vssd1 vssd1 vccd1 vccd1 _08659_/B sky130_fd_sc_hd__and2_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_8_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13693_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ _11922_/A _10536_/A1 _10536_/B2 _11997_/A vssd1 vssd1 vccd1 vccd1 _07610_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08589_ _07238_/X _13168_/A1 _07477_/X _07239_/Y vssd1 vssd1 vccd1 vccd1 _08590_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08077__A1 _10522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10620_ _10620_/A _10620_/B vssd1 vssd1 vccd1 vccd1 _10620_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__08077__B2 _09885_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10551_ _10686_/B _10550_/C _10550_/A vssd1 vssd1 vccd1 vccd1 _10552_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__11620__A2 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10482_ _12825_/S _10478_/X _10479_/X _10481_/Y vssd1 vssd1 vccd1 vccd1 dest_val[6]
+ sky130_fd_sc_hd__a22o_4
X_13270_ hold294/A hold35/X vssd1 vssd1 vccd1 vccd1 _13473_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__11908__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12221_ reg1_val[22] curr_PC[22] vssd1 vssd1 vccd1 vccd1 _12222_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_122_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12152_ _06876_/B _09520_/X _11688_/B reg1_val[21] vssd1 vssd1 vccd1 vccd1 _12152_/Y
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__07575__C _10078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09329__A1 _07366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11103_ _11104_/A _11104_/B _11104_/C vssd1 vssd1 vccd1 vccd1 _11103_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09329__B2 _07557_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12083_ _12173_/A _12083_/B vssd1 vssd1 vccd1 vccd1 _12085_/B sky130_fd_sc_hd__and2_1
X_11034_ _12253_/A _11034_/B vssd1 vssd1 vccd1 vccd1 _11038_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08001__A1 _09173_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08001__B2 _11047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11394__A _12093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07760__B1 _08950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12985_ _12985_/A _12985_/B vssd1 vssd1 vccd1 vccd1 _12986_/B sky130_fd_sc_hd__nand2_2
XANTENNA__08304__A2 _11047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10647__B1 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11936_ _12029_/A _11936_/B vssd1 vssd1 vccd1 vccd1 _11938_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11867_ _11958_/A _11867_/B _11867_/C vssd1 vssd1 vccd1 vccd1 _11867_/X sky130_fd_sc_hd__and3_1
XFILLER_0_7_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12656__C _12754_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13606_ hold159/X _13140_/C _13568_/A vssd1 vssd1 vccd1 vccd1 hold160/A sky130_fd_sc_hd__o21a_1
X_10818_ _12087_/A fanout20/X fanout18/X _12103_/A vssd1 vssd1 vccd1 vccd1 _10819_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09265__B1 _13135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08208__A _10236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11798_ _12163_/A _12163_/B vssd1 vssd1 vccd1 vccd1 _11896_/C sky130_fd_sc_hd__or2_1
XANTENNA__07112__A _13748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13537_ hold259/X _13536_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13537_/X sky130_fd_sc_hd__mux2_1
X_10749_ _06973_/B _12793_/A2 _11586_/B vssd1 vssd1 vccd1 vccd1 _10749_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13468_ _13547_/A hold284/X vssd1 vssd1 vccd1 vccd1 _13709_/D sky130_fd_sc_hd__and2_1
XFILLER_0_23_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13364__A2 _13542_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12419_ _12668_/A _12419_/B vssd1 vssd1 vccd1 vccd1 _12421_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13399_ _07305_/B _13419_/A2 hold89/X vssd1 vssd1 vccd1 vccd1 _13681_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_23_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07960_ _07962_/A _07962_/B vssd1 vssd1 vccd1 vccd1 _07960_/X sky130_fd_sc_hd__and2_1
X_06911_ reg1_val[16] _06911_/B vssd1 vssd1 vccd1 vccd1 _06912_/B sky130_fd_sc_hd__and2_1
X_07891_ _07892_/A _07892_/B vssd1 vssd1 vccd1 vccd1 _07891_/X sky130_fd_sc_hd__and2_4
X_09630_ _09630_/A _09630_/B vssd1 vssd1 vccd1 vccd1 _09631_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06842_ _06928_/B _13025_/B vssd1 vssd1 vccd1 vccd1 _06842_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_4_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09561_ _09562_/A _09562_/B vssd1 vssd1 vccd1 vccd1 _09811_/B sky130_fd_sc_hd__and2b_1
X_06773_ instruction[0] pred_val instruction[2] vssd1 vssd1 vccd1 vccd1 _07123_/A
+ sky130_fd_sc_hd__and3b_1
X_08512_ _08512_/A _08512_/B vssd1 vssd1 vccd1 vccd1 _08565_/B sky130_fd_sc_hd__nand2_2
XANTENNA__10638__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09492_ reg1_val[6] reg1_val[25] _09493_/S vssd1 vssd1 vccd1 vccd1 _09492_/X sky130_fd_sc_hd__mux2_1
X_08443_ _09591_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08448_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout151_A _07406_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10648__A _11076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout249_A _06744_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08374_ _09501_/A _07300_/Y _11638_/A _08271_/A vssd1 vssd1 vccd1 vccd1 _08375_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08059__A1 _08821_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08059__B2 _08821_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08118__A _09381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07022__A _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07325_ _11126_/A reg1_val[14] _07328_/B _07328_/C vssd1 vssd1 vccd1 vccd1 _07513_/A
+ sky130_fd_sc_hd__or4_2
XANTENNA__11602__A2 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07256_ _07594_/B _09254_/D _07255_/X _07251_/Y vssd1 vssd1 vccd1 vccd1 _07256_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_0_104_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07187_ _07188_/C _07187_/B _07523_/A _07476_/A vssd1 vssd1 vccd1 vccd1 _07192_/B
+ sky130_fd_sc_hd__and4b_2
XFILLER_0_60_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12315__B1 _09521_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07692__A _09950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09731__A1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09731__B2 _07833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09828_ _09828_/A _09828_/B _10150_/A _10298_/A vssd1 vssd1 vccd1 vccd1 _09828_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__12103__A _12103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout64_A _11731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09759_ _11076_/A _09759_/B vssd1 vssd1 vccd1 vccd1 _09763_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12618__B2 _11823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12770_ _12773_/A _12773_/B vssd1 vssd1 vccd1 vccd1 _12770_/X sky130_fd_sc_hd__and2_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _12253_/A _11721_/B vssd1 vssd1 vccd1 vccd1 _11722_/B sky130_fd_sc_hd__xnor2_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12476__C _12476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _11652_/A _11652_/B vssd1 vssd1 vccd1 vccd1 _11654_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout50 _07223_/Y vssd1 vssd1 vccd1 vccd1 fanout50/X sky130_fd_sc_hd__clkbuf_4
Xfanout61 _10518_/A vssd1 vssd1 vccd1 vccd1 _12764_/B sky130_fd_sc_hd__clkbuf_8
Xfanout72 _07546_/X vssd1 vssd1 vccd1 vccd1 _08704_/B sky130_fd_sc_hd__buf_8
X_10603_ _10599_/X _10602_/X _10603_/S vssd1 vssd1 vccd1 vccd1 _10603_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11054__B1 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout83 fanout84/X vssd1 vssd1 vccd1 vccd1 fanout83/X sky130_fd_sc_hd__buf_6
X_11583_ _11693_/A2 _11691_/B hold195/A vssd1 vssd1 vccd1 vccd1 _11583_/Y sky130_fd_sc_hd__a21oi_1
Xfanout94 _10050_/A vssd1 vssd1 vccd1 vccd1 _11719_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13322_ _13642_/Q _13463_/B2 _13450_/B hold243/X vssd1 vssd1 vccd1 vccd1 hold244/A
+ sky130_fd_sc_hd__a22o_1
X_10534_ _10679_/B _10534_/B vssd1 vssd1 vccd1 vccd1 _10550_/A sky130_fd_sc_hd__and2_1
XFILLER_0_107_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13346__A2 _13506_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13253_ hold66/X hold289/X vssd1 vssd1 vccd1 vccd1 _13253_/X sky130_fd_sc_hd__and2b_1
X_10465_ hold287/A _12314_/A _10610_/B _12796_/A1 vssd1 vssd1 vccd1 vccd1 _10465_/X
+ sky130_fd_sc_hd__a31o_2
X_12204_ _12365_/A _12365_/B vssd1 vssd1 vccd1 vccd1 _12440_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10396_ _10397_/A _10397_/B vssd1 vssd1 vccd1 vccd1 _10398_/A sky130_fd_sc_hd__and2_1
X_13184_ _11922_/A _13194_/A2 hold117/X _13539_/A vssd1 vssd1 vccd1 vccd1 _13628_/D
+ sky130_fd_sc_hd__o211a_1
X_12135_ _12133_/X _12134_/X _12578_/A vssd1 vssd1 vccd1 vccd1 _12136_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07981__B1 wire101/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12066_ _09523_/Y _12055_/Y _12056_/X _12060_/Y _12065_/X vssd1 vssd1 vccd1 vccd1
+ _12066_/X sky130_fd_sc_hd__a311o_1
XANTENNA__09722__A1 _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ _10992_/Y _10993_/X _11003_/X _11016_/X vssd1 vssd1 vccd1 vccd1 _11017_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__12321__A3 _12235_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12609__A1 _09145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12609__B2 _12667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12968_ _12968_/A _12968_/B vssd1 vssd1 vccd1 vccd1 _12970_/A sky130_fd_sc_hd__nor2_2
XANTENNA__12667__B _12764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11919_ _11920_/A _11920_/B vssd1 vssd1 vccd1 vccd1 _11921_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12899_ _12900_/A _12900_/B _12900_/C vssd1 vssd1 vccd1 vccd1 _12907_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_74_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11045__B1 _07877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07110_ _07110_/A _07110_/B vssd1 vssd1 vccd1 vccd1 _07123_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11596__B2 _10889_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09468__S _09493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08090_ _08090_/A _08090_/B vssd1 vssd1 vccd1 vccd1 _08111_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_27_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10915__B _11825_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07041_ _06955_/Y _07040_/X _11122_/A vssd1 vssd1 vccd1 vccd1 _07041_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08992_ _08167_/A _08235_/A _08167_/C vssd1 vssd1 vccd1 vccd1 _08994_/B sky130_fd_sc_hd__a21o_1
X_07943_ _07943_/A _07943_/B vssd1 vssd1 vccd1 vccd1 _07944_/B sky130_fd_sc_hd__xnor2_4
X_07874_ _07874_/A _07874_/B vssd1 vssd1 vccd1 vccd1 _07884_/A sky130_fd_sc_hd__nand2_1
X_09613_ _09613_/A _09812_/A _09613_/C vssd1 vssd1 vccd1 vccd1 _09812_/B sky130_fd_sc_hd__nor3_1
X_06825_ instruction[35] _12981_/C vssd1 vssd1 vccd1 vccd1 _13029_/B sky130_fd_sc_hd__and2_4
X_09544_ _09881_/A _10726_/A vssd1 vssd1 vccd1 vccd1 _09656_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06756_ reg1_val[22] vssd1 vssd1 vccd1 vccd1 _07357_/A sky130_fd_sc_hd__inv_2
XANTENNA__09232__A _10078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11284__B1 _11708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09475_ reg1_val[13] reg1_val[18] _09493_/S vssd1 vssd1 vccd1 vccd1 _09475_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_65_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08426_ _08485_/A _08485_/B vssd1 vssd1 vccd1 vccd1 _08503_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_93_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08357_ _08357_/A _08357_/B vssd1 vssd1 vccd1 vccd1 _08411_/A sky130_fd_sc_hd__or2_1
XFILLER_0_18_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07308_ _07312_/B _10649_/A _10537_/A vssd1 vssd1 vccd1 vccd1 _07308_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_6_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07255__A2 _07213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08288_ _08288_/A _08288_/B _08288_/C vssd1 vssd1 vccd1 vccd1 _08293_/A sky130_fd_sc_hd__and3_1
XFILLER_0_6_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13328__A2 _13506_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07239_ _07240_/A _07240_/B vssd1 vssd1 vccd1 vccd1 _07239_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__13201__B _13207_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12536__B1 _09519_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10250_ _10250_/A _10250_/B vssd1 vssd1 vccd1 vccd1 _10252_/B sky130_fd_sc_hd__xnor2_2
X_10181_ _10170_/Y _10180_/Y _12648_/A vssd1 vssd1 vccd1 vccd1 _10181_/X sky130_fd_sc_hd__mux2_1
Xfanout240 _12327_/A vssd1 vssd1 vccd1 vccd1 _12971_/S sky130_fd_sc_hd__buf_8
Xfanout251 _13141_/A vssd1 vssd1 vccd1 vccd1 _13463_/B2 sky130_fd_sc_hd__buf_4
Xfanout262 _12979_/A vssd1 vssd1 vccd1 vccd1 _12956_/A sky130_fd_sc_hd__buf_8
Xfanout273 _13444_/C1 vssd1 vssd1 vccd1 vccd1 _13459_/A sky130_fd_sc_hd__clkbuf_4
Xfanout284 _06762_/Y vssd1 vssd1 vccd1 vccd1 _12738_/S sky130_fd_sc_hd__buf_2
XANTENNA__11511__A1 _12557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout295 _12578_/A vssd1 vssd1 vccd1 vccd1 _10734_/A sky130_fd_sc_hd__buf_4
XANTENNA__09841__S _10004_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11511__B2 _12557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12822_ _12823_/A _12823_/B _12823_/C vssd1 vssd1 vccd1 vccd1 _12830_/B sky130_fd_sc_hd__a21o_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12753_ _12753_/A _12753_/B vssd1 vssd1 vccd1 vccd1 _12753_/Y sky130_fd_sc_hd__nor2_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ fanout29/X _09146_/Y fanout5/A fanout27/X vssd1 vssd1 vccd1 vccd1 _11705_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _12571_/X _12682_/D _12683_/X vssd1 vssd1 vccd1 vccd1 _12684_/X sky130_fd_sc_hd__a21o_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11635_ wire101/X fanout9/A fanout4/X _13180_/A1 vssd1 vssd1 vccd1 vccd1 _11636_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13567__A2 _13584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07597__A _10787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11566_ _11958_/A _11566_/B vssd1 vssd1 vccd1 vccd1 _11566_/Y sky130_fd_sc_hd__nor2_1
X_13305_ _13233_/B _13548_/B _13233_/A vssd1 vssd1 vccd1 vccd1 _13553_/A sky130_fd_sc_hd__o21bai_1
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10517_ wire122/X fanout9/X fanout4/X _10637_/A vssd1 vssd1 vccd1 vccd1 _10518_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11497_ _11498_/A _11498_/B vssd1 vssd1 vccd1 vccd1 _11646_/A sky130_fd_sc_hd__and2_1
XANTENNA__12008__A _12092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13236_ _13236_/A _13236_/B vssd1 vssd1 vccd1 vccd1 _13544_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10448_ _12515_/S _10589_/B _10447_/X vssd1 vssd1 vccd1 vccd1 _10449_/B sky130_fd_sc_hd__a21o_1
X_13167_ hold62/X _13191_/B vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__or2_1
XFILLER_0_0_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10379_ _10379_/A _10379_/B vssd1 vssd1 vccd1 vccd1 _10380_/B sky130_fd_sc_hd__xor2_2
X_12118_ _12120_/A _12120_/B _12120_/C vssd1 vssd1 vccd1 vccd1 _12121_/A sky130_fd_sc_hd__a21o_1
X_13098_ _13098_/A _13102_/D vssd1 vssd1 vccd1 vccd1 loadstore_address[23] sky130_fd_sc_hd__xnor2_4
XFILLER_0_46_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12049_ reg1_val[20] curr_PC[20] vssd1 vssd1 vccd1 vccd1 _12050_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10305__A2 _10727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09171__A2 _11047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07590_ _09951_/A _07590_/B vssd1 vssd1 vccd1 vccd1 _07603_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09459__A0 _11126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08131__A0 _10119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12463__C1 _09529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09260_ _09260_/A _09260_/B vssd1 vssd1 vccd1 vccd1 _09261_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__08682__A1 _08873_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08891__A _09674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08682__B2 _08891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08211_ _08214_/A _08214_/B vssd1 vssd1 vccd1 vccd1 _08290_/A sky130_fd_sc_hd__nand2_1
X_09191_ _09190_/A _09190_/B _09192_/A vssd1 vssd1 vccd1 vccd1 _09191_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_62_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07890__C1 _09254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08142_ _08140_/A _08140_/B _08177_/A vssd1 vssd1 vccd1 vccd1 _08150_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__08434__A1 _08873_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08434__B2 _08891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08073_ _11708_/A _08073_/B vssd1 vssd1 vccd1 vccd1 _08080_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07024_ _09694_/A _10004_/S vssd1 vssd1 vccd1 vccd1 _07024_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08198__B1 _08907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08737__A2 _08866_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08975_ _08844_/A _08842_/X _08976_/A vssd1 vssd1 vccd1 vccd1 _08975_/Y sky130_fd_sc_hd__a21oi_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__buf_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ _07927_/A _07927_/B vssd1 vssd1 vccd1 vccd1 _07926_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12297__A2 _12372_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09162__A2 _07643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07857_ _10049_/A2 _08246_/B _09885_/B1 fanout21/X vssd1 vssd1 vccd1 vccd1 _07858_/B
+ sky130_fd_sc_hd__o22a_1
X_06808_ instruction[39] _12981_/C vssd1 vssd1 vccd1 vccd1 _13054_/B sky130_fd_sc_hd__and2_4
X_07788_ _07788_/A _07788_/B vssd1 vssd1 vccd1 vccd1 _07798_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_78_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09527_ _07091_/B _11586_/B _09523_/Y hold188/A _09526_/X vssd1 vssd1 vccd1 vccd1
+ _09527_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09458_ _09454_/X _09457_/X _10005_/S vssd1 vssd1 vccd1 vccd1 _09458_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout27_A _07453_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08409_ _08416_/A _08416_/B _08399_/X vssd1 vssd1 vccd1 vccd1 _08466_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_47_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09389_ _09389_/A _09389_/B vssd1 vssd1 vccd1 vccd1 _09390_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12754__C _12754_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11420_ _11802_/B _11420_/B vssd1 vssd1 vccd1 vccd1 _11426_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07228__A2 _07213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09622__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11351_ _11864_/A _09032_/X _09034_/C _10866_/B vssd1 vssd1 vccd1 vccd1 _11352_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10302_ _10302_/A _10302_/B vssd1 vssd1 vccd1 vccd1 _10303_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11282_ _11282_/A _12614_/A vssd1 vssd1 vccd1 vccd1 _11285_/B sky130_fd_sc_hd__nand2_1
X_13021_ _13019_/Y _13021_/B vssd1 vssd1 vccd1 vccd1 _13022_/B sky130_fd_sc_hd__nand2b_2
X_10233_ _10233_/A _10233_/B vssd1 vssd1 vccd1 vccd1 _10234_/B sky130_fd_sc_hd__or2_1
XANTENNA__09137__A _09591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10164_ _10165_/A _10165_/B vssd1 vssd1 vccd1 vccd1 _10164_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_100_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10095_ _10095_/A _10095_/B vssd1 vssd1 vccd1 vccd1 _10099_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07880__A _11731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12805_ _12806_/A _12806_/B vssd1 vssd1 vccd1 vccd1 _12816_/A sky130_fd_sc_hd__nand2_1
X_10997_ _10876_/A _10873_/Y _10875_/B vssd1 vssd1 vccd1 vccd1 _10999_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12736_ _12736_/A _12736_/B vssd1 vssd1 vccd1 vccd1 _12736_/Y sky130_fd_sc_hd__nor2_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12667_ _12667_/A _12764_/B vssd1 vssd1 vccd1 vccd1 _12668_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12748__B1 _12748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11618_ _11712_/A _11618_/B vssd1 vssd1 vccd1 vccd1 _11619_/B sky130_fd_sc_hd__nor2_1
X_12598_ _12598_/A _12598_/B _12598_/C vssd1 vssd1 vccd1 vccd1 _12598_/X sky130_fd_sc_hd__or3_1
XFILLER_0_108_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11549_ _11549_/A _11549_/B vssd1 vssd1 vccd1 vccd1 _11551_/C sky130_fd_sc_hd__xor2_2
XFILLER_0_123_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13219_ hold273/A hold42/X vssd1 vssd1 vccd1 vccd1 _13569_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__10481__A _12825_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10526__A2 _11423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_10_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13684_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10631__D _10981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08760_ _08786_/A _08786_/B vssd1 vssd1 vccd1 vccd1 _08760_/Y sky130_fd_sc_hd__nand2_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07790__A _09591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07711_ _07964_/A _07964_/B vssd1 vssd1 vccd1 vccd1 _07965_/A sky130_fd_sc_hd__or2_1
X_08691_ _08699_/A _08699_/B _08679_/X vssd1 vssd1 vccd1 vccd1 _08722_/A sky130_fd_sc_hd__a21o_2
X_07642_ _07642_/A _07876_/A vssd1 vssd1 vccd1 vccd1 _07642_/X sky130_fd_sc_hd__and2_1
X_07573_ _10537_/A _07575_/B vssd1 vssd1 vccd1 vccd1 _10934_/A sky130_fd_sc_hd__nor2_1
X_09312_ _09313_/A _09313_/B vssd1 vssd1 vccd1 vccd1 _09828_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_87_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09243_ _09940_/A _09243_/B vssd1 vssd1 vccd1 vccd1 _09246_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout231_A _11688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09174_ _10266_/A _09174_/B vssd1 vssd1 vccd1 vccd1 _09176_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07030__A _09501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08125_ _08125_/A _08125_/B _08125_/C vssd1 vssd1 vccd1 vccd1 _08130_/A sky130_fd_sc_hd__or3_1
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08056_ _09381_/A fanout39/X _08118_/B _08873_/B2 vssd1 vssd1 vccd1 vccd1 _08057_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_113_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07007_ reg1_val[3] _10457_/S vssd1 vssd1 vccd1 vccd1 _07007_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_12_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10517__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07918__B1 _07557_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09383__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08958_ _09004_/A _09004_/B vssd1 vssd1 vccd1 vccd1 _09005_/A sky130_fd_sc_hd__nor2_1
XANTENNA__13467__B2 _13542_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07909_ _07909_/A _07909_/B vssd1 vssd1 vccd1 vccd1 _07911_/B sky130_fd_sc_hd__xnor2_2
X_08889_ _08889_/A _08889_/B _08889_/C vssd1 vssd1 vccd1 vccd1 _08897_/A sky130_fd_sc_hd__and3_1
XFILLER_0_98_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10920_ _07282_/X fanout38/X fanout36/X _12087_/A vssd1 vssd1 vccd1 vccd1 _10921_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07697__A2 _08118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06873__A2_N _06906_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10851_ _10852_/A _10852_/B _10852_/C vssd1 vssd1 vccd1 vccd1 _10851_/X sky130_fd_sc_hd__a21o_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13570_ _13570_/A _13570_/B vssd1 vssd1 vccd1 vccd1 _13570_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10782_ _10783_/A _10783_/B _10781_/X vssd1 vssd1 vccd1 vccd1 _10962_/B sky130_fd_sc_hd__o21ba_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ reg1_val[26] curr_PC[26] vssd1 vssd1 vccd1 vccd1 _12521_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_109_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06888__A2_N _06906_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12452_ _12452_/A _12452_/B vssd1 vssd1 vccd1 vccd1 _12452_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_35_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10205__A1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11403_ _12092_/A _11403_/B vssd1 vssd1 vccd1 vccd1 _11521_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10205__B2 _07833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11402__B1 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12781__A _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12383_ _12382_/A _12382_/B _12382_/Y _09506_/X vssd1 vssd1 vccd1 vccd1 _12383_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11953__A1 _12695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11334_ _11334_/A _11334_/B vssd1 vssd1 vccd1 vccd1 _11337_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07621__A2 _09955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07594__B _07594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11265_ curr_PC[11] curr_PC[12] _11265_/C vssd1 vssd1 vccd1 vccd1 _11266_/B sky130_fd_sc_hd__and3_1
XFILLER_0_30_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13004_ reg1_val[5] _13005_/B vssd1 vssd1 vccd1 vccd1 _13004_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09374__A2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10216_ _10217_/A _10217_/B _10217_/C vssd1 vssd1 vccd1 vccd1 _10218_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11196_ _11058_/X _11062_/A _07477_/X _11802_/B vssd1 vssd1 vccd1 vccd1 _11326_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10147_ _10148_/A _10148_/B vssd1 vssd1 vccd1 vccd1 _10147_/X sky130_fd_sc_hd__and2_1
XANTENNA__13458__B2 _13463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09126__A2 _10235_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10078_ _10078_/A _10078_/B vssd1 vssd1 vccd1 vccd1 _10080_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09834__B1 _11866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09330__A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12719_ fanout10/X _12718_/Y _12717_/Y _12764_/B vssd1 vssd1 vccd1 vccd1 _12769_/S
+ sky130_fd_sc_hd__o2bb2a_1
X_13699_ _13700_/CLK _13699_/D vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09930_ _09931_/B _09931_/C _10542_/A vssd1 vssd1 vccd1 vccd1 _09932_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_21_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09861_ _13642_/Q hold188/A _10606_/A2 vssd1 vssd1 vccd1 vccd1 _09862_/B sky130_fd_sc_hd__o21ai_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08812_ _08846_/A _08816_/B _08805_/Y vssd1 vssd1 vccd1 vccd1 _08815_/B sky130_fd_sc_hd__a21bo_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _12094_/A _09792_/B vssd1 vssd1 vccd1 vccd1 _09800_/A sky130_fd_sc_hd__xnor2_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ _08755_/A _08755_/B _08756_/B vssd1 vssd1 vccd1 vccd1 _08743_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09505__A _10734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12657__C1 _12799_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout279_A _13444_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08674_ _08677_/A _08677_/B vssd1 vssd1 vccd1 vccd1 _08674_/X sky130_fd_sc_hd__and2_1
XFILLER_0_68_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07625_ fanout39/X _07366_/X _08118_/B _07557_/Y vssd1 vssd1 vccd1 vccd1 _07626_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06887__B1 _06906_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07556_ _07556_/A _07557_/B vssd1 vssd1 vccd1 vccd1 _07556_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_119_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10386__A _11709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07487_ _12094_/A _07493_/B vssd1 vssd1 vccd1 vccd1 _07487_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_119_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09226_ _09135_/A _09135_/B _09138_/Y vssd1 vssd1 vccd1 vccd1 _09230_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_91_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07398__C _09703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09157_ _12754_/A _12754_/B _07637_/B vssd1 vssd1 vccd1 vccd1 _09157_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_16_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08108_ _08108_/A _08108_/B vssd1 vssd1 vccd1 vccd1 _08164_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08800__A1 _08950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09088_ _09087_/A _09087_/B _09082_/A _09082_/B _09082_/C vssd1 vssd1 vccd1 vccd1
+ _12583_/B sky130_fd_sc_hd__a2111o_1
XANTENNA__08800__B2 _08866_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08039_ _08039_/A _08039_/B vssd1 vssd1 vccd1 vccd1 _08098_/A sky130_fd_sc_hd__xor2_1
XANTENNA_fanout94_A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11050_ _11050_/A _11050_/B vssd1 vssd1 vccd1 vccd1 _11051_/B sky130_fd_sc_hd__and2_1
X_10001_ _09671_/X _09673_/X _10005_/S vssd1 vssd1 vccd1 vccd1 _10001_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_99_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11952_ _12035_/B _11952_/B vssd1 vssd1 vccd1 vccd1 _12164_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__12663__A2 _10889_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10903_ _12551_/A _10903_/B vssd1 vssd1 vccd1 vccd1 _10910_/A sky130_fd_sc_hd__xnor2_1
X_11883_ hold259/A _12058_/A _11969_/B _11882_/Y _12748_/B1 vssd1 vssd1 vccd1 vccd1
+ _11889_/D sky130_fd_sc_hd__a311o_1
X_13622_ _13717_/CLK _13622_/D vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__dfxtp_1
X_10834_ _10834_/A _10834_/B vssd1 vssd1 vccd1 vccd1 _10847_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_66_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13553_ _13553_/A _13553_/B vssd1 vssd1 vccd1 vccd1 _13553_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__11623__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10765_ _12825_/S _10761_/X _10762_/X _10764_/Y vssd1 vssd1 vccd1 vccd1 dest_val[8]
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_81_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12504_ _12505_/A _12505_/B _12505_/C vssd1 vssd1 vccd1 vccd1 _12506_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13484_ _13484_/A _13484_/B vssd1 vssd1 vccd1 vccd1 _13484_/Y sky130_fd_sc_hd__xnor2_1
X_10696_ _10696_/A _10696_/B vssd1 vssd1 vccd1 vccd1 _10697_/B sky130_fd_sc_hd__or2_1
XFILLER_0_23_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13376__B1 _13584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12435_ _12435_/A _12435_/B vssd1 vssd1 vccd1 vccd1 _12437_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09595__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12366_ _12208_/A _12368_/C _12364_/X vssd1 vssd1 vccd1 vccd1 _12629_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11317_ _11318_/B _11318_/A vssd1 vssd1 vccd1 vccd1 _11438_/B sky130_fd_sc_hd__nand2b_1
X_12297_ _12296_/A _12372_/D _11955_/A vssd1 vssd1 vccd1 vccd1 _12297_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_38_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11248_ hold209/A _13651_/Q _11248_/C vssd1 vssd1 vccd1 vccd1 _11366_/B sky130_fd_sc_hd__or3_1
XANTENNA__11154__A2 _11802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11179_ fanout47/X fanout20/X fanout18/X fanout46/X vssd1 vssd1 vccd1 vccd1 _11180_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06949__A _11126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07410_ _07410_/A _07535_/B vssd1 vssd1 vccd1 vccd1 _07414_/D sky130_fd_sc_hd__nand2_1
X_08390_ _08454_/A _08454_/B vssd1 vssd1 vccd1 vccd1 _08455_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_70_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07341_ _07336_/Y _07340_/X _07637_/B vssd1 vssd1 vccd1 vccd1 _07414_/B sky130_fd_sc_hd__a21o_2
XANTENNA__11614__B1 _11708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09283__A1 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09283__B2 _08395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07272_ _07535_/B _07270_/X _07271_/X vssd1 vssd1 vccd1 vccd1 _07274_/B sky130_fd_sc_hd__o21ai_2
X_09011_ _10160_/B _10160_/C vssd1 vssd1 vccd1 vccd1 _10306_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_116_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11917__A1 _07198_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11917__B2 _11997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold101 hold101/A vssd1 vssd1 vccd1 vccd1 hold101/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 hold112/A vssd1 vssd1 vccd1 vccd1 hold112/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 hold123/A vssd1 vssd1 vccd1 vccd1 hold123/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11393__A2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08794__B1 _09216_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold134 hold134/A vssd1 vssd1 vccd1 vccd1 hold134/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 hold145/A vssd1 vssd1 vccd1 vccd1 hold145/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 hold156/A vssd1 vssd1 vccd1 vccd1 hold156/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold167 hold167/A vssd1 vssd1 vccd1 vccd1 hold167/X sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ _09914_/B _09914_/A vssd1 vssd1 vccd1 vccd1 _10134_/B sky130_fd_sc_hd__nand2b_1
Xhold178 hold178/A vssd1 vssd1 vccd1 vccd1 hold178/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 hold189/A vssd1 vssd1 vccd1 vccd1 hold189/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09844_ _09457_/X _09461_/X _10005_/S vssd1 vssd1 vccd1 vccd1 _09844_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_95_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08010__A2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ _09773_/X _09775_/B vssd1 vssd1 vccd1 vccd1 _09776_/B sky130_fd_sc_hd__nand2b_2
X_06987_ _10590_/A _10589_/A vssd1 vssd1 vccd1 vccd1 _10449_/A sky130_fd_sc_hd__nor2_1
X_08726_ _08726_/A _08726_/B vssd1 vssd1 vccd1 vccd1 _09044_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_68_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08657_ _08980_/A _08980_/B _08983_/A vssd1 vssd1 vccd1 vccd1 _08657_/X sky130_fd_sc_hd__a21o_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07608_ _07671_/A _07671_/B vssd1 vssd1 vccd1 vccd1 _07672_/A sky130_fd_sc_hd__nand2_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08588_ _08588_/A _08588_/B vssd1 vssd1 vccd1 vccd1 _08643_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07539_ _07537_/B _07537_/C _11076_/A vssd1 vssd1 vccd1 vccd1 _11157_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__08077__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10550_ _10550_/A _10686_/B _10550_/C vssd1 vssd1 vccd1 vccd1 _10552_/B sky130_fd_sc_hd__and3_1
XFILLER_0_106_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09209_ _09198_/A _09198_/B _09199_/X vssd1 vssd1 vccd1 vccd1 _09313_/A sky130_fd_sc_hd__a21o_2
XANTENNA__13358__B1 _13506_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10481_ _12825_/S _10763_/C vssd1 vssd1 vccd1 vccd1 _10481_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11908__A1 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12220_ reg1_val[22] curr_PC[22] vssd1 vssd1 vccd1 vccd1 _12222_/A sky130_fd_sc_hd__or2_1
XANTENNA__11908__B2 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12151_ _12151_/A _12151_/B vssd1 vssd1 vccd1 vccd1 _12151_/X sky130_fd_sc_hd__or2_1
X_11102_ _11104_/A _11104_/B _11104_/C vssd1 vssd1 vccd1 vccd1 _11105_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__09329__A2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12082_ _12082_/A _12082_/B vssd1 vssd1 vccd1 vccd1 _12083_/B sky130_fd_sc_hd__or2_1
XANTENNA__08537__B1 _08778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11033_ _12087_/A fanout38/X fanout36/X _12103_/A vssd1 vssd1 vccd1 vccd1 _11034_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08001__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09145__A _09254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07760__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07760__B2 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12984_ _12985_/A _12985_/B vssd1 vssd1 vccd1 vccd1 _12984_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10647__A1 _10538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11935_ _11935_/A _11935_/B _11935_/C vssd1 vssd1 vccd1 vccd1 _11936_/B sky130_fd_sc_hd__and3_1
XFILLER_0_86_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11866_ _11866_/A _11866_/B vssd1 vssd1 vccd1 vccd1 _11866_/Y sky130_fd_sc_hd__nand2_1
X_13605_ _13605_/A _13605_/B hold144/X vssd1 vssd1 vccd1 vccd1 hold145/A sky130_fd_sc_hd__and3_1
X_10817_ _12421_/A _10817_/B vssd1 vssd1 vccd1 vccd1 _10821_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11797_ _12406_/B1 _11792_/X _11793_/Y _11796_/Y vssd1 vssd1 vccd1 vccd1 dest_val[17]
+ sky130_fd_sc_hd__o31a_4
XFILLER_0_6_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07112__B _13744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13536_ _13536_/A _13536_/B vssd1 vssd1 vccd1 vccd1 _13536_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10748_ _10748_/A _12056_/B hold163/A vssd1 vssd1 vccd1 vccd1 _10748_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_125_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13467_ hold283/X _13555_/A2 _13466_/X _13542_/B2 vssd1 vssd1 vccd1 vccd1 hold284/A
+ sky130_fd_sc_hd__a22o_1
X_10679_ _10679_/A _10679_/B _10679_/C vssd1 vssd1 vccd1 vccd1 _10680_/B sky130_fd_sc_hd__and3_1
XFILLER_0_125_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12418_ _12614_/A fanout12/X _12667_/A fanout16/X vssd1 vssd1 vccd1 vccd1 _12419_/B
+ sky130_fd_sc_hd__a22o_1
X_13398_ hold5/X _13416_/A2 _13420_/B1 hold64/X _13383_/A vssd1 vssd1 vccd1 vccd1
+ hold89/A sky130_fd_sc_hd__o221a_1
XFILLER_0_49_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12349_ _12426_/B _12349_/B vssd1 vssd1 vccd1 vccd1 _12351_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_11_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12324__B2 _10866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06910_ _06910_/A vssd1 vssd1 vccd1 vccd1 _06912_/A sky130_fd_sc_hd__inv_2
X_07890_ _07521_/A _07595_/A _07595_/B _09254_/B vssd1 vssd1 vccd1 vccd1 _07892_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_65_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06841_ instruction[34] _12981_/C vssd1 vssd1 vccd1 vccd1 _13025_/B sky130_fd_sc_hd__and2_4
XFILLER_0_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09560_ _09811_/A _09560_/B vssd1 vssd1 vccd1 vccd1 _09562_/B sky130_fd_sc_hd__nor2_2
X_06772_ instruction[22] instruction[15] _07135_/S vssd1 vssd1 vccd1 vccd1 reg1_idx[4]
+ sky130_fd_sc_hd__mux2_8
X_08511_ _08518_/A _08518_/B vssd1 vssd1 vccd1 vccd1 _08512_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__10638__A1 _07477_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09491_ _09489_/X _09490_/X _09688_/S vssd1 vssd1 vccd1 vccd1 _09491_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10638__B2 _07472_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08442_ _13149_/A fanout84/X _08580_/B _08923_/B1 vssd1 vssd1 vccd1 vccd1 _08443_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_58_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13588__B1 _13568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08373_ _08951_/A _08373_/B vssd1 vssd1 vccd1 vccd1 _08418_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13024__B _13025_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08059__A2 _11732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08118__B _08118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07267__A0 _13015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07022__B _10007_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07324_ _07531_/A _07571_/A _07324_/C vssd1 vssd1 vccd1 vccd1 _11372_/A sky130_fd_sc_hd__and3_1
XFILLER_0_73_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07255_ _07217_/A _07213_/A _07213_/B _07214_/Y _07251_/A vssd1 vssd1 vccd1 vccd1
+ _07255_/X sky130_fd_sc_hd__a41o_1
XFILLER_0_116_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07186_ _07476_/A _07186_/B _07186_/C _07187_/B vssd1 vssd1 vccd1 vccd1 _07521_/B
+ sky130_fd_sc_hd__and4_2
XANTENNA__08767__B1 _09910_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09664__S _09703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10603__S _10603_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09827_ _09650_/A _09650_/B _09826_/X vssd1 vssd1 vccd1 vccd1 _09827_/X sky130_fd_sc_hd__a21o_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09731__A2 wire122/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12103__B _12666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09758_ fanout47/X fanout68/X fanout66/X fanout45/X vssd1 vssd1 vccd1 vccd1 _09759_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12079__B1 _07699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12618__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08709_ _08907_/A _09173_/B2 _11047_/A _08197_/A vssd1 vssd1 vccd1 vccd1 _08710_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_68_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11826__B1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09689_ _09687_/X _09688_/X _10005_/S vssd1 vssd1 vccd1 vccd1 _09689_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_69_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _12557_/A fanout38/X fanout36/X _12557_/B vssd1 vssd1 vccd1 vccd1 _11721_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07213__A _07213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11651_ _11652_/B _11652_/A vssd1 vssd1 vccd1 vccd1 _11651_/Y sky130_fd_sc_hd__nand2b_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout40 _12087_/A vssd1 vssd1 vccd1 vccd1 fanout40/X sky130_fd_sc_hd__buf_6
Xfanout51 _07217_/Y vssd1 vssd1 vccd1 vccd1 fanout51/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__07258__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10602_ _10457_/S _10600_/X _10601_/X vssd1 vssd1 vccd1 vccd1 _10602_/X sky130_fd_sc_hd__a21o_1
Xfanout62 _10518_/A vssd1 vssd1 vccd1 vccd1 _11802_/B sky130_fd_sc_hd__buf_4
XANTENNA__11054__A1 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11054__B2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11582_ hold193/A hold297/A _11582_/C vssd1 vssd1 vccd1 vccd1 _11691_/B sky130_fd_sc_hd__or3_1
XFILLER_0_9_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout84 _07520_/X vssd1 vssd1 vccd1 vccd1 fanout84/X sky130_fd_sc_hd__buf_8
XFILLER_0_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout95 _07381_/X vssd1 vssd1 vccd1 vccd1 _10050_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13321_ _13459_/A hold189/X vssd1 vssd1 vccd1 vccd1 hold190/A sky130_fd_sc_hd__and2_1
X_10533_ _10533_/A _10533_/B vssd1 vssd1 vccd1 vccd1 _10534_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_107_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_588 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13252_ hold251/X hold90/X vssd1 vssd1 vccd1 vccd1 _13518_/B sky130_fd_sc_hd__nand2b_1
X_10464_ _12314_/A _10610_/B hold287/A vssd1 vssd1 vccd1 vccd1 _10464_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_122_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12203_ _12203_/A _12203_/B _12203_/C vssd1 vssd1 vccd1 vccd1 _12365_/B sky130_fd_sc_hd__and3_1
XFILLER_0_60_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13183_ hold116/X _13191_/B vssd1 vssd1 vccd1 vccd1 hold117/A sky130_fd_sc_hd__or2_1
X_10395_ _10395_/A _10395_/B vssd1 vssd1 vccd1 vccd1 _10397_/B sky130_fd_sc_hd__xnor2_1
X_12134_ _12046_/A _07050_/Y _07055_/Y vssd1 vssd1 vccd1 vccd1 _12134_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_102_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07981__A1 _08933_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07981__B2 _07175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12065_ _12710_/B2 _11131_/X _11143_/X _12537_/B2 _12064_/X vssd1 vssd1 vccd1 vccd1
+ _12065_/X sky130_fd_sc_hd__a221o_1
X_11016_ _12537_/B2 _11001_/X _12143_/B _12710_/B2 _11014_/Y vssd1 vssd1 vccd1 vccd1
+ _11016_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_126_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12609__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12967_ _12979_/A _12967_/B vssd1 vssd1 vccd1 vccd1 _12968_/B sky130_fd_sc_hd__nor2_1
X_11918_ _12666_/A _11918_/B vssd1 vssd1 vccd1 vccd1 _11920_/B sky130_fd_sc_hd__xnor2_1
X_12898_ _12907_/A _12898_/B vssd1 vssd1 vccd1 vccd1 _12900_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11849_ _11849_/A _11849_/B vssd1 vssd1 vccd1 vccd1 _11851_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07249__B1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11045__B2 _11423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13519_ _13519_/A _13519_/B vssd1 vssd1 vccd1 vccd1 _13519_/Y sky130_fd_sc_hd__xnor2_1
X_07040_ _06962_/Y _07039_/Y _10992_/A vssd1 vssd1 vccd1 vccd1 _07040_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_113_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12545__A1 _07108_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09484__S _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08991_ _08990_/A _08990_/B _09003_/A vssd1 vssd1 vccd1 vccd1 _08991_/X sky130_fd_sc_hd__a21o_1
X_07942_ _07943_/B _07943_/A vssd1 vssd1 vccd1 vccd1 _09190_/B sky130_fd_sc_hd__and2b_1
X_07873_ _07873_/A _07873_/B vssd1 vssd1 vccd1 vccd1 _07945_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__13019__B _13020_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08921__B1 _09910_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09612_ _09726_/B _09611_/B _09611_/C vssd1 vssd1 vccd1 vccd1 _09613_/C sky130_fd_sc_hd__a21oi_1
X_06824_ _06824_/A _06824_/B vssd1 vssd1 vccd1 vccd1 _12642_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07017__B _09496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09543_ _10342_/A _09541_/X _09542_/X vssd1 vssd1 vccd1 vccd1 dest_val[0] sky130_fd_sc_hd__o21ai_4
XANTENNA__09513__A _13744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06755_ reg1_val[21] vssd1 vssd1 vccd1 vccd1 _07348_/A sky130_fd_sc_hd__inv_2
XANTENNA__11808__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09474_ reg1_val[12] reg1_val[19] _09493_/S vssd1 vssd1 vccd1 vccd1 _09474_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_66_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08425_ _09659_/B _08425_/B vssd1 vssd1 vccd1 vccd1 _08485_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08356_ _08368_/A _08368_/B vssd1 vssd1 vccd1 vccd1 _08357_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_46_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12233__B1 _12796_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07307_ _10537_/A _10649_/A _07306_/X vssd1 vssd1 vccd1 vccd1 _07307_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__11587__A2 _11587_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08287_ _08287_/A _08287_/B vssd1 vssd1 vccd1 vccd1 _08288_/C sky130_fd_sc_hd__nor2_1
XANTENNA__07660__B1 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07238_ _07240_/A _07240_/B _08951_/A vssd1 vssd1 vccd1 vccd1 _07238_/X sky130_fd_sc_hd__mux2_8
XFILLER_0_116_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07169_ reg1_val[4] _07168_/X _07572_/S vssd1 vssd1 vccd1 vccd1 _07172_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_14_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10180_ _10458_/S _10179_/X _10175_/X vssd1 vssd1 vccd1 vccd1 _10180_/Y sky130_fd_sc_hd__a21oi_2
Xfanout230 _09705_/X vssd1 vssd1 vccd1 vccd1 _12314_/A sky130_fd_sc_hd__clkbuf_8
Xfanout241 _07106_/Y vssd1 vssd1 vccd1 vccd1 _12327_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__07208__A _07535_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout252 _13141_/A vssd1 vssd1 vccd1 vccd1 _13542_/B2 sky130_fd_sc_hd__buf_4
Xfanout263 _13082_/A vssd1 vssd1 vccd1 vccd1 _12979_/A sky130_fd_sc_hd__buf_4
Xfanout274 _13444_/C1 vssd1 vssd1 vccd1 vccd1 _13543_/A sky130_fd_sc_hd__buf_4
Xfanout285 _06748_/Y vssd1 vssd1 vccd1 vccd1 _08197_/A sky130_fd_sc_hd__buf_6
XANTENNA__11511__A2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout296 instruction[7] vssd1 vssd1 vccd1 vccd1 _12578_/A sky130_fd_sc_hd__buf_4
X_12821_ _12830_/A _12821_/B vssd1 vssd1 vccd1 vccd1 _12823_/C sky130_fd_sc_hd__nand2_1
XANTENNA__07479__B1 _08486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12752_ hold224/A _12374_/A _12750_/X _12795_/A1 vssd1 vssd1 vccd1 vccd1 _12753_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _11601_/X _12163_/A _12695_/A vssd1 vssd1 vccd1 vccd1 _11703_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_84_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _12567_/X _12626_/A _12626_/B vssd1 vssd1 vccd1 vccd1 _12683_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_127_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _10944_/A _11508_/B _11509_/X vssd1 vssd1 vccd1 vccd1 _11637_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07597__B _10787_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11565_ _07094_/B _11463_/B _06927_/B vssd1 vssd1 vccd1 vccd1 _11566_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_64_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13304_ _13544_/A _13544_/B _13236_/A vssd1 vssd1 vccd1 vccd1 _13548_/B sky130_fd_sc_hd__a21oi_1
X_10516_ _10516_/A _10516_/B vssd1 vssd1 vccd1 vccd1 _10554_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_107_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11496_ _11719_/A _11496_/B vssd1 vssd1 vccd1 vccd1 _11498_/B sky130_fd_sc_hd__xnor2_1
X_13235_ hold275/A hold85/X vssd1 vssd1 vccd1 vccd1 _13236_/B sky130_fd_sc_hd__and2b_1
X_10447_ _10734_/A _10447_/B _10447_/C vssd1 vssd1 vccd1 vccd1 _10447_/X sky130_fd_sc_hd__and3_1
X_13166_ _13166_/A1 _13194_/A2 hold106/X _13543_/A vssd1 vssd1 vccd1 vccd1 _13619_/D
+ sky130_fd_sc_hd__o211a_1
X_10378_ _10379_/A _10379_/B vssd1 vssd1 vccd1 vccd1 _10378_/X sky130_fd_sc_hd__and2_1
X_12117_ _12117_/A _12117_/B vssd1 vssd1 vccd1 vccd1 _12120_/C sky130_fd_sc_hd__xnor2_1
X_13097_ reg1_val[23] _13129_/B vssd1 vssd1 vccd1 vccd1 _13102_/D sky130_fd_sc_hd__xnor2_4
XANTENNA__09156__B1 _13129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12048_ reg1_val[20] curr_PC[20] vssd1 vssd1 vccd1 vccd1 _12050_/A sky130_fd_sc_hd__or2_1
XANTENNA__13554__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09333__A _11731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08891__B _08891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08682__A2 _09216_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08210_ _08746_/A _08210_/B vssd1 vssd1 vccd1 vccd1 _08214_/B sky130_fd_sc_hd__xnor2_2
X_09190_ _09190_/A _09190_/B vssd1 vssd1 vccd1 vccd1 _09192_/B sky130_fd_sc_hd__nor2_2
XANTENNA__11018__B2 _11866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08141_ _08176_/A _08176_/B vssd1 vssd1 vccd1 vccd1 _08177_/A sky130_fd_sc_hd__or2_1
XFILLER_0_43_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08434__A2 _09173_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08072_ _09216_/B2 fanout24/X _08486_/B _08868_/B1 vssd1 vssd1 vccd1 vccd1 _08073_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_125_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07023_ _07025_/B _07025_/C _12985_/A vssd1 vssd1 vccd1 vccd1 _07026_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08974_ _08974_/A _08974_/B vssd1 vssd1 vccd1 vccd1 _09028_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09147__B1 _10536_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ _09179_/B _07925_/B vssd1 vssd1 vccd1 vccd1 _07927_/B sky130_fd_sc_hd__nand2_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09698__A1 _12525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12869__A _13029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07856_ _10263_/A _07856_/B vssd1 vssd1 vccd1 vccd1 _07864_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09243__A _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06807_ _13129_/A _09254_/A vssd1 vssd1 vccd1 vccd1 _12740_/A sky130_fd_sc_hd__xor2_4
X_07787_ _07851_/A _07851_/B vssd1 vssd1 vccd1 vccd1 _07787_/X sky130_fd_sc_hd__and2_1
XFILLER_0_78_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09526_ _09501_/A _11688_/B _09521_/Y hold245/A vssd1 vssd1 vccd1 vccd1 _09526_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_78_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09457_ _09455_/X _09456_/X _09674_/S vssd1 vssd1 vccd1 vccd1 _09457_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08408_ _08408_/A _08408_/B vssd1 vssd1 vccd1 vccd1 _08416_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__07698__A _10119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09388_ _09389_/A _09389_/B vssd1 vssd1 vccd1 vccd1 _09388_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_53_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12757__A1 _13129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08339_ _10263_/A _08339_/B vssd1 vssd1 vccd1 vccd1 _08406_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__09622__A1 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09622__B2 _08395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11350_ _11864_/A _09032_/X _09034_/C vssd1 vssd1 vccd1 vccd1 _11352_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10301_ _09988_/X _10297_/X _10300_/Y vssd1 vssd1 vccd1 vccd1 _10302_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_61_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11281_ _11281_/A _11281_/B vssd1 vssd1 vccd1 vccd1 _11288_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13020_ reg1_val[8] _13020_/B vssd1 vssd1 vccd1 vccd1 _13021_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13182__A1 wire101/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10232_ _10233_/A _10233_/B vssd1 vssd1 vccd1 vccd1 _10392_/B sky130_fd_sc_hd__nand2_1
X_10163_ _10734_/A _07007_/Y _07033_/X _10162_/Y vssd1 vssd1 vccd1 vccd1 _10165_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_100_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10094_ _10235_/A1 _07891_/X fanout10/X _10235_/B2 vssd1 vssd1 vccd1 vccd1 _10095_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11683__A _12525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12804_ _09694_/A curr_PC[1] _12825_/S vssd1 vssd1 vccd1 vccd1 _12806_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_69_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10996_ reg1_val[10] curr_PC[10] vssd1 vssd1 vccd1 vccd1 _10999_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _12735_/A1 _12732_/Y _12733_/X _09429_/X vssd1 vssd1 vccd1 vccd1 _12736_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_123_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _12666_/A _12666_/B vssd1 vssd1 vccd1 vccd1 _12670_/A sky130_fd_sc_hd__xnor2_1
X_11617_ _11617_/A _11617_/B vssd1 vssd1 vccd1 vccd1 _11618_/B sky130_fd_sc_hd__and2_1
XFILLER_0_115_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12597_ hold249/A _12786_/B1 _12653_/B _12596_/Y _12748_/B1 vssd1 vssd1 vccd1 vccd1
+ _12597_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_4_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12212__A3 _12372_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11548_ _11549_/A _11549_/B vssd1 vssd1 vccd1 vccd1 _11660_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_12_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11479_ reg1_val[14] _07527_/A _11586_/B vssd1 vssd1 vccd1 vccd1 _11479_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13218_ hold42/X hold273/A vssd1 vssd1 vccd1 vccd1 _13218_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_110_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _13149_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13149_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07710_ _07710_/A _07710_/B vssd1 vssd1 vccd1 vccd1 _07964_/B sky130_fd_sc_hd__xnor2_1
X_08690_ _08690_/A _08690_/B vssd1 vssd1 vccd1 vccd1 _08699_/B sky130_fd_sc_hd__xor2_4
XANTENNA__11487__B2 _11866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07641_ _07641_/A _07641_/B _07641_/C _07641_/D vssd1 vssd1 vccd1 vccd1 _07876_/A
+ sky130_fd_sc_hd__nand4_2
X_07572_ reg1_val[10] _11010_/A _07572_/S vssd1 vssd1 vccd1 vccd1 _07575_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_48_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09311_ _09311_/A _09311_/B vssd1 vssd1 vccd1 vccd1 _09313_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_75_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09242_ fanout24/X fanout76/X fanout74/X fanout23/X vssd1 vssd1 vccd1 vccd1 _09243_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10462__A2 _12793_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09173_ _10049_/A2 fanout21/X _08246_/B _09173_/B2 vssd1 vssd1 vccd1 vccd1 _09174_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_43_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08124_ _08123_/B _08123_/C _09949_/A vssd1 vssd1 vccd1 vccd1 _08125_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__07030__B _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11411__B2 _11281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06969__A2 _06936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08055_ _08113_/A _08113_/B _08050_/Y vssd1 vssd1 vccd1 vccd1 _08068_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__10672__A _11281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07006_ _06928_/A _06936_/B _13000_/B _07004_/X vssd1 vssd1 vccd1 vccd1 _07419_/A
+ sky130_fd_sc_hd__a31o_4
XANTENNA__13164__A1 wire122/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11175__B1 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07918__A1 _08118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07918__B2 fanout39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10922__B1 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ _09950_/A _09006_/B vssd1 vssd1 vccd1 vccd1 _09004_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13467__A2 _13555_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07908_ _07908_/A _07908_/B vssd1 vssd1 vccd1 vccd1 _07909_/B sky130_fd_sc_hd__xnor2_2
X_08888_ _08877_/A _08876_/C _08876_/B vssd1 vssd1 vccd1 vccd1 _08889_/C sky130_fd_sc_hd__a21o_1
X_07839_ _07968_/A _08028_/A _07968_/C vssd1 vssd1 vccd1 vccd1 _07969_/A sky130_fd_sc_hd__a21o_1
XANTENNA__13207__B _13207_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10850_ _10852_/A _10852_/B _10852_/C vssd1 vssd1 vccd1 vccd1 _10853_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09509_ _09509_/A _09520_/B vssd1 vssd1 vccd1 vccd1 _09509_/X sky130_fd_sc_hd__or2_4
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10781_ _10962_/A _10781_/B vssd1 vssd1 vccd1 vccd1 _10781_/X sky130_fd_sc_hd__or2_1
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ _12461_/A _12458_/Y _12460_/B vssd1 vssd1 vccd1 vccd1 _12524_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_109_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12451_ _07077_/X _12450_/X _12515_/S vssd1 vssd1 vccd1 vccd1 _12452_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11402_ _07198_/Y fanout15/X fanout31/X _12189_/A vssd1 vssd1 vccd1 vccd1 _11403_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07606__B1 _08806_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09847__S _10004_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10205__A2 _07477_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11402__A1 _07198_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12382_ _12382_/A _12382_/B vssd1 vssd1 vccd1 vccd1 _12382_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_105_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11402__B2 _12189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11333_ _11334_/A _11334_/B vssd1 vssd1 vccd1 vccd1 _11449_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09148__A _09949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11264_ curr_PC[12] _11382_/C vssd1 vssd1 vccd1 vccd1 _11264_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08052__A _10078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11166__B1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13003_ _13002_/A _12999_/Y _13001_/B vssd1 vssd1 vccd1 vccd1 _13007_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_30_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10215_ _10215_/A _10215_/B vssd1 vssd1 vccd1 vccd1 _10217_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_120_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11195_ _11195_/A _11195_/B vssd1 vssd1 vccd1 vccd1 _11202_/A sky130_fd_sc_hd__xnor2_1
X_10146_ _10148_/A _10148_/B vssd1 vssd1 vccd1 vccd1 _10146_/X sky130_fd_sc_hd__or2_1
XFILLER_0_27_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13458__A2 _13450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10077_ _08833_/B _10787_/B _10787_/C _07307_/Y fanout44/X vssd1 vssd1 vccd1 vccd1
+ _10078_/B sky130_fd_sc_hd__o32a_1
XANTENNA__12418__B1 _12667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap81 _11309_/A vssd1 vssd1 vccd1 vccd1 _13172_/A1 sky130_fd_sc_hd__buf_6
XFILLER_0_85_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10979_ _10981_/C _11106_/A vssd1 vssd1 vccd1 vccd1 _11227_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12718_ fanout5/X _12718_/B vssd1 vssd1 vccd1 vccd1 _12718_/Y sky130_fd_sc_hd__nor2_1
X_13698_ _13700_/CLK hold97/X vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12649_ _12648_/A _10022_/A _12648_/Y _09529_/B vssd1 vssd1 vccd1 vccd1 _12661_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_72_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08270__B1 _08328_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09860_ _09860_/A _09860_/B vssd1 vssd1 vccd1 vccd1 _09860_/Y sky130_fd_sc_hd__nand2_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10904__B1 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09492__S _09493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _08811_/A _08811_/B vssd1 vssd1 vccd1 vccd1 _08816_/B sky130_fd_sc_hd__xnor2_1
X_09791_ fanout21/X _07522_/Y _11423_/A _08246_/B vssd1 vssd1 vccd1 vccd1 _09792_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08742_ _08742_/A _08742_/B vssd1 vssd1 vccd1 vccd1 _08756_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12657__B1 _12657_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08673_ _08746_/A _08673_/B vssd1 vssd1 vccd1 vccd1 _08677_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout174_A _10236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07624_ _10050_/A _07624_/B vssd1 vssd1 vccd1 vccd1 _07628_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07555_ _11709_/A _07555_/B vssd1 vssd1 vccd1 vccd1 _07563_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06864__B _12981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07486_ _07486_/A _07486_/B _07486_/C _07486_/D vssd1 vssd1 vccd1 vccd1 _07493_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__08137__A _10236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09225_ _09225_/A _09225_/B vssd1 vssd1 vccd1 vccd1 _09297_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_8_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10986__A3 _10984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12882__A _13042_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09667__S _09674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09156_ reg1_val[29] _12656_/A _13129_/A vssd1 vssd1 vccd1 vccd1 _12754_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08107_ _08105_/Y _08998_/B _08035_/X vssd1 vssd1 vccd1 vccd1 _09001_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_71_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09087_ _09087_/A _09087_/B vssd1 vssd1 vccd1 vccd1 _09087_/X sky130_fd_sc_hd__and2_1
XANTENNA__08800__A2 _10522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08038_ _08038_/A _08038_/B vssd1 vssd1 vccd1 vccd1 _08101_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11148__B1 _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11010__B _12235_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10000_ _09670_/X _09682_/X _10004_/S vssd1 vssd1 vccd1 vccd1 _10000_/X sky130_fd_sc_hd__mux2_1
X_09989_ _09989_/A _10298_/A _09989_/C _10433_/A vssd1 vssd1 vccd1 vccd1 _09989_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__10123__A1 _09955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11951_ _11559_/B _11950_/X _11949_/Y vssd1 vssd1 vccd1 vccd1 _11952_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_98_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10902_ fanout34/X _07543_/X _07548_/X fanout32/X vssd1 vssd1 vccd1 vccd1 _10903_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_58_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11882_ _12058_/A _11969_/B hold259/A vssd1 vssd1 vccd1 vccd1 _11882_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10833_ _10832_/B _10832_/C _10832_/A vssd1 vssd1 vccd1 vccd1 _10834_/B sky130_fd_sc_hd__a21oi_1
X_13621_ _13717_/CLK _13621_/D vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10577__A _10577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11623__A1 _11997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10764_ _12825_/S _11020_/C vssd1 vssd1 vccd1 vccd1 _10764_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13552_ _13229_/X _13552_/B vssd1 vssd1 vccd1 vccd1 _13553_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__08047__A _10095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11623__B2 _11922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12503_ _12568_/B _12503_/B vssd1 vssd1 vccd1 vccd1 _12505_/C sky130_fd_sc_hd__or2_1
X_13483_ _13265_/X _13483_/B vssd1 vssd1 vccd1 vccd1 _13484_/B sky130_fd_sc_hd__nand2b_1
X_10695_ _10696_/A _10696_/B vssd1 vssd1 vccd1 vccd1 _10798_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07886__A _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12434_ _12435_/A _12435_/B vssd1 vssd1 vccd1 vccd1 _12505_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_23_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12365_ _12365_/A _12365_/B _12442_/A vssd1 vssd1 vccd1 vccd1 _12368_/C sky130_fd_sc_hd__or3_2
XFILLER_0_50_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11316_ _11438_/A _11316_/B vssd1 vssd1 vccd1 vccd1 _11318_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12296_ _12296_/A _12372_/D vssd1 vssd1 vccd1 vccd1 _12296_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11139__B1 _12657_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08004__B1 _08580_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11247_ _11244_/X _11246_/Y _12648_/A _11241_/X vssd1 vssd1 vccd1 vccd1 _11247_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_120_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11178_ _11709_/A _11178_/B vssd1 vssd1 vccd1 vccd1 _11182_/A sky130_fd_sc_hd__xnor2_2
X_10129_ _10130_/A _10130_/B vssd1 vssd1 vccd1 vccd1 _10129_/X sky130_fd_sc_hd__and2_1
XFILLER_0_89_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13562__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13603__A2 _13584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07340_ _07357_/A _07377_/A _07337_/B _07334_/D _07334_/B vssd1 vssd1 vccd1 vccd1
+ _07340_/X sky130_fd_sc_hd__a41o_1
XFILLER_0_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09283__A2 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07271_ reg1_val[6] _07572_/S vssd1 vssd1 vccd1 vccd1 _07271_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09010_ _09010_/A _09010_/B vssd1 vssd1 vccd1 vccd1 _10160_/C sky130_fd_sc_hd__xor2_2
XFILLER_0_72_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10934__B fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11917__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold102 hold102/A vssd1 vssd1 vccd1 vccd1 hold102/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold113 hold113/A vssd1 vssd1 vccd1 vccd1 hold113/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08794__A1 _08821_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold124 hold124/A vssd1 vssd1 vccd1 vccd1 hold124/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08794__B2 _08821_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold135 hold135/A vssd1 vssd1 vccd1 vccd1 hold135/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 hold146/A vssd1 vssd1 vccd1 vccd1 hold146/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 hold157/A vssd1 vssd1 vccd1 vccd1 hold157/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold168 hold168/A vssd1 vssd1 vccd1 vccd1 hold168/X sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ _09912_/A _09912_/B vssd1 vssd1 vccd1 vccd1 _09914_/B sky130_fd_sc_hd__xnor2_1
Xhold179 hold179/A vssd1 vssd1 vccd1 vccd1 hold179/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09843_ _09454_/X _09479_/X _10004_/S vssd1 vssd1 vccd1 vccd1 _09843_/X sky130_fd_sc_hd__mux2_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08420__A _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06887__A2_N _06980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _09774_/A _09774_/B vssd1 vssd1 vccd1 vccd1 _09775_/B sky130_fd_sc_hd__or2_1
X_06986_ reg1_val[6] _07556_/A vssd1 vssd1 vccd1 vccd1 _06986_/Y sky130_fd_sc_hd__nand2_1
X_08725_ _08725_/A _09051_/B vssd1 vssd1 vccd1 vccd1 _09046_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10105__A1 _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08656_ _08982_/A _08982_/B _08982_/C vssd1 vssd1 vccd1 vccd1 _08983_/A sky130_fd_sc_hd__a21oi_2
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09251__A _09371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07607_ _10078_/A _07607_/B vssd1 vssd1 vccd1 vccd1 _07671_/B sky130_fd_sc_hd__xor2_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ _08588_/A _08588_/B vssd1 vssd1 vccd1 vccd1 _08587_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_49_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07538_ _07517_/A _07517_/B _11076_/A _07537_/B _07537_/C vssd1 vssd1 vccd1 vccd1
+ _07538_/X sky130_fd_sc_hd__o2111a_2
XFILLER_0_48_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07469_ _07473_/A _07473_/B _11709_/A vssd1 vssd1 vccd1 vccd1 _11282_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_107_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09208_ _09825_/A _10435_/A vssd1 vssd1 vccd1 vccd1 _12743_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10480_ curr_PC[6] _10480_/B vssd1 vssd1 vccd1 vccd1 _10763_/C sky130_fd_sc_hd__and2_1
XFILLER_0_72_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11908__A2 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09139_ _09139_/A _09139_/B vssd1 vssd1 vccd1 vccd1 _09153_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11021__A _12825_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12150_ hold174/A _12311_/B1 _12227_/B _12533_/B1 vssd1 vssd1 vccd1 vccd1 _12151_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_114_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11101_ _11101_/A _11101_/B vssd1 vssd1 vccd1 vccd1 _11104_/C sky130_fd_sc_hd__xor2_1
X_12081_ _12082_/A _12082_/B vssd1 vssd1 vccd1 vccd1 _12173_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10860__A _11106_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08537__A1 _08866_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08537__B2 _09216_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11032_ _12421_/A _11032_/B vssd1 vssd1 vccd1 vccd1 _11041_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07760__A2 _08866_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12983_ _12987_/A _12983_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[0] sky130_fd_sc_hd__nor2_8
XANTENNA__09498__C1 _10603_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10647__A2 _07891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11934_ _11935_/A _11935_/B _11935_/C vssd1 vssd1 vccd1 vccd1 _12029_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09161__A _09161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11865_ _11864_/A _11864_/B _11864_/C _11864_/D vssd1 vssd1 vccd1 vccd1 _11866_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13604_ hold15/X _13597_/B hold143/X vssd1 vssd1 vccd1 vccd1 hold144/A sky130_fd_sc_hd__a21o_1
X_10816_ _07299_/Y _07422_/Y fanout70/X _07416_/X vssd1 vssd1 vccd1 vccd1 _10817_/B
+ sky130_fd_sc_hd__o22a_1
X_11796_ _11893_/B _11795_/Y _10342_/A vssd1 vssd1 vccd1 vccd1 _11796_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07276__A1 _10542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13535_ _13240_/X _13535_/B vssd1 vssd1 vccd1 vccd1 _13536_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_55_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10747_ _12056_/B _10748_/A hold163/A vssd1 vssd1 vccd1 vccd1 _10747_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_0_54_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_11_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10678_ _10679_/A _10679_/B _10679_/C vssd1 vssd1 vccd1 vccd1 _10838_/A sky130_fd_sc_hd__a21oi_2
X_13466_ hold264/X _13465_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13466_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12417_ _12417_/A _12417_/B vssd1 vssd1 vccd1 vccd1 _12423_/A sky130_fd_sc_hd__xnor2_1
X_13397_ hold5/X _13420_/B1 _07267_/X _13419_/A2 _13396_/Y vssd1 vssd1 vccd1 vccd1
+ hold6/A sky130_fd_sc_hd__o221a_1
XFILLER_0_23_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12348_ _12348_/A _12348_/B vssd1 vssd1 vccd1 vccd1 _12349_/B sky130_fd_sc_hd__or2_1
XFILLER_0_120_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11866__A _11866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10770__A _11708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12279_ _12280_/A _12280_/B vssd1 vssd1 vccd1 vccd1 _12362_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11585__B _12235_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13521__B2 _13542_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06840_ _06840_/A _06840_/B vssd1 vssd1 vccd1 vccd1 _12516_/A sky130_fd_sc_hd__nand2_1
X_06771_ instruction[19] instruction[12] _07135_/S vssd1 vssd1 vccd1 vccd1 reg1_idx[1]
+ sky130_fd_sc_hd__mux2_8
X_08510_ _08510_/A _08510_/B vssd1 vssd1 vccd1 vccd1 _08518_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09490_ reg1_val[5] reg1_val[26] _09493_/S vssd1 vssd1 vccd1 vccd1 _09490_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10638__A2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08441_ _08746_/A _08441_/B vssd1 vssd1 vccd1 vccd1 _08448_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11106__A _11106_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08372_ _08866_/B2 fanout76/X fanout74/X _08950_/B vssd1 vssd1 vccd1 vccd1 _08373_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11599__B1 _12867_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07323_ reg1_val[12] reg1_val[13] vssd1 vssd1 vccd1 vccd1 _07328_/C sky130_fd_sc_hd__or2_1
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout137_A _12695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13321__A _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07254_ _07287_/A _07254_/B _07254_/C vssd1 vssd1 vccd1 vccd1 _09254_/D sky130_fd_sc_hd__or3_4
XFILLER_0_26_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07185_ _07186_/B _07186_/C _07185_/C vssd1 vssd1 vccd1 vccd1 _07476_/C sky130_fd_sc_hd__and3_1
XANTENNA__08767__A1 _08806_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08767__B2 _08806_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10326__A1 _12314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09826_ _09426_/A _09426_/B _09650_/A _09650_/B vssd1 vssd1 vccd1 vccd1 _09826_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12079__A1 _12557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ _10537_/A _09757_/B vssd1 vssd1 vccd1 vccd1 _09765_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12079__B2 _12557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06969_ _06928_/A _06936_/B _13025_/B _06967_/X vssd1 vssd1 vccd1 vccd1 _07449_/A
+ sky130_fd_sc_hd__a31oi_4
X_08708_ _09371_/A _08708_/B vssd1 vssd1 vccd1 vccd1 _08744_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11826__A1 _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09688_ _09490_/X _09492_/X _09688_/S vssd1 vssd1 vccd1 vccd1 _09688_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11826__B2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _10944_/A _08640_/B vssd1 vssd1 vccd1 vccd1 _08639_/Y sky130_fd_sc_hd__nand2_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _11650_/A _11650_/B vssd1 vssd1 vccd1 vccd1 _11652_/B sky130_fd_sc_hd__xnor2_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout30 _07421_/X vssd1 vssd1 vccd1 vccd1 _07833_/B sky130_fd_sc_hd__buf_6
XFILLER_0_76_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout41 _07289_/X vssd1 vssd1 vccd1 vccd1 _12087_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07258__A1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10601_ _11575_/S _10601_/B _10601_/C vssd1 vssd1 vccd1 vccd1 _10601_/X sky130_fd_sc_hd__and3_1
Xfanout52 _07217_/Y vssd1 vssd1 vccd1 vccd1 _12557_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__07258__B2 _08328_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout63 _09265_/Y vssd1 vssd1 vccd1 vccd1 _10518_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__11054__A2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11581_ _12058_/A _11881_/D hold296/A vssd1 vssd1 vccd1 vccd1 _11581_/Y sky130_fd_sc_hd__a21oi_1
Xfanout74 _07543_/X vssd1 vssd1 vccd1 vccd1 fanout74/X sky130_fd_sc_hd__buf_8
XANTENNA__10855__A _10981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout85 _07478_/Y vssd1 vssd1 vccd1 vccd1 fanout85/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10262__B1 _07453_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout96 _12094_/A vssd1 vssd1 vccd1 vccd1 _10266_/A sky130_fd_sc_hd__clkbuf_16
X_13320_ hold188/X _13463_/B2 _13450_/B _13642_/Q vssd1 vssd1 vccd1 vccd1 hold189/A
+ sky130_fd_sc_hd__a22o_1
X_10532_ _10533_/A _10533_/B vssd1 vssd1 vccd1 vccd1 _10679_/B sky130_fd_sc_hd__or2_1
XANTENNA__08207__B1 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10463_ hold294/A hold283/A _10463_/C vssd1 vssd1 vccd1 vccd1 _10610_/B sky130_fd_sc_hd__or3_2
X_13251_ hold90/X hold251/X vssd1 vssd1 vccd1 vccd1 _13251_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_60_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12202_ _12202_/A vssd1 vssd1 vccd1 vccd1 _12365_/A sky130_fd_sc_hd__inv_2
X_13182_ wire101/X _13194_/A2 hold38/X _13539_/A vssd1 vssd1 vccd1 vccd1 _13627_/D
+ sky130_fd_sc_hd__o211a_1
X_10394_ _10395_/B _10395_/A vssd1 vssd1 vccd1 vccd1 _10394_/X sky130_fd_sc_hd__and2b_1
X_12133_ _12046_/A _12044_/X _06869_/B vssd1 vssd1 vccd1 vccd1 _12133_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_102_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07981__A2 _11922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09707__B1 _12796_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12064_ _07349_/X _07481_/X _12235_/C _12063_/X vssd1 vssd1 vccd1 vccd1 _12064_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08060__A _10239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11015_ _10603_/S _10319_/X _09537_/B vssd1 vssd1 vccd1 vccd1 _12143_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_max_cap102_A _07300_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12966_ _12979_/A _12967_/B vssd1 vssd1 vccd1 vccd1 _12968_/A sky130_fd_sc_hd__and2_1
XFILLER_0_87_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11917_ _07198_/Y fanout8/X fanout3/X _11997_/A vssd1 vssd1 vccd1 vccd1 _11918_/B
+ sky130_fd_sc_hd__a22o_1
X_12897_ _13054_/B _12897_/B vssd1 vssd1 vccd1 vccd1 _12898_/B sky130_fd_sc_hd__or2_1
XFILLER_0_28_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11848_ _11944_/A _11848_/B vssd1 vssd1 vccd1 vccd1 _11851_/A sky130_fd_sc_hd__nand2_1
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07249__A1 _08821_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07249__B2 _08821_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11779_ _11779_/A _11779_/B vssd1 vssd1 vccd1 vccd1 _11779_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_82_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13141__A _13141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12793__A2 _12793_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13518_ _13251_/X _13518_/B vssd1 vssd1 vccd1 vccd1 _13519_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_82_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13449_ _13547_/A hold246/X vssd1 vssd1 vccd1 vccd1 _13705_/D sky130_fd_sc_hd__and2_1
XFILLER_0_113_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08990_ _08990_/A _08990_/B vssd1 vssd1 vccd1 vccd1 _09003_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_11_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07941_ _09190_/A _07941_/B vssd1 vssd1 vccd1 vccd1 _07943_/B sky130_fd_sc_hd__or2_2
X_07872_ _07872_/A _07872_/B vssd1 vssd1 vccd1 vccd1 _07873_/B sky130_fd_sc_hd__nor2_2
XANTENNA__08921__A1 _07238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09611_ _09726_/B _09611_/B _09611_/C vssd1 vssd1 vccd1 vccd1 _09812_/A sky130_fd_sc_hd__and3_1
XANTENNA__08921__B2 _07239_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06823_ _06824_/A _06824_/B vssd1 vssd1 vccd1 vccd1 _06848_/D sky130_fd_sc_hd__and2_1
XFILLER_0_92_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09542_ curr_PC[0] _12825_/S vssd1 vssd1 vccd1 vccd1 _09542_/X sky130_fd_sc_hd__or2_1
X_06754_ reg1_val[20] vssd1 vssd1 vccd1 vccd1 _07483_/A sky130_fd_sc_hd__inv_2
XANTENNA__11808__A1 _12557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11808__B2 _07597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07314__A _10078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13035__B _13036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09473_ _09469_/X _09472_/X _10005_/S vssd1 vssd1 vccd1 vccd1 _09473_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_66_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout254_A _13141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08424_ _08271_/A _07544_/Y _11638_/A _09501_/A vssd1 vssd1 vccd1 vccd1 _08425_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10492__B1 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08355_ _08355_/A _08355_/B vssd1 vssd1 vccd1 vccd1 _08368_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13430__B1 _13444_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07306_ _10537_/A _07312_/B vssd1 vssd1 vccd1 vccd1 _07306_/X sky130_fd_sc_hd__and2b_1
X_08286_ _08286_/A _08286_/B vssd1 vssd1 vccd1 vccd1 _08287_/B sky130_fd_sc_hd__and2_1
XFILLER_0_61_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08145__A _11286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07237_ _09371_/A _07240_/A _07236_/X vssd1 vssd1 vccd1 vccd1 _07237_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__07660__A1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07660__B2 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12890__A _13048_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07984__A _09950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07168_ reg1_val[4] _07265_/D vssd1 vssd1 vccd1 vccd1 _07168_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_112_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07099_ _07099_/A _07099_/B _07099_/C vssd1 vssd1 vccd1 vccd1 _07099_/X sky130_fd_sc_hd__or3_1
XFILLER_0_100_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout220 _07363_/B vssd1 vssd1 vccd1 vccd1 _11576_/A sky130_fd_sc_hd__clkbuf_8
Xfanout231 _11688_/B vssd1 vssd1 vccd1 vccd1 _12657_/B1 sky130_fd_sc_hd__buf_4
Xfanout242 _12406_/B1 vssd1 vssd1 vccd1 vccd1 _10342_/A sky130_fd_sc_hd__buf_8
Xfanout253 _13141_/A vssd1 vssd1 vccd1 vccd1 _13563_/B2 sky130_fd_sc_hd__clkbuf_4
Xfanout264 _13082_/A vssd1 vssd1 vccd1 vccd1 _13129_/B sky130_fd_sc_hd__buf_8
Xfanout275 _13444_/C1 vssd1 vssd1 vccd1 vccd1 _13539_/A sky130_fd_sc_hd__clkbuf_4
Xfanout286 _06748_/Y vssd1 vssd1 vccd1 vccd1 _08328_/B2 sky130_fd_sc_hd__clkbuf_4
X_09809_ _09635_/A _09635_/B _09634_/A vssd1 vssd1 vccd1 vccd1 _09819_/A sky130_fd_sc_hd__a21o_2
Xfanout297 instruction[6] vssd1 vssd1 vccd1 vccd1 _13744_/A sky130_fd_sc_hd__clkbuf_8
X_12820_ _12995_/B _12820_/B vssd1 vssd1 vccd1 vccd1 _12821_/B sky130_fd_sc_hd__or2_1
XANTENNA__07479__A1 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07479__B2 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _12374_/A _12750_/X hold224/A vssd1 vssd1 vccd1 vccd1 _12753_/A sky130_fd_sc_hd__a21oi_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _12406_/B1 _11699_/X _11700_/X _11701_/Y vssd1 vssd1 vccd1 vccd1 dest_val[16]
+ sky130_fd_sc_hd__a2bb2o_4
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _12127_/B _12682_/B _12682_/C _12682_/D vssd1 vssd1 vccd1 vccd1 _12686_/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _11633_/A _11633_/B vssd1 vssd1 vccd1 vccd1 _11642_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10235__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11564_ _09048_/B _11562_/X _11563_/Y vssd1 vssd1 vccd1 vccd1 _11564_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_25_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11983__B1 _11982_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13303_ _13239_/B _13540_/B _13237_/X vssd1 vssd1 vccd1 vccd1 _13544_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_24_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10515_ _10515_/A _10515_/B _10515_/C vssd1 vssd1 vccd1 vccd1 _10516_/B sky130_fd_sc_hd__and3_1
XFILLER_0_107_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11495_ _12087_/A fanout34/X fanout32/X _12103_/A vssd1 vssd1 vccd1 vccd1 _11496_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07894__A _08907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10446_ _06994_/A _07003_/B _10308_/X _06996_/B vssd1 vssd1 vccd1 vccd1 _10589_/B
+ sky130_fd_sc_hd__a31oi_1
X_13234_ hold85/X hold275/A vssd1 vssd1 vccd1 vccd1 _13236_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_0_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10377_ _11719_/A _10377_/B vssd1 vssd1 vccd1 vccd1 _10379_/B sky130_fd_sc_hd__xnor2_2
X_13165_ hold105/X _13191_/B vssd1 vssd1 vccd1 vccd1 hold106/A sky130_fd_sc_hd__or2_1
XFILLER_0_20_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12116_ _12117_/A _12117_/B vssd1 vssd1 vccd1 vccd1 _12203_/B sky130_fd_sc_hd__nand2_1
X_13096_ _13093_/A _13095_/B _13093_/B vssd1 vssd1 vccd1 vccd1 _13098_/A sky130_fd_sc_hd__a21bo_1
X_12047_ _12046_/A _12046_/B _12046_/Y _12047_/C1 vssd1 vssd1 vccd1 vccd1 _12047_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07118__B _07118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12463__A1 _12782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12949_ _12947_/X _12949_/B vssd1 vssd1 vccd1 vccd1 _12961_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_87_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08419__B1 _08486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07890__A1 _07521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08140_ _08140_/A _08140_/B vssd1 vssd1 vccd1 vccd1 _08176_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10226__B1 _07877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11974__B1 _12533_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08071_ _08071_/A _08071_/B vssd1 vssd1 vccd1 vccd1 _08088_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_70_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09495__S _10007_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07022_ _09694_/A _10007_/S vssd1 vssd1 vccd1 vccd1 _07022_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13176__C1 _13543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08973_ _08974_/A _08973_/B vssd1 vssd1 vccd1 vccd1 _09023_/B sky130_fd_sc_hd__and2_1
XANTENNA__09147__A1 _08271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09147__B2 _09501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ _07924_/A _07924_/B vssd1 vssd1 vccd1 vccd1 _07925_/B sky130_fd_sc_hd__nand2_1
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
X_07855_ fanout28/X _10915_/A _11047_/A _08395_/B vssd1 vssd1 vccd1 vccd1 _07856_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06867__B _07201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06806_ _09254_/A vssd1 vssd1 vccd1 vccd1 _09146_/A sky130_fd_sc_hd__inv_2
X_07786_ _07786_/A _07786_/B vssd1 vssd1 vccd1 vccd1 _07851_/B sky130_fd_sc_hd__xnor2_2
X_09525_ _13744_/A instruction[5] _09525_/C vssd1 vssd1 vccd1 vccd1 _09525_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__13480__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10465__B1 _12796_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09456_ reg1_val[12] reg1_val[19] _09463_/S vssd1 vssd1 vccd1 vccd1 _09456_/X sky130_fd_sc_hd__mux2_1
X_08407_ _08405_/B _08472_/B _08405_/A vssd1 vssd1 vccd1 vccd1 _08416_/A sky130_fd_sc_hd__a21bo_2
X_09387_ _09387_/A _09387_/B vssd1 vssd1 vccd1 vccd1 _09389_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_46_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12757__A2 _09254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08338_ _09671_/S fanout28/X _08395_/B _08873_/B2 vssd1 vssd1 vccd1 vccd1 _08339_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_46_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09622__A2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08269_ _09948_/A _08269_/B vssd1 vssd1 vccd1 vccd1 _08274_/A sky130_fd_sc_hd__xnor2_1
X_10300_ _09983_/X _10146_/X _10147_/X vssd1 vssd1 vccd1 vccd1 _10300_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11280_ fanout83/X fanout10/X fanout5/X _08580_/B vssd1 vssd1 vccd1 vccd1 _11281_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_14_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10231_ _11825_/A _10231_/B vssd1 vssd1 vccd1 vccd1 _10233_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13182__A2 _13194_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07219__A _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10162_ _07010_/B _10161_/X _10734_/A vssd1 vssd1 vccd1 vccd1 _10162_/Y sky130_fd_sc_hd__a21oi_1
X_10093_ _10093_/A _10093_/B vssd1 vssd1 vccd1 vccd1 _10100_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09153__B _09153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12803_ _12809_/A _12803_/B vssd1 vssd1 vccd1 vccd1 new_PC[0] sky130_fd_sc_hd__and2_4
X_10995_ reg1_val[10] curr_PC[10] vssd1 vssd1 vccd1 vccd1 _10995_/X sky130_fd_sc_hd__and2_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12734_ _12735_/A1 _12733_/X _12732_/Y vssd1 vssd1 vccd1 vccd1 _12736_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06793__A _13135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ fanout8/X fanout7/X fanout3/X _09145_/Y vssd1 vssd1 vccd1 vccd1 _12666_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11616_ _11617_/A _11617_/B vssd1 vssd1 vccd1 vccd1 _11712_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10759__A1 _12537_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12596_ _12786_/B1 _12653_/B hold249/A vssd1 vssd1 vccd1 vccd1 _12596_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10759__B2 _12710_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08821__B1 _08923_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11547_ _11441_/A _11441_/B _11442_/Y vssd1 vssd1 vccd1 vccd1 _11549_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11478_ hold193/A _11478_/B vssd1 vssd1 vccd1 vccd1 _11478_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13217_ _13579_/B _13217_/B vssd1 vssd1 vccd1 vccd1 _13311_/B sky130_fd_sc_hd__nor2_1
X_10429_ _10429_/A _10429_/B vssd1 vssd1 vccd1 vccd1 _10432_/B sky130_fd_sc_hd__xnor2_4
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ hold11/X _13193_/B _13147_/Y _13459_/A vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__o211a_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ _13079_/A _13081_/D vssd1 vssd1 vccd1 vccd1 loadstore_address[19] sky130_fd_sc_hd__xnor2_4
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07640_ _07641_/A _07641_/B _07641_/C _07641_/D vssd1 vssd1 vccd1 vccd1 _07642_/A
+ sky130_fd_sc_hd__a22o_1
X_07571_ _07571_/A _07571_/B vssd1 vssd1 vccd1 vccd1 _11010_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_87_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09310_ _09310_/A _09310_/B vssd1 vssd1 vccd1 vccd1 _09311_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_48_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09241_ _10944_/A _09241_/B vssd1 vssd1 vccd1 vccd1 _09248_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09172_ _11507_/A _09172_/B vssd1 vssd1 vccd1 vccd1 _09176_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08123_ _09949_/A _08123_/B _08123_/C vssd1 vssd1 vccd1 vccd1 _08125_/B sky130_fd_sc_hd__and3_1
XFILLER_0_22_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11411__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout217_A _09496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08054_ _08054_/A _08054_/B vssd1 vssd1 vccd1 vccd1 _08113_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06969__A3 _13025_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08423__A _08951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07005_ _06928_/A _06936_/B _13000_/B _07004_/X vssd1 vssd1 vccd1 vccd1 _10457_/S
+ sky130_fd_sc_hd__a31oi_4
XFILLER_0_101_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13164__A2 _13194_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11175__A1 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11175__B2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07918__A2 _07491_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10922__A1 _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10922__B2 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13475__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ _09659_/A _09660_/A vssd1 vssd1 vccd1 vccd1 _09006_/B sky130_fd_sc_hd__and2_1
XANTENNA__09254__A _09254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07907_ _07908_/A _07908_/B vssd1 vssd1 vccd1 vccd1 _07907_/Y sky130_fd_sc_hd__nand2_1
X_08887_ _08887_/A _08887_/B vssd1 vssd1 vccd1 vccd1 _08889_/B sky130_fd_sc_hd__xnor2_1
X_07838_ _07838_/A _07838_/B vssd1 vssd1 vccd1 vccd1 _07968_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__11883__C1 _12748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07769_ _07970_/A _07970_/B _07766_/C vssd1 vssd1 vccd1 vccd1 _07770_/C sky130_fd_sc_hd__a21oi_1
X_09508_ _09509_/A _09520_/B vssd1 vssd1 vccd1 vccd1 _09508_/Y sky130_fd_sc_hd__nor2_1
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10780_ _10780_/A _10780_/B _10780_/C vssd1 vssd1 vccd1 vccd1 _10781_/B sky130_fd_sc_hd__and3_1
XANTENNA_fanout32_A _07699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _09688_/S _09436_/X _09438_/Y _10005_/S vssd1 vssd1 vccd1 vccd1 _09439_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07221__B _07521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12450_ _12382_/A _12380_/X _06847_/B vssd1 vssd1 vccd1 vccd1 _12450_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_124_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11401_ _11401_/A _11401_/B vssd1 vssd1 vccd1 vccd1 _11417_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07606__A1 _10536_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07606__B2 _11922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12381_ _07059_/X _12380_/X _12515_/S vssd1 vssd1 vccd1 vccd1 _12382_/B sky130_fd_sc_hd__mux2_1
XANTENNA__11402__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_80 reg1_val[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11332_ _11332_/A _11332_/B vssd1 vssd1 vccd1 vccd1 _11334_/B sky130_fd_sc_hd__xor2_1
X_11263_ _10730_/B _11230_/X _11231_/Y _11262_/X vssd1 vssd1 vccd1 vccd1 _11263_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11166__A1 _11732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11166__B2 _07310_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13002_ _13002_/A _13002_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[4] sky130_fd_sc_hd__xnor2_4
X_10214_ _10215_/B vssd1 vssd1 vccd1 vccd1 _10214_/Y sky130_fd_sc_hd__inv_2
X_11194_ _11195_/A _11195_/B vssd1 vssd1 vccd1 vccd1 _11326_/B sky130_fd_sc_hd__and2b_1
X_10145_ _10145_/A _10145_/B vssd1 vssd1 vccd1 vccd1 _10148_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__07385__A3 _07634_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10076_ _10507_/A _10076_/B vssd1 vssd1 vccd1 vccd1 _10080_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09531__A1 _10007_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07542__B1 _07521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12418__A1 _12614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12418__B2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10978_ _10721_/Y _10851_/X _10853_/B vssd1 vssd1 vccd1 vccd1 _10978_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_128_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07412__A _12253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12717_ _12717_/A fanout5/X vssd1 vssd1 vccd1 vccd1 _12717_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_85_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13697_ _13700_/CLK _13697_/D vssd1 vssd1 vccd1 vccd1 hold130/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12648_ _12648_/A _12648_/B vssd1 vssd1 vccd1 vccd1 _12648_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_53_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12579_ _12516_/A _12514_/Y _06840_/A vssd1 vssd1 vccd1 vccd1 _12579_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13146__A2 _13193_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10904__A1 _13180_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10904__B2 wire101/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08810_ _08845_/A _08845_/B vssd1 vssd1 vccd1 vccd1 _08846_/A sky130_fd_sc_hd__and2_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _09557_/A _09556_/Y _09554_/Y vssd1 vssd1 vccd1 vccd1 _09804_/A sky130_fd_sc_hd__a21bo_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08741_ _08766_/A _08766_/B _08755_/A vssd1 vssd1 vccd1 vccd1 _08756_/A sky130_fd_sc_hd__o21ai_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08672_ _13149_/A _10538_/A _08778_/B _08923_/B1 vssd1 vssd1 vccd1 vccd1 _08673_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07623_ fanout35/X _08873_/B2 _07699_/B _13149_/A vssd1 vssd1 vccd1 vccd1 _07624_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07025__C _07025_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13606__B1 _13568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10948__A _11709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07554_ _10915_/A fanout24/X _07471_/Y _08486_/B vssd1 vssd1 vccd1 vccd1 _07555_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_75_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07485_ _07486_/A _07486_/B _07486_/C _07486_/D vssd1 vssd1 vccd1 vccd1 _11991_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09224_ _09225_/B _09225_/A vssd1 vssd1 vccd1 vccd1 _09224_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_91_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13385__A2 _13444_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09155_ reg1_val[29] _13129_/A _12656_/A vssd1 vssd1 vccd1 vccd1 _12754_/A sky130_fd_sc_hd__or3_4
XFILLER_0_90_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08106_ _08999_/A _08999_/B vssd1 vssd1 vccd1 vccd1 _08998_/B sky130_fd_sc_hd__or2_1
XANTENNA__07468__S _11709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09086_ _09092_/A _09086_/B _09086_/C vssd1 vssd1 vccd1 vccd1 _09087_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_114_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08037_ _08037_/A _08037_/B vssd1 vssd1 vccd1 vccd1 _08101_/A sky130_fd_sc_hd__and2_1
XFILLER_0_102_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11699__A2 _11793_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ _09824_/A _09824_/B _09987_/Y vssd1 vssd1 vccd1 vccd1 _09988_/X sky130_fd_sc_hd__a21bo_1
X_08939_ _09161_/A _07238_/X _07239_/Y _07399_/Y vssd1 vssd1 vccd1 vccd1 _08940_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10659__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11950_ _11950_/A _12125_/B vssd1 vssd1 vccd1 vccd1 _11950_/X sky130_fd_sc_hd__and2_1
XANTENNA__10123__A2 _10518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10901_ _10843_/A _10843_/B _10844_/Y vssd1 vssd1 vccd1 vccd1 _10974_/A sky130_fd_sc_hd__o21ai_1
X_11881_ hold257/A hold292/A hold296/A _11881_/D vssd1 vssd1 vccd1 vccd1 _11969_/B
+ sky130_fd_sc_hd__or4_1
X_13620_ _13717_/CLK _13620_/D vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__dfxtp_1
X_10832_ _10832_/A _10832_/B _10832_/C vssd1 vssd1 vccd1 vccd1 _10834_/A sky130_fd_sc_hd__and3_1
XANTENNA__10577__B _10631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07232__A _07572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13551_ _13591_/A hold256/X vssd1 vssd1 vccd1 vccd1 _13727_/D sky130_fd_sc_hd__and2_1
X_10763_ curr_PC[7] curr_PC[8] _10763_/C vssd1 vssd1 vccd1 vccd1 _11020_/C sky130_fd_sc_hd__and3_2
XANTENNA__11623__A2 _07643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12502_ _12502_/A _12502_/B _12502_/C vssd1 vssd1 vccd1 vccd1 _12503_/B sky130_fd_sc_hd__nor3_1
X_13482_ _13591_/A hold277/X vssd1 vssd1 vccd1 vccd1 _13712_/D sky130_fd_sc_hd__and2_1
XFILLER_0_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10694_ _12094_/A _10694_/B vssd1 vssd1 vccd1 vccd1 _10696_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12433_ _12353_/A _12352_/B _12352_/A vssd1 vssd1 vccd1 vccd1 _12435_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_120_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12364_ _12202_/A _12288_/A _12287_/A vssd1 vssd1 vccd1 vccd1 _12364_/X sky130_fd_sc_hd__a21o_1
X_11315_ _11315_/A _11315_/B _11315_/C vssd1 vssd1 vccd1 vccd1 _11316_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_105_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12295_ _12442_/A _12295_/B vssd1 vssd1 vccd1 vccd1 _12372_/D sky130_fd_sc_hd__xnor2_4
XFILLER_0_50_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11139__B2 _11126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08004__A1 _09885_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08004__B2 _10049_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11246_ _12525_/A _11246_/B vssd1 vssd1 vccd1 vccd1 _11246_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_max_cap81_A _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11177_ fanout23/X _10787_/B _10787_/C fanout25/X _12557_/B vssd1 vssd1 vccd1 vccd1
+ _11178_/B sky130_fd_sc_hd__o32a_1
XANTENNA__07407__A _09496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10128_ _10128_/A _10128_/B vssd1 vssd1 vccd1 vccd1 _10130_/B sky130_fd_sc_hd__nor2_2
X_10059_ _10060_/A _10060_/B _10060_/C vssd1 vssd1 vccd1 vccd1 _10282_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__07126__B _07129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11614__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07270_ _07320_/C _07270_/B vssd1 vssd1 vccd1 vccd1 _07270_/X sky130_fd_sc_hd__and2_1
XFILLER_0_57_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11378__B2 _09493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold103 hold103/A vssd1 vssd1 vccd1 vccd1 hold103/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 hold114/A vssd1 vssd1 vccd1 vccd1 hold114/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08794__A2 _08866_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold125 hold125/A vssd1 vssd1 vccd1 vccd1 hold125/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold136 hold136/A vssd1 vssd1 vccd1 vccd1 hold136/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 hold147/A vssd1 vssd1 vccd1 vccd1 hold147/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 hold158/A vssd1 vssd1 vccd1 vccd1 hold158/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09911_ _09912_/A _09912_/B vssd1 vssd1 vccd1 vccd1 _10134_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_111_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold169 hold169/A vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09842_ _09840_/X _09841_/X _10600_/S vssd1 vssd1 vccd1 vccd1 _09842_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13319__A _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _09774_/A _09774_/B vssd1 vssd1 vccd1 vccd1 _09773_/X sky130_fd_sc_hd__and2_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06985_ reg1_val[6] _07556_/A vssd1 vssd1 vccd1 vccd1 _10589_/A sky130_fd_sc_hd__and2_1
X_08724_ _08724_/A _08724_/B vssd1 vssd1 vccd1 vccd1 _08724_/X sky130_fd_sc_hd__xor2_1
X_08655_ _08655_/A _08655_/B vssd1 vssd1 vccd1 vccd1 _08982_/C sky130_fd_sc_hd__xor2_1
XANTENNA__06875__B _06875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07606_ _10536_/A1 wire101/A _08806_/B1 _11922_/A vssd1 vssd1 vccd1 vccd1 _07607_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08586_ _09659_/B _08586_/B vssd1 vssd1 vccd1 vccd1 _08588_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_49_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07537_ _11076_/A _07537_/B _07537_/C vssd1 vssd1 vccd1 vccd1 _07546_/A sky130_fd_sc_hd__and3_1
XFILLER_0_63_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07987__A _09371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09678__S _09703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07468_ _07474_/A _07474_/B _11709_/A vssd1 vssd1 vccd1 vccd1 _07468_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09207_ _09094_/B _09205_/X _09206_/X _09092_/X _09204_/X vssd1 vssd1 vccd1 vccd1
+ _10435_/A sky130_fd_sc_hd__o221a_2
XANTENNA__13358__A2 _13463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07399_ _10007_/S _07400_/B vssd1 vssd1 vccd1 vccd1 _07399_/Y sky130_fd_sc_hd__xnor2_4
X_09138_ _09139_/A _09139_/B vssd1 vssd1 vccd1 vccd1 _09138_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09431__B1 _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09069_ _09060_/B _09060_/C _09068_/X vssd1 vssd1 vccd1 vccd1 _09071_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12832__S _12867_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11100_ _11101_/B _11101_/A vssd1 vssd1 vccd1 vccd1 _11222_/B sky130_fd_sc_hd__nand2b_1
X_12080_ _12417_/A _12080_/B vssd1 vssd1 vccd1 vccd1 _12082_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08537__A2 _10538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11031_ wire101/X fanout14/X fanout31/X _11922_/A vssd1 vssd1 vccd1 vccd1 _11032_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09426__B _09426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12982_ _12982_/A _12982_/B vssd1 vssd1 vccd1 vccd1 _12983_/B sky130_fd_sc_hd__nor2_2
X_11933_ _11933_/A _11933_/B vssd1 vssd1 vccd1 vccd1 _11935_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__10588__A _10734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09161__B fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11864_ _11864_/A _11864_/B _11864_/C _11864_/D vssd1 vssd1 vccd1 vccd1 _11864_/X
+ sky130_fd_sc_hd__and4_1
X_13603_ hold143/X _13584_/B hold192/A _13599_/D vssd1 vssd1 vccd1 vccd1 _13605_/B
+ sky130_fd_sc_hd__a22o_1
X_10815_ _12252_/A _10815_/B vssd1 vssd1 vccd1 vccd1 _10823_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11795_ curr_PC[16] _11794_/C curr_PC[17] vssd1 vssd1 vccd1 vccd1 _11795_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10804__B1 _07543_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13534_ _13539_/A hold260/X vssd1 vssd1 vccd1 vccd1 _13723_/D sky130_fd_sc_hd__and2_1
X_10746_ hold180/A _10882_/C vssd1 vssd1 vccd1 vccd1 _10748_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13465_ _13465_/A _13465_/B vssd1 vssd1 vccd1 vccd1 _13465_/Y sky130_fd_sc_hd__xnor2_1
X_10677_ _10811_/A _10677_/B vssd1 vssd1 vccd1 vccd1 _10679_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_23_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07028__A2 _06928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12416_ fanout35/X fanout10/X fanout5/X _07401_/Y vssd1 vssd1 vccd1 vccd1 _12417_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13396_ _06743_/Y _13141_/A rst vssd1 vssd1 vccd1 vccd1 _13396_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10032__A1 _12314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12347_ _12348_/A _12348_/B vssd1 vssd1 vccd1 vccd1 _12426_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_49_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12278_ _12278_/A _12278_/B vssd1 vssd1 vccd1 vccd1 _12280_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13139__A _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11229_ _11452_/A _11229_/B vssd1 vssd1 vccd1 vccd1 _11600_/A sky130_fd_sc_hd__xor2_4
XANTENNA__13521__A2 _13555_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06770_ instruction[18] instruction[11] _07135_/S vssd1 vssd1 vccd1 vccd1 reg1_idx[0]
+ sky130_fd_sc_hd__mux2_8
XFILLER_0_65_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11296__B1 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08440_ _08868_/B1 _10538_/A _08778_/B _10522_/A vssd1 vssd1 vccd1 vccd1 _08441_/B
+ sky130_fd_sc_hd__o22a_1
X_08371_ _08371_/A _08371_/B vssd1 vssd1 vccd1 vccd1 _08408_/A sky130_fd_sc_hd__xor2_4
XANTENNA__11106__B _11225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07322_ reg1_val[12] reg1_val[13] vssd1 vssd1 vccd1 vccd1 _07324_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_45_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07253_ _07287_/A _07254_/B _07254_/C vssd1 vssd1 vccd1 vccd1 _07595_/A sky130_fd_sc_hd__nor3_4
XANTENNA__12548__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07184_ _07472_/A _07455_/A _10889_/A _07184_/D vssd1 vssd1 vccd1 vccd1 _07185_/C
+ sky130_fd_sc_hd__nor4_1
XFILLER_0_41_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10023__A1 _12537_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08767__A2 _07399_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10023__B2 _12759_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09825_ _09825_/A _09986_/A _10150_/A _10298_/A vssd1 vssd1 vccd1 vccd1 _10435_/B
+ sky130_fd_sc_hd__or4_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09756_ _12413_/A _10536_/A1 _10536_/B2 _12496_/A vssd1 vssd1 vccd1 vccd1 _09757_/B
+ sky130_fd_sc_hd__a22o_1
X_06968_ _06928_/A _06936_/B _13025_/B _06967_/X vssd1 vssd1 vccd1 vccd1 _07184_/D
+ sky130_fd_sc_hd__a31o_2
XANTENNA__06886__A _06886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12079__A2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08707_ _07239_/Y wire122/A _10637_/A _07238_/X vssd1 vssd1 vccd1 vccd1 _08708_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11287__B1 _11286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09687_ _09486_/X _09489_/X _09688_/S vssd1 vssd1 vccd1 vccd1 _09687_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11826__A2 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06899_ reg1_val[17] _11793_/A vssd1 vssd1 vccd1 vccd1 _11867_/B sky130_fd_sc_hd__nand2_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _08686_/A _08686_/B _08634_/Y vssd1 vssd1 vccd1 vccd1 _08662_/A sky130_fd_sc_hd__o21ai_4
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08569_ _08569_/A _08569_/B vssd1 vssd1 vccd1 vccd1 _09068_/B sky130_fd_sc_hd__xnor2_1
Xfanout20 fanout21/X vssd1 vssd1 vccd1 vccd1 fanout20/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout31 _07421_/X vssd1 vssd1 vccd1 vccd1 fanout31/X sky130_fd_sc_hd__buf_4
Xfanout42 _07282_/X vssd1 vssd1 vccd1 vccd1 fanout42/X sky130_fd_sc_hd__buf_8
X_10600_ _10004_/X _10007_/X _10600_/S vssd1 vssd1 vccd1 vccd1 _10600_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13512__A _13543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07258__A2 _08907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout53 _07204_/Y vssd1 vssd1 vccd1 vccd1 fanout53/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_64_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11580_ hold296/A _12058_/A _11881_/D vssd1 vssd1 vccd1 vccd1 _11580_/X sky130_fd_sc_hd__and3_1
XFILLER_0_119_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout64 _11731_/A vssd1 vssd1 vccd1 vccd1 _12668_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_107_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10855__B _10981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout75 _10787_/A vssd1 vssd1 vccd1 vccd1 fanout75/X sky130_fd_sc_hd__buf_8
XFILLER_0_91_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout86 _11709_/A vssd1 vssd1 vccd1 vccd1 _09940_/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__10262__A1 _10814_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10262__B2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10531_ _10531_/A _10531_/B vssd1 vssd1 vccd1 vccd1 _10533_/B sky130_fd_sc_hd__xnor2_1
Xfanout97 _11512_/A vssd1 vssd1 vccd1 vccd1 _12094_/A sky130_fd_sc_hd__buf_12
XANTENNA_fanout9_A fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11032__A _12421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08207__A1 _08873_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13250_ _13248_/X _13250_/B vssd1 vssd1 vccd1 vccd1 _13523_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__08207__B2 _08891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10462_ _06986_/Y _12793_/A2 _11586_/B vssd1 vssd1 vccd1 vccd1 _10462_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__13200__A1 _07257_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12201_ _12203_/A _12203_/B _12203_/C vssd1 vssd1 vccd1 vccd1 _12202_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13181_ hold37/X _13191_/B vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__or2_1
X_10393_ _10393_/A _10393_/B vssd1 vssd1 vccd1 vccd1 _10395_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_103_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11762__A1 _11553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12132_ _12131_/A _12131_/B _12131_/Y _10866_/B vssd1 vssd1 vccd1 vccd1 _12132_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12063_ _12046_/A _12709_/A2 _09515_/Y _06869_/B _12062_/Y vssd1 vssd1 vccd1 vccd1
+ _12063_/X sky130_fd_sc_hd__a221o_1
X_11014_ _11014_/A _11014_/B _11014_/C vssd1 vssd1 vccd1 vccd1 _11014_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__06796__A _06928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09172__A _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12965_ reg1_val[25] curr_PC[25] _12978_/S vssd1 vssd1 vccd1 vccd1 _12967_/B sky130_fd_sc_hd__mux2_1
X_11916_ _12016_/B _11916_/B vssd1 vssd1 vccd1 vccd1 _11924_/A sky130_fd_sc_hd__nand2_1
X_12896_ _13054_/B _12897_/B vssd1 vssd1 vccd1 vccd1 _12907_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_68_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11847_ _11847_/A _11847_/B vssd1 vssd1 vccd1 vccd1 _11848_/B sky130_fd_sc_hd__or2_1
XFILLER_0_74_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07249__A2 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ _11776_/Y _11778_/B vssd1 vssd1 vccd1 vccd1 _11779_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_82_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07420__A _10457_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13517_ _13543_/A hold252/X vssd1 vssd1 vccd1 vccd1 _13719_/D sky130_fd_sc_hd__and2_1
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10729_ _12130_/A _11151_/A _11151_/B vssd1 vssd1 vccd1 vccd1 _10729_/X sky130_fd_sc_hd__and3_1
XFILLER_0_125_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13448_ _13463_/B2 _13446_/Y _13447_/X _13450_/B hold245/X vssd1 vssd1 vccd1 vccd1
+ hold246/A sky130_fd_sc_hd__a32o_1
XFILLER_0_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13379_ _13605_/A hold225/X vssd1 vssd1 vccd1 vccd1 _13671_/D sky130_fd_sc_hd__and2_1
Xclkbuf_4_7_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13731_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07940_ _07940_/A _07940_/B _07940_/C vssd1 vssd1 vccd1 vccd1 _07941_/B sky130_fd_sc_hd__and3_1
X_07871_ _07870_/A _07870_/C _07870_/B vssd1 vssd1 vccd1 vccd1 _07872_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__08382__B1 _08580_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09610_ _09610_/A _09610_/B vssd1 vssd1 vccd1 vccd1 _09611_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__08921__A2 _07399_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06822_ reg1_val[28] _09254_/C vssd1 vssd1 vccd1 vccd1 _06824_/B sky130_fd_sc_hd__nand2_1
X_09541_ _13145_/A _11793_/B _09540_/X vssd1 vssd1 vccd1 vccd1 _09541_/X sky130_fd_sc_hd__o21a_1
XANTENNA__11269__B1 _07877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06753_ reg1_val[18] vssd1 vssd1 vccd1 vccd1 _07442_/A sky130_fd_sc_hd__inv_2
XFILLER_0_92_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12466__C1 _12748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11808__A2 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08134__B1 _08778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09472_ _09470_/X _09471_/X _09688_/S vssd1 vssd1 vccd1 vccd1 _09472_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08423_ _08951_/A _08423_/B vssd1 vssd1 vccd1 vccd1 _08485_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10492__A1 _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10492__B2 _12103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout247_A _06886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08354_ _08353_/A _08415_/A vssd1 vssd1 vccd1 vccd1 _08368_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_74_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12233__A2 _12314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07305_ _10095_/A _07305_/B vssd1 vssd1 vccd1 vccd1 _07312_/B sky130_fd_sc_hd__and2_1
XFILLER_0_128_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08285_ _08178_/A _08178_/B _08178_/C vssd1 vssd1 vccd1 vccd1 _08288_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_116_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07236_ _08951_/A _07240_/B vssd1 vssd1 vccd1 vccd1 _07236_/X sky130_fd_sc_hd__and2_1
XANTENNA__11992__B2 _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07660__A2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07167_ _07535_/B _07164_/X _07165_/X vssd1 vssd1 vccd1 vccd1 _08203_/A sky130_fd_sc_hd__o21a_4
XFILLER_0_42_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07098_ _07098_/A _07098_/B _07098_/C _07098_/D vssd1 vssd1 vccd1 vccd1 _07099_/C
+ sky130_fd_sc_hd__or4_1
Xfanout210 _13145_/A vssd1 vssd1 vccd1 vccd1 _09688_/S sky130_fd_sc_hd__clkbuf_8
Xfanout221 _10603_/S vssd1 vssd1 vccd1 vccd1 _10458_/S sky130_fd_sc_hd__clkbuf_8
Xfanout232 _09525_/Y vssd1 vssd1 vccd1 vccd1 _11688_/B sky130_fd_sc_hd__clkbuf_8
Xfanout243 _07108_/D vssd1 vssd1 vccd1 vccd1 _12406_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout254 _13141_/A vssd1 vssd1 vccd1 vccd1 _13599_/D sky130_fd_sc_hd__buf_4
Xfanout265 _13082_/A vssd1 vssd1 vccd1 vccd1 _13136_/A sky130_fd_sc_hd__clkbuf_8
Xfanout276 _13444_/C1 vssd1 vssd1 vccd1 vccd1 _13547_/A sky130_fd_sc_hd__buf_4
Xfanout287 reg1_val[7] vssd1 vssd1 vccd1 vccd1 _13015_/A sky130_fd_sc_hd__buf_6
X_09808_ _09808_/A _09808_/B vssd1 vssd1 vccd1 vccd1 _09821_/A sky130_fd_sc_hd__xor2_4
XANTENNA__13507__A _13543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout298 instruction[4] vssd1 vssd1 vccd1 vccd1 _13748_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout62_A _10518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09739_ _09740_/B _09740_/A vssd1 vssd1 vccd1 vccd1 _09739_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__11027__A _11027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12750_ hold197/A _12750_/B vssd1 vssd1 vccd1 vccd1 _12750_/X sky130_fd_sc_hd__or2_1
XANTENNA__07479__A2 _11047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09873__B1 _11587_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ curr_PC[16] _11794_/C _12825_/S vssd1 vssd1 vccd1 vccd1 _11701_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _12681_/A _12728_/A vssd1 vssd1 vccd1 vccd1 _12682_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_37_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _11743_/B _11632_/B vssd1 vssd1 vccd1 vccd1 _11633_/B sky130_fd_sc_hd__or2_1
XANTENNA__13421__A1 _11913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08336__A _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10235__A1 _10235_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10235__B2 _10235_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11563_ _09048_/B _11562_/X _11866_/A vssd1 vssd1 vccd1 vccd1 _11563_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_64_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11983__A1 _10866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13302_ _13535_/B _13536_/A _13240_/X vssd1 vssd1 vccd1 vccd1 _13540_/B sky130_fd_sc_hd__a21o_1
X_10514_ _10515_/A _10515_/B _10515_/C vssd1 vssd1 vccd1 vccd1 _10516_/A sky130_fd_sc_hd__a21oi_1
X_11494_ _11825_/A _11494_/B vssd1 vssd1 vccd1 vccd1 _11498_/A sky130_fd_sc_hd__xnor2_1
X_13233_ _13233_/A _13233_/B vssd1 vssd1 vccd1 vccd1 _13548_/A sky130_fd_sc_hd__nor2_1
X_10445_ _10445_/A _10445_/B vssd1 vssd1 vccd1 vccd1 _10445_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__07894__B _10787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11196__C1 _11802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13164_ wire122/X _13194_/A2 hold112/X _13539_/A vssd1 vssd1 vccd1 vccd1 _13618_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10376_ fanout34/X _11047_/A _07478_/Y fanout32/X vssd1 vssd1 vccd1 vccd1 _10377_/B
+ sky130_fd_sc_hd__o22a_1
X_12115_ _12203_/A _12115_/B vssd1 vssd1 vccd1 vccd1 _12117_/B sky130_fd_sc_hd__and2_1
X_13095_ _13102_/C _13095_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[22] sky130_fd_sc_hd__xnor2_4
XFILLER_0_20_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12046_ _12046_/A _12046_/B vssd1 vssd1 vccd1 vccd1 _12046_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07167__A1 _07535_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06914__A1 _06936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07415__A _12421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12948_ _12956_/A _12948_/B vssd1 vssd1 vccd1 vccd1 _12949_/B sky130_fd_sc_hd__or2_1
XANTENNA__09864__B1 _12515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10474__A1 _12648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12879_ _12879_/A _12879_/B _12879_/C vssd1 vssd1 vccd1 vccd1 _12880_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_87_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08419__A1 _09671_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08419__B2 _08873_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08246__A _09671_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10226__B2 _07495_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08070_ _08090_/A _08090_/B vssd1 vssd1 vccd1 vccd1 _08070_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07021_ _07025_/B _07025_/C vssd1 vssd1 vccd1 vccd1 _10004_/S sky130_fd_sc_hd__nand2_8
XFILLER_0_70_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08972_ _09023_/A _08971_/A _08971_/B _08883_/X _08882_/X vssd1 vssd1 vccd1 vccd1
+ _08974_/B sky130_fd_sc_hd__a311o_1
X_07923_ _07924_/A _07924_/B vssd1 vssd1 vccd1 vccd1 _09179_/B sky130_fd_sc_hd__or2_1
XANTENNA__09147__A2 _12667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13327__A _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07854_ _07620_/A _07620_/B _07618_/X vssd1 vssd1 vccd1 vccd1 _07873_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10162__B1 _10734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07325__A _11126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06805_ _06804_/Y _06872_/B1 _06873_/B1 reg2_val[30] vssd1 vssd1 vccd1 vccd1 _09254_/A
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_97_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07785_ _07786_/B _07786_/A vssd1 vssd1 vccd1 vccd1 _07785_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_97_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09524_ _09524_/A _09524_/B vssd1 vssd1 vccd1 vccd1 _09524_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11257__A3 _12235_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09455_ reg1_val[13] reg1_val[18] _09463_/S vssd1 vssd1 vccd1 vccd1 _09455_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11662__B1 _11552_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08406_ _08406_/A _08406_/B vssd1 vssd1 vccd1 vccd1 _08472_/B sky130_fd_sc_hd__xnor2_4
X_09386_ _09386_/A _09386_/B vssd1 vssd1 vccd1 vccd1 _09387_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07060__A _13129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08337_ _08340_/A _08340_/B vssd1 vssd1 vccd1 vccd1 _08337_/X sky130_fd_sc_hd__and2_1
XFILLER_0_74_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09428__A_N _13748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09686__S _10007_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08268_ _08821_/B2 fanout76/X fanout74/X _08821_/A1 vssd1 vssd1 vccd1 vccd1 _08269_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_34_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07219_ _08197_/A _09694_/A vssd1 vssd1 vccd1 vccd1 _07219_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08199_ _09949_/A _08199_/B _08199_/C vssd1 vssd1 vccd1 vccd1 _08201_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_104_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10230_ _10374_/B2 fanout9/X fanout4/X _10349_/A1 vssd1 vssd1 vccd1 vccd1 _10231_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07219__B _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10161_ _07015_/Y _09865_/B _07016_/Y _07008_/Y vssd1 vssd1 vccd1 vccd1 _10161_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_30_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10092_ _10093_/A _10093_/B vssd1 vssd1 vccd1 vccd1 _10222_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07235__A _09950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12802_ _12982_/B _12802_/B vssd1 vssd1 vccd1 vccd1 _12803_/B sky130_fd_sc_hd__or2_1
X_10994_ reg1_val[10] curr_PC[10] vssd1 vssd1 vccd1 vccd1 _10999_/A sky130_fd_sc_hd__or2_1
XFILLER_0_69_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12733_ _12733_/A _12733_/B _12733_/C _12635_/Y vssd1 vssd1 vccd1 vccd1 _12733_/X
+ sky130_fd_sc_hd__or4b_2
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06793__B _07398_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _12638_/X _12643_/X _12662_/X _12663_/X vssd1 vssd1 vccd1 vccd1 dest_val[28]
+ sky130_fd_sc_hd__a31oi_4
XANTENNA__08066__A _08951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11615_ _11708_/A _07473_/A fanout7/X _11614_/Y vssd1 vssd1 vccd1 vccd1 _11617_/B
+ sky130_fd_sc_hd__a31o_1
X_12595_ hold273/A _12595_/B vssd1 vssd1 vccd1 vccd1 _12653_/B sky130_fd_sc_hd__or2_1
XFILLER_0_37_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11546_ _11546_/A _11546_/B vssd1 vssd1 vccd1 vccd1 _11549_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_123_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08821__A1 _08821_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08821__B2 _08821_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11477_ hold297/A _11582_/C _11693_/A2 vssd1 vssd1 vccd1 vccd1 _11478_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13216_ hold249/A hold28/X vssd1 vssd1 vccd1 vccd1 _13217_/B sky130_fd_sc_hd__and2b_1
X_10428_ _10428_/A _10428_/B vssd1 vssd1 vccd1 vccd1 _10429_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_21_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08585__B1 _13174_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13147_ _13147_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13147_/Y sky130_fd_sc_hd__nand2_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ _10359_/A _10359_/B vssd1 vssd1 vccd1 vccd1 _10360_/B sky130_fd_sc_hd__xor2_4
XANTENNA__07129__B _07129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13078_ reg1_val[19] _13129_/B vssd1 vssd1 vccd1 vccd1 _13081_/D sky130_fd_sc_hd__xnor2_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13330__B1 _13506_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12029_ _12029_/A _12029_/B _12029_/C vssd1 vssd1 vccd1 vccd1 _12030_/B sky130_fd_sc_hd__or3_1
XANTENNA__13147__A _13147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13581__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07570_ _13015_/A _07320_/C _07320_/D reg1_val[10] vssd1 vssd1 vccd1 vccd1 _07571_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_73_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09240_ _11732_/A fanout79/X fanout70/X fanout83/X vssd1 vssd1 vccd1 vccd1 _09241_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10937__C _11027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09171_ fanout28/X _11047_/A fanout85/X _08395_/B vssd1 vssd1 vccd1 vccd1 _09172_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08122_ _08907_/A _08197_/B _08197_/C vssd1 vssd1 vccd1 vccd1 _08123_/C sky130_fd_sc_hd__or3_1
XFILLER_0_113_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08704__A _09674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08053_ _08053_/A vssd1 vssd1 vccd1 vccd1 _08113_/A sky130_fd_sc_hd__inv_2
XFILLER_0_113_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07004_ reg2_val[3] _07110_/A vssd1 vssd1 vccd1 vccd1 _07004_/X sky130_fd_sc_hd__and2_1
XFILLER_0_3_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11175__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10922__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08955_ _09694_/A _09701_/B _13147_/A _08197_/A vssd1 vssd1 vccd1 vccd1 _09660_/A
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08328__B1 _10814_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06878__B _12981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07906_ _10095_/A _07906_/B vssd1 vssd1 vccd1 vccd1 _07908_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09254__B _09254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08886_ _08882_/X _09023_/A vssd1 vssd1 vccd1 vccd1 _09021_/A sky130_fd_sc_hd__and2b_1
X_07837_ _08027_/A _08027_/B vssd1 vssd1 vccd1 vccd1 _08028_/A sky130_fd_sc_hd__or2_1
XANTENNA__12896__A _13054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07768_ _12421_/A _07768_/B vssd1 vssd1 vccd1 vccd1 _07770_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09270__A _10522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09507_ instruction[3] _13748_/A _09507_/C vssd1 vssd1 vccd1 vccd1 _09507_/X sky130_fd_sc_hd__or3_4
XFILLER_0_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11635__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07699_ _09381_/A _07699_/B vssd1 vssd1 vccd1 vccd1 _07700_/B sky130_fd_sc_hd__nor2_1
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07303__A1 _07572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11305__A _11825_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09438_ _09688_/S _09438_/B vssd1 vssd1 vccd1 vccd1 _09438_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_109_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09369_ _09369_/A _09369_/B vssd1 vssd1 vccd1 vccd1 _09379_/A sky130_fd_sc_hd__xnor2_1
X_11400_ _11400_/A _11400_/B vssd1 vssd1 vccd1 vccd1 _11401_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07606__A2 wire101/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12380_ _12303_/A _12301_/X _06856_/A vssd1 vssd1 vccd1 vccd1 _12380_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_34_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_70 _10751_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_81 reg1_val[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11331_ _11331_/A _11331_/B vssd1 vssd1 vccd1 vccd1 _11332_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09429__B _13748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11262_ _11866_/A _11233_/Y _11238_/X _11261_/X vssd1 vssd1 vccd1 vccd1 _11262_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_30_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13001_ _12999_/Y _13001_/B vssd1 vssd1 vccd1 vccd1 _13002_/B sky130_fd_sc_hd__and2b_1
XANTENNA__11166__A2 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10213_ _10213_/A _10213_/B vssd1 vssd1 vccd1 vccd1 _10215_/B sky130_fd_sc_hd__or2_1
XFILLER_0_120_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11193_ _11193_/A _11193_/B vssd1 vssd1 vccd1 vccd1 _11195_/B sky130_fd_sc_hd__xor2_1
XANTENNA__10374__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ _10144_/A _10144_/B vssd1 vssd1 vccd1 vccd1 _10145_/B sky130_fd_sc_hd__xor2_4
XANTENNA__08319__B1 _07556_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10075_ fanout47/X fanout75/X _08704_/B fanout45/X vssd1 vssd1 vccd1 vccd1 _10076_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12418__A2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10977_ _10977_/A _10977_/B vssd1 vssd1 vccd1 vccd1 _11225_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_69_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12716_ _11823_/A _12668_/B _12671_/B vssd1 vssd1 vccd1 vccd1 _12723_/A sky130_fd_sc_hd__o21ai_2
X_13696_ _13700_/CLK hold72/X vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12647_ _12647_/A _12698_/C vssd1 vssd1 vccd1 vccd1 _12648_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12745__S _12782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12578_ _12578_/A _12578_/B _12578_/C vssd1 vssd1 vccd1 vccd1 _12578_/X sky130_fd_sc_hd__and3_1
XFILLER_0_4_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11529_ _11530_/A _11530_/B vssd1 vssd1 vccd1 vccd1 _11531_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13576__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10904__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09355__A _09575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08740_ _08766_/A _08766_/B vssd1 vssd1 vccd1 vccd1 _08755_/B sky130_fd_sc_hd__or2_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08671_ _08715_/A _08715_/B _08667_/Y vssd1 vssd1 vccd1 vccd1 _08677_/A sky130_fd_sc_hd__o21ai_2
X_07622_ _12421_/A _07622_/B vssd1 vssd1 vccd1 vccd1 _07630_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07553_ _07911_/A _07553_/B vssd1 vssd1 vccd1 vccd1 _07566_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11125__A _11126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07484_ _07486_/C _07486_/D vssd1 vssd1 vccd1 vccd1 _07484_/X sky130_fd_sc_hd__and2_1
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09223_ _09223_/A _09223_/B vssd1 vssd1 vccd1 vccd1 _09225_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09154_ _09154_/A _09154_/B vssd1 vssd1 vccd1 vccd1 _09168_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_44_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08105_ _08997_/A _08997_/B vssd1 vssd1 vccd1 vccd1 _08105_/Y sky130_fd_sc_hd__nand2_1
X_09085_ _09086_/B _09086_/C _09092_/A vssd1 vssd1 vccd1 vccd1 _09087_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_44_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08036_ _08036_/A _08036_/B vssd1 vssd1 vccd1 vccd1 _08037_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10356__B1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09987_ _09650_/A _09650_/B _09824_/A _09824_/B vssd1 vssd1 vccd1 vccd1 _09987_/Y
+ sky130_fd_sc_hd__o22ai_1
X_08938_ _08938_/A _08938_/B _08938_/C vssd1 vssd1 vccd1 vccd1 _08964_/B sky130_fd_sc_hd__and3_1
XANTENNA__10659__A1 _07299_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08869_ _09950_/A _08869_/B vssd1 vssd1 vccd1 vccd1 _08901_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10659__B2 _10814_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10900_ _10900_/A _10900_/B vssd1 vssd1 vccd1 vccd1 _10900_/Y sky130_fd_sc_hd__nand2_1
X_11880_ hold203/A _12311_/B1 _11972_/B _11879_/Y _12533_/B1 vssd1 vssd1 vccd1 vccd1
+ _11889_/C sky130_fd_sc_hd__a311o_1
X_10831_ _10830_/A _10830_/B _10964_/B _10829_/Y vssd1 vssd1 vccd1 vccd1 _10832_/C
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10226__A2_N fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10577__C _10857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13550_ hold255/X _13550_/A2 _13549_/X _13563_/B2 vssd1 vssd1 vccd1 vccd1 hold256/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10762_ curr_PC[6] curr_PC[7] _10480_/B curr_PC[8] vssd1 vssd1 vccd1 vccd1 _10762_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_27_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12501_ _12502_/A _12502_/B _12502_/C vssd1 vssd1 vccd1 vccd1 _12568_/B sky130_fd_sc_hd__o21a_1
X_13481_ hold276/X _13550_/A2 _13480_/X _13563_/B2 vssd1 vssd1 vccd1 vccd1 hold277/A
+ sky130_fd_sc_hd__a22o_1
X_10693_ fanout42/X fanout20/X fanout18/X _12087_/A vssd1 vssd1 vccd1 vccd1 _10694_/B
+ sky130_fd_sc_hd__o22a_1
X_12432_ _12505_/A _12432_/B vssd1 vssd1 vccd1 vccd1 _12435_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12363_ _12363_/A _12363_/B vssd1 vssd1 vccd1 vccd1 _12508_/A sky130_fd_sc_hd__or2_2
XFILLER_0_50_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11314_ _11315_/A _11315_/B _11315_/C vssd1 vssd1 vccd1 vccd1 _11438_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_105_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12294_ _11559_/B _11950_/X _12293_/B _12292_/Y _12293_/X vssd1 vssd1 vccd1 vccd1
+ _12295_/B sky130_fd_sc_hd__a311o_2
XFILLER_0_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11139__A2 _11793_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11245_ _11242_/X _11243_/Y _11125_/X _11129_/B vssd1 vssd1 vccd1 vccd1 _11246_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_120_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08004__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10898__A1 _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11176_ _11913_/A _11176_/B vssd1 vssd1 vccd1 vccd1 _11185_/A sky130_fd_sc_hd__xnor2_1
X_10127_ _10127_/A _10127_/B vssd1 vssd1 vccd1 vccd1 _10128_/B sky130_fd_sc_hd__and2_1
XANTENNA__09903__A _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10058_ _10058_/A _10058_/B vssd1 vssd1 vccd1 vccd1 _10060_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__11600__D_N _11561_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13748_ _13748_/A vssd1 vssd1 vccd1 vccd1 sign_extend sky130_fd_sc_hd__buf_12
XFILLER_0_57_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13679_ _13684_/CLK _13679_/D vssd1 vssd1 vccd1 vccd1 hold161/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10035__C1 _10034_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold104 hold104/A vssd1 vssd1 vccd1 vccd1 hold104/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold115 hold115/A vssd1 vssd1 vccd1 vccd1 hold115/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 hold126/A vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold137 hold137/A vssd1 vssd1 vccd1 vccd1 hold137/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 hold148/A vssd1 vssd1 vccd1 vccd1 hold148/X sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ _09910_/A1 _10518_/A _09754_/B _09752_/Y vssd1 vssd1 vccd1 vccd1 _09912_/B
+ sky130_fd_sc_hd__a31o_1
Xhold159 hold159/A vssd1 vssd1 vccd1 vccd1 hold159/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09841_ _09445_/X _09464_/X _10004_/S vssd1 vssd1 vccd1 vccd1 _09841_/X sky130_fd_sc_hd__mux2_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ _10507_/A _09772_/B vssd1 vssd1 vccd1 vccd1 _09774_/B sky130_fd_sc_hd__xnor2_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06984_ reg1_val[6] _07556_/A vssd1 vssd1 vccd1 vccd1 _10590_/A sky130_fd_sc_hd__nor2_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ _08724_/A _08724_/B _08726_/A _08726_/B vssd1 vssd1 vccd1 vccd1 _08723_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout277_A _13444_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08654_ _08694_/A _08694_/B vssd1 vssd1 vccd1 vccd1 _08982_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_96_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07605_ _10095_/A _07605_/B vssd1 vssd1 vccd1 vccd1 _07671_/A sky130_fd_sc_hd__xnor2_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13054__B _13054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08585_ _08271_/A _13172_/A1 _13174_/A1 _09501_/A vssd1 vssd1 vccd1 vccd1 _08586_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07536_ _07537_/B _07537_/C vssd1 vssd1 vccd1 vccd1 _07536_/X sky130_fd_sc_hd__and2_1
XFILLER_0_76_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07052__B _07230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07467_ _11508_/A _07467_/B vssd1 vssd1 vccd1 vccd1 _07474_/B sky130_fd_sc_hd__or2_1
XFILLER_0_9_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10694__A _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09206_ _09086_/B _09086_/C _09318_/A _09318_/C vssd1 vssd1 vccd1 vccd1 _09206_/X
+ sky130_fd_sc_hd__a211o_1
X_07398_ _11463_/A _07398_/B _09703_/B vssd1 vssd1 vccd1 vccd1 _07400_/B sky130_fd_sc_hd__and3_4
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09137_ _09591_/A _09137_/B vssd1 vssd1 vccd1 vccd1 _09139_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_44_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09431__A1 _12695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09068_ _09068_/A _09068_/B vssd1 vssd1 vccd1 vccd1 _09068_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08019_ _08039_/A _08039_/B vssd1 vssd1 vccd1 vccd1 _08019_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_13_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10329__B1 _10326_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout92_A _11514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11030_ _11209_/B _11030_/B vssd1 vssd1 vccd1 vccd1 _11068_/A sky130_fd_sc_hd__and2_1
X_12981_ instruction[25] _12982_/A _12981_/C vssd1 vssd1 vccd1 vccd1 _12987_/A sky130_fd_sc_hd__and3_4
XFILLER_0_99_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11932_ _11933_/A _11933_/B vssd1 vssd1 vccd1 vccd1 _12014_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10501__B1 _08580_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08339__A _10263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11863_ _11862_/A _12163_/C _11955_/A vssd1 vssd1 vccd1 vccd1 _11863_/X sky130_fd_sc_hd__a21o_1
X_10814_ _10814_/A1 fanout38/X fanout36/X fanout42/X vssd1 vssd1 vccd1 vccd1 _10815_/B
+ sky130_fd_sc_hd__o22a_1
X_13602_ hold15/X _13597_/X _13601_/Y _13605_/A vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__o211a_1
X_11794_ curr_PC[16] curr_PC[17] _11794_/C vssd1 vssd1 vccd1 vccd1 _11893_/B sky130_fd_sc_hd__and3_1
XANTENNA__10804__A1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10745_ _10742_/X _10744_/X _12648_/A vssd1 vssd1 vccd1 vccd1 _10745_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10804__B2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13533_ hold259/X _13555_/A2 _13532_/X _13542_/B2 vssd1 vssd1 vccd1 vccd1 hold260/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13464_ _13547_/A hold265/X vssd1 vssd1 vccd1 vccd1 _13708_/D sky130_fd_sc_hd__and2_1
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10676_ _10676_/A _10676_/B vssd1 vssd1 vccd1 vccd1 _10677_/B sky130_fd_sc_hd__or2_1
XFILLER_0_35_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12415_ _12411_/A _12332_/B _12335_/A vssd1 vssd1 vccd1 vccd1 _12429_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__07028__A3 _12806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13395_ _07274_/B _13207_/B hold162/X vssd1 vssd1 vccd1 vccd1 _13679_/D sky130_fd_sc_hd__a21boi_1
XFILLER_0_23_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12346_ _12346_/A vssd1 vssd1 vccd1 vccd1 _12348_/B sky130_fd_sc_hd__inv_2
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12277_ _12278_/A _12278_/B vssd1 vssd1 vccd1 vccd1 _12358_/B sky130_fd_sc_hd__nand2b_1
X_11228_ _10724_/A _11227_/Y _11226_/X vssd1 vssd1 vccd1 vccd1 _11229_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11159_ _11307_/A _11307_/B vssd1 vssd1 vccd1 vccd1 _11161_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_65_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06976__B _13015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11296__A1 _12557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11296__B2 _12557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07153__A _12578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08370_ _08370_/A _08370_/B vssd1 vssd1 vccd1 vccd1 _08466_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_92_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13442__C1 _13444_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07321_ _11126_/A reg1_val[12] _07328_/B vssd1 vssd1 vccd1 vccd1 _07321_/X sky130_fd_sc_hd__or3_1
XANTENNA__12796__A1 _12796_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11403__A _12092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07252_ _07252_/A _07252_/B _07252_/C _07252_/D vssd1 vssd1 vccd1 vccd1 _07254_/C
+ sky130_fd_sc_hd__or4_2
XANTENNA__12548__A1 _12667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12548__B2 _12614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07183_ _10889_/A _07184_/D vssd1 vssd1 vccd1 vccd1 _07183_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_30_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10023__A2 _10010_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07328__A _11126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12720__A1 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09824_ _09824_/A _09824_/B vssd1 vssd1 vccd1 vccd1 _10433_/A sky130_fd_sc_hd__xnor2_4
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09755_ _09755_/A _09755_/B vssd1 vssd1 vccd1 vccd1 _09788_/A sky130_fd_sc_hd__xnor2_1
X_06967_ reg2_val[8] _06980_/B vssd1 vssd1 vccd1 vccd1 _06967_/X sky130_fd_sc_hd__and2_1
XANTENNA__10689__A _11913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06886__B _12995_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08706_ _08717_/A _08717_/B vssd1 vssd1 vccd1 vccd1 _08719_/A sky130_fd_sc_hd__nand2b_1
X_09686_ _09530_/X _09685_/X _10007_/S vssd1 vssd1 vccd1 vccd1 _09686_/X sky130_fd_sc_hd__mux2_1
X_06898_ _06896_/Y _06906_/B1 _06980_/B reg2_val[17] vssd1 vssd1 vccd1 vccd1 _07300_/A
+ sky130_fd_sc_hd__a2bb2o_2
X_08637_ _08637_/A _08637_/B vssd1 vssd1 vccd1 vccd1 _08686_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ _08566_/X _08567_/X _08515_/X vssd1 vssd1 vccd1 vccd1 _08568_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12236__B1 _09520_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout10 _09146_/Y vssd1 vssd1 vccd1 vccd1 fanout10/X sky130_fd_sc_hd__clkbuf_8
Xfanout21 _07488_/X vssd1 vssd1 vccd1 vccd1 fanout21/X sky130_fd_sc_hd__buf_8
X_07519_ _07517_/A _07517_/B _07517_/C _07517_/D vssd1 vssd1 vccd1 vccd1 _11410_/A
+ sky130_fd_sc_hd__o22ai_2
Xfanout32 _07699_/B vssd1 vssd1 vccd1 vccd1 fanout32/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout43 fanout44/X vssd1 vssd1 vccd1 vccd1 _12557_/B sky130_fd_sc_hd__clkbuf_8
X_08499_ _08521_/B _08521_/A vssd1 vssd1 vccd1 vccd1 _08499_/Y sky130_fd_sc_hd__nand2b_1
Xfanout54 _07204_/Y vssd1 vssd1 vccd1 vccd1 fanout54/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__09652__B2 _09426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout65 _07868_/Y vssd1 vssd1 vccd1 vccd1 _11731_/A sky130_fd_sc_hd__buf_12
XFILLER_0_92_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12409__A _12666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout76 _11423_/A vssd1 vssd1 vccd1 vccd1 fanout76/X sky130_fd_sc_hd__buf_6
XFILLER_0_9_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10530_ _10531_/A _10531_/B vssd1 vssd1 vccd1 vccd1 _10679_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10262__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout87 _07438_/X vssd1 vssd1 vccd1 vccd1 _11709_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout98 _10119_/A vssd1 vssd1 vccd1 vccd1 _12253_/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__12128__B _12164_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10461_ hold237/A _10606_/A2 _10604_/B _12533_/B1 vssd1 vssd1 vccd1 vccd1 _10461_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08207__A2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13200__A2 _13598_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12200_ _12200_/A _12200_/B vssd1 vssd1 vccd1 vccd1 _12203_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_60_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13180_ _13180_/A1 _13194_/A2 hold56/X _13539_/A vssd1 vssd1 vccd1 vccd1 _13626_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10392_ _10392_/A _10392_/B vssd1 vssd1 vccd1 vccd1 _10393_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_60_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12131_ _12131_/A _12131_/B vssd1 vssd1 vccd1 vccd1 _12131_/Y sky130_fd_sc_hd__nor2_1
X_12062_ _06869_/A _09520_/X _12061_/X vssd1 vssd1 vccd1 vccd1 _12062_/Y sky130_fd_sc_hd__o21ai_1
X_11013_ _07093_/B _09509_/X _11010_/Y _11012_/X vssd1 vssd1 vccd1 vccd1 _11014_/C
+ sky130_fd_sc_hd__o211a_1
XANTENNA__06796__B _13042_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12964_ _12964_/A _12964_/B vssd1 vssd1 vccd1 vccd1 new_PC[24] sky130_fd_sc_hd__xor2_4
XFILLER_0_87_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11915_ _11915_/A _11915_/B vssd1 vssd1 vccd1 vccd1 _11916_/B sky130_fd_sc_hd__nand2_1
X_12895_ reg1_val[14] curr_PC[14] _12978_/S vssd1 vssd1 vccd1 vccd1 _12897_/B sky130_fd_sc_hd__mux2_1
X_11846_ _11847_/A _11847_/B vssd1 vssd1 vccd1 vccd1 _11944_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_51_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ reg1_val[17] curr_PC[17] vssd1 vssd1 vccd1 vccd1 _11778_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10789__B1 _11286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10728_ _12130_/A _11151_/B _11151_/A vssd1 vssd1 vccd1 vccd1 _10730_/C sky130_fd_sc_hd__a21o_1
X_13516_ hold251/X _13555_/A2 _13515_/X _13542_/B2 vssd1 vssd1 vccd1 vccd1 hold252/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10659_ _07299_/Y fanout39/X fanout36/X _10814_/A1 vssd1 vssd1 vccd1 vccd1 _10660_/B
+ sky130_fd_sc_hd__o22a_1
X_13447_ hold13/X fanout2/X _13704_/Q vssd1 vssd1 vccd1 vccd1 _13447_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_125_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13378_ hold197/X _13599_/D _13584_/B hold224/X vssd1 vssd1 vccd1 vccd1 hold225/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12329_ _12329_/A fanout7/X vssd1 vssd1 vccd1 vccd1 _12329_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09159__B1 _11823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07148__A _12971_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08906__B1 _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07870_ _07870_/A _07870_/B _07870_/C vssd1 vssd1 vccd1 vccd1 _07872_/A sky130_fd_sc_hd__and3_1
XANTENNA__08382__A1 _08923_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09363__A _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08382__B2 _08866_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06821_ _06824_/A vssd1 vssd1 vccd1 vccd1 _06821_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_92_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09540_ _09432_/X _09433_/X _09539_/X _07152_/X vssd1 vssd1 vccd1 vccd1 _09540_/X
+ sky130_fd_sc_hd__a31o_1
X_06752_ reg1_val[14] vssd1 vssd1 vccd1 vccd1 _06923_/A sky130_fd_sc_hd__inv_2
XANTENNA__11269__B2 _07548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08134__A1 _09173_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08134__B2 _11047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09471_ _11126_/A reg1_val[20] _09493_/S vssd1 vssd1 vccd1 vccd1 _09471_/X sky130_fd_sc_hd__mux2_1
X_08422_ _08866_/B2 fanout82/X fanout76/X _08950_/B vssd1 vssd1 vccd1 vccd1 _08423_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07893__B1 _08328_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10492__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08353_ _08353_/A _08353_/B _08353_/C vssd1 vssd1 vccd1 vccd1 _08415_/A sky130_fd_sc_hd__or3_1
XFILLER_0_58_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13430__A2 _06744_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07304_ _10095_/A _07305_/B vssd1 vssd1 vccd1 vccd1 _10649_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_74_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08284_ _08294_/A _08294_/B vssd1 vssd1 vccd1 vccd1 _08284_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_73_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06999__A2 _06936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07235_ _09950_/A _07235_/B vssd1 vssd1 vccd1 vccd1 _07240_/B sky130_fd_sc_hd__and2_2
XANTENNA__11992__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09398__B1 _10915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13194__A1 _12331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07166_ _07535_/B _07164_/X _07165_/X vssd1 vssd1 vccd1 vccd1 _07166_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_0_41_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07097_ _10736_/A _07097_/B _09701_/A _07091_/Y vssd1 vssd1 vccd1 vccd1 _07098_/D
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout200 _08203_/A vssd1 vssd1 vccd1 vccd1 _09371_/A sky130_fd_sc_hd__buf_12
Xfanout211 _09381_/A vssd1 vssd1 vccd1 vccd1 _13145_/A sky130_fd_sc_hd__buf_4
Xfanout222 _06998_/X vssd1 vssd1 vccd1 vccd1 _10603_/S sky130_fd_sc_hd__clkbuf_4
Xfanout233 _12781_/A vssd1 vssd1 vccd1 vccd1 _11866_/A sky130_fd_sc_hd__buf_4
Xfanout244 _12782_/B vssd1 vssd1 vccd1 vccd1 _12525_/A sky130_fd_sc_hd__buf_4
Xfanout255 hold109/X vssd1 vssd1 vccd1 vccd1 _13141_/A sky130_fd_sc_hd__buf_4
XANTENNA__09273__A _11731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout266 _06894_/B vssd1 vssd1 vccd1 vccd1 _12981_/C sky130_fd_sc_hd__buf_4
X_09807_ _09807_/A _09807_/B vssd1 vssd1 vccd1 vccd1 _09808_/B sky130_fd_sc_hd__nor2_2
Xfanout277 _13444_/C1 vssd1 vssd1 vccd1 vccd1 _13591_/A sky130_fd_sc_hd__buf_2
Xfanout288 reg1_val[30] vssd1 vssd1 vccd1 vccd1 _13129_/A sky130_fd_sc_hd__buf_8
X_07999_ _08486_/B _10522_/A _08868_/B1 fanout24/X vssd1 vssd1 vccd1 vccd1 _08000_/B
+ sky130_fd_sc_hd__o22a_1
X_09738_ _09738_/A _09738_/B vssd1 vssd1 vccd1 vccd1 _09740_/B sky130_fd_sc_hd__xnor2_4
X_09669_ _09665_/X _09668_/X _10600_/S vssd1 vssd1 vccd1 vccd1 _09669_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09873__A1 _09496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ curr_PC[16] _11794_/C vssd1 vssd1 vccd1 vccd1 _11700_/X sky130_fd_sc_hd__or2_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _12680_/A _12680_/B vssd1 vssd1 vccd1 vccd1 _12765_/A sky130_fd_sc_hd__nand2_2
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10866__B _10866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07521__A _07521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _11631_/A _11631_/B vssd1 vssd1 vccd1 vccd1 _11632_/B sky130_fd_sc_hd__and2_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13421__A2 _13445_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11562_ _11562_/A _11562_/B vssd1 vssd1 vccd1 vccd1 _11562_/X sky130_fd_sc_hd__or2_1
XANTENNA__10235__A2 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10513_ _10513_/A _10513_/B vssd1 vssd1 vccd1 vccd1 _10515_/C sky130_fd_sc_hd__xor2_1
X_13301_ _13244_/B _13531_/B _13244_/A vssd1 vssd1 vccd1 vccd1 _13536_/A sky130_fd_sc_hd__o21bai_1
XFILLER_0_24_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11493_ _13180_/A1 fanout8/X fanout3/X _11638_/A vssd1 vssd1 vccd1 vccd1 _11494_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13232_ hold266/X hold48/X vssd1 vssd1 vccd1 vccd1 _13233_/B sky130_fd_sc_hd__and2b_1
X_10444_ _10306_/B _10306_/C _11864_/A vssd1 vssd1 vccd1 vccd1 _10445_/B sky130_fd_sc_hd__o21a_1
XANTENNA__07894__C _10787_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11196__B1 _07477_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08061__B1 _08271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13163_ hold111/X _13191_/B vssd1 vssd1 vccd1 vccd1 hold112/A sky130_fd_sc_hd__or2_1
XFILLER_0_0_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10375_ _10522_/B _10375_/B vssd1 vssd1 vccd1 vccd1 _10379_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10943__B1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12114_ _12114_/A _12114_/B vssd1 vssd1 vccd1 vccd1 _12115_/B sky130_fd_sc_hd__or2_1
X_13094_ _13086_/Y _13090_/B _13088_/B vssd1 vssd1 vccd1 vccd1 _13095_/B sky130_fd_sc_hd__o21ai_4
X_12045_ _07050_/Y _12044_/X _12515_/S vssd1 vssd1 vccd1 vccd1 _12046_/B sky130_fd_sc_hd__mux2_1
XANTENNA__12696__B1 _11866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06914__A2 _13082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12448__B1 _10730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12947_ _12956_/A _12948_/B vssd1 vssd1 vccd1 vccd1 _12947_/X sky130_fd_sc_hd__and2_1
XANTENNA__10474__A2 _09529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12878_ _12879_/A _12879_/B _12879_/C vssd1 vssd1 vccd1 vccd1 _12886_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08419__A2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11829_ _11829_/A _11829_/B vssd1 vssd1 vccd1 vccd1 _11830_/B sky130_fd_sc_hd__xnor2_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08246__B _08246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07020_ _07025_/B _07025_/C vssd1 vssd1 vccd1 vccd1 _07020_/X sky130_fd_sc_hd__and2_1
XANTENNA__13176__A1 _11527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08971_ _08971_/A _08971_/B vssd1 vssd1 vccd1 vccd1 _09021_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_87_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07922_ _09179_/A _07922_/B vssd1 vssd1 vccd1 vccd1 _07924_/B sky130_fd_sc_hd__nand2_1
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09552__B1 _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07853_ _07784_/A _07784_/B _07785_/Y vssd1 vssd1 vccd1 vccd1 _07959_/A sky130_fd_sc_hd__a21bo_2
X_06804_ _06886_/A _13059_/B vssd1 vssd1 vccd1 vccd1 _06804_/Y sky130_fd_sc_hd__nor2_1
X_07784_ _07784_/A _07784_/B vssd1 vssd1 vccd1 vccd1 _07786_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09523_ instruction[3] _09523_/B vssd1 vssd1 vccd1 vccd1 _09523_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_78_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09454_ _09452_/X _09453_/X _09688_/S vssd1 vssd1 vccd1 vccd1 _09454_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10465__A2 _12314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08405_ _08405_/A _08405_/B vssd1 vssd1 vccd1 vccd1 _08472_/A sky130_fd_sc_hd__nand2_2
X_09385_ _09386_/A _09386_/B vssd1 vssd1 vccd1 vccd1 _09385_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_19_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08336_ _09940_/A _08336_/B vssd1 vssd1 vccd1 vccd1 _08340_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11798__A _12163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08267_ _08309_/A _08309_/B vssd1 vssd1 vccd1 vccd1 _08279_/B sky130_fd_sc_hd__and2_1
XFILLER_0_46_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07218_ _12982_/A _12985_/A vssd1 vssd1 vccd1 vccd1 _08271_/A sky130_fd_sc_hd__nor2_8
XFILLER_0_6_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08198_ _07283_/A _07283_/B _08907_/A vssd1 vssd1 vccd1 vccd1 _08199_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_14_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07149_ _13744_/A _09516_/A vssd1 vssd1 vccd1 vccd1 _09520_/B sky130_fd_sc_hd__or2_2
XFILLER_0_30_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09791__B1 _11423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10160_ _11562_/A _10160_/B _10160_/C vssd1 vssd1 vccd1 vccd1 _10160_/X sky130_fd_sc_hd__or3_1
X_10091_ _10091_/A _10091_/B vssd1 vssd1 vccd1 vccd1 _10093_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_100_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12801_ _12982_/B _12802_/B vssd1 vssd1 vccd1 vccd1 _12809_/A sky130_fd_sc_hd__nand2_1
X_10993_ _10992_/A _10992_/B _12047_/C1 vssd1 vssd1 vccd1 vccd1 _10993_/X sky130_fd_sc_hd__o21a_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07857__B1 _09885_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _12765_/B _12732_/B vssd1 vssd1 vccd1 vccd1 _12732_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_38_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _07062_/B _10889_/B _07108_/D vssd1 vssd1 vccd1 vccd1 _12663_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_38_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07609__B1 _10536_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11614_ _07473_/B fanout7/X _11708_/A vssd1 vssd1 vccd1 vccd1 _11614_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12594_ _13668_/Q _12374_/A _12650_/B _12795_/A1 vssd1 vssd1 vccd1 vccd1 _12594_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_52_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11545_ _11546_/A _11546_/B vssd1 vssd1 vccd1 vccd1 _11660_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08821__A2 _08866_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07397__S _12551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13158__A1 _07556_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11501__A _11731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11476_ hold300/A _11476_/B vssd1 vssd1 vccd1 vccd1 _11476_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10427_ _10428_/A _10428_/B vssd1 vssd1 vccd1 vccd1 _10427_/X sky130_fd_sc_hd__and2_1
X_13215_ hold28/X hold249/X vssd1 vssd1 vccd1 vccd1 _13579_/B sky130_fd_sc_hd__and2b_1
XANTENNA__10117__A _10266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08585__A1 _08271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08585__B2 _09501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10358_ _10359_/A _10359_/B vssd1 vssd1 vccd1 vccd1 _10358_/X sky130_fd_sc_hd__and2_1
X_13146_ hold13/X _13193_/B _13145_/Y _13547_/A vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__o211a_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13077_ _13074_/A _13076_/B _13074_/B vssd1 vssd1 vccd1 vccd1 _13079_/A sky130_fd_sc_hd__a21bo_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10289_ _10290_/B _10290_/A vssd1 vssd1 vccd1 vccd1 _10289_/Y sky130_fd_sc_hd__nand2b_1
X_12028_ _12029_/A _12029_/B _12029_/C vssd1 vssd1 vccd1 vccd1 _12120_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__13147__B _13193_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06984__B _07556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09170_ _07864_/A _07863_/B _07861_/X vssd1 vssd1 vccd1 vccd1 _09182_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_8_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08121_ _07198_/A _07198_/B _08197_/A vssd1 vssd1 vccd1 vccd1 _08123_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08273__B1 _09659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08704__B _08704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08052_ _10078_/A _08052_/B vssd1 vssd1 vccd1 vccd1 _08053_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07003_ _07001_/Y _07003_/B vssd1 vssd1 vccd1 vccd1 _10165_/A sky130_fd_sc_hd__and2b_1
XANTENNA__07100__S _13744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout105_A _07276_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08954_ _08954_/A _08954_/B vssd1 vssd1 vccd1 vccd1 _09004_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08328__B2 _08328_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07905_ fanout53/X _10235_/A1 _10235_/B2 fanout47/X vssd1 vssd1 vccd1 vccd1 _07906_/B
+ sky130_fd_sc_hd__o22a_1
X_08885_ _08885_/A _08885_/B vssd1 vssd1 vccd1 vccd1 _09023_/A sky130_fd_sc_hd__or2_1
XANTENNA__07055__B _07201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07836_ _07836_/A _07836_/B vssd1 vssd1 vccd1 vccd1 _08027_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_79_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09551__A _11731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07767_ _09161_/A fanout14/X _07833_/B _09604_/A vssd1 vssd1 vccd1 vccd1 _07768_/B
+ sky130_fd_sc_hd__a22o_1
X_09506_ _13744_/A _09516_/A _09525_/C vssd1 vssd1 vccd1 vccd1 _09506_/X sky130_fd_sc_hd__and3b_4
XANTENNA__11635__A1 wire101/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07698_ _10119_/A _07698_/B vssd1 vssd1 vccd1 vccd1 _07704_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11635__B2 _13180_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09437_ _08197_/A _13135_/A _09463_/S vssd1 vssd1 vccd1 vccd1 _09438_/B sky130_fd_sc_hd__mux2_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09368_ _09368_/A _09368_/B vssd1 vssd1 vccd1 vccd1 _09369_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_35_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout18_A _07493_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08319_ _07492_/Y _07545_/Y _07556_/Y _07541_/X vssd1 vssd1 vccd1 vccd1 _08320_/B
+ sky130_fd_sc_hd__a22o_1
X_09299_ _09299_/A _09299_/B vssd1 vssd1 vccd1 vccd1 _09304_/A sky130_fd_sc_hd__or2_4
XANTENNA_60 reg2_val[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12417__A _12417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_71 _11774_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_82 reg1_val[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11330_ _11331_/A _11331_/B vssd1 vssd1 vccd1 vccd1 _11330_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_6_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11261_ _12537_/B2 _11241_/X _11247_/X _12760_/A1 _11260_/X vssd1 vssd1 vccd1 vccd1
+ _11261_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_120_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13000_ reg1_val[4] _13000_/B vssd1 vssd1 vccd1 vccd1 _13001_/B sky130_fd_sc_hd__nand2_1
X_10212_ _10212_/A _10212_/B vssd1 vssd1 vccd1 vccd1 _10213_/B sky130_fd_sc_hd__nor2_1
X_11192_ _11193_/A _11193_/B vssd1 vssd1 vccd1 vccd1 _11326_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10374__A1 _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10374__B2 _10374_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10143_ _10144_/A _10144_/B vssd1 vssd1 vccd1 vccd1 _10143_/X sky130_fd_sc_hd__and2_1
XANTENNA__08319__A1 _07492_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08319__B2 _07541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10074_ _10074_/A vssd1 vssd1 vccd1 vccd1 _10082_/A sky130_fd_sc_hd__inv_2
Xmax_cap73 _07544_/Y vssd1 vssd1 vccd1 vccd1 _11527_/A sky130_fd_sc_hd__buf_6
XFILLER_0_69_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ _10976_/A _10976_/B _10976_/C vssd1 vssd1 vccd1 vccd1 _10977_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_84_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12715_ _09254_/B _12799_/A2 _12690_/Y _12714_/X _12971_/S vssd1 vssd1 vccd1 vccd1
+ dest_val[29] sky130_fd_sc_hd__o221a_4
X_13695_ _13700_/CLK hold148/X vssd1 vssd1 vccd1 vccd1 hold146/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12646_ _12589_/A _12586_/Y _12588_/B vssd1 vssd1 vccd1 vccd1 _12698_/C sky130_fd_sc_hd__o21ai_2
XFILLER_0_26_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12327__A _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12577_ _12635_/C _12575_/X _12576_/Y vssd1 vssd1 vccd1 vccd1 _12577_/X sky130_fd_sc_hd__o21a_1
XANTENNA__11231__A _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11528_ _11528_/A _11528_/B vssd1 vssd1 vccd1 vccd1 _11530_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11459_ _11458_/A _11458_/B _11955_/A vssd1 vssd1 vccd1 vccd1 _11459_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08540__A _10236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ _13129_/A _13129_/B vssd1 vssd1 vccd1 vccd1 _13131_/A sky130_fd_sc_hd__or2_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08670_ _08670_/A _08670_/B vssd1 vssd1 vccd1 vccd1 _08715_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09371__A _09371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07621_ fanout14/X _09955_/A _07833_/B _10104_/A vssd1 vssd1 vccd1 vccd1 _07622_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07552_ _07552_/A _07552_/B vssd1 vssd1 vccd1 vccd1 _07553_/B sky130_fd_sc_hd__or2_1
XFILLER_0_76_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07483_ _07483_/A _07637_/B vssd1 vssd1 vccd1 vccd1 _07486_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_29_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09222_ _09119_/A _09119_/B _09120_/Y vssd1 vssd1 vccd1 vccd1 _09223_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_33_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09153_ _09153_/A _09153_/B vssd1 vssd1 vccd1 vccd1 _09154_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_56_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10456__S _10456_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08104_ _08104_/A _08104_/B vssd1 vssd1 vccd1 vccd1 _08997_/B sky130_fd_sc_hd__xor2_4
X_09084_ _09080_/A _09080_/B _09080_/C _09081_/A _09003_/A vssd1 vssd1 vccd1 vccd1
+ _09086_/C sky130_fd_sc_hd__a311o_2
XFILLER_0_71_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08035_ _08999_/A _08999_/B vssd1 vssd1 vccd1 vccd1 _08035_/X sky130_fd_sc_hd__and2_1
XFILLER_0_114_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13542__B2 _13542_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10356__A1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10356__B2 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09986_ _09986_/A _10150_/A _10298_/A _10433_/A vssd1 vssd1 vccd1 vccd1 _10579_/B
+ sky130_fd_sc_hd__or4_1
X_08937_ _08938_/A _08938_/C _08938_/B vssd1 vssd1 vccd1 vccd1 _08937_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_99_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10659__A2 fanout39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08868_ _08907_/A _09216_/B2 _08868_/B1 _08197_/A vssd1 vssd1 vccd1 vccd1 _08869_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_99_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07819_ _07819_/A _07819_/B vssd1 vssd1 vccd1 vccd1 _07830_/B sky130_fd_sc_hd__and2_1
X_08799_ _08799_/A _08799_/B vssd1 vssd1 vccd1 vccd1 _08820_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10830_ _10830_/A _10830_/B _10964_/B _10829_/Y vssd1 vssd1 vccd1 vccd1 _10832_/B
+ sky130_fd_sc_hd__or4bb_1
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10577__D _10981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10761_ _11866_/A _10731_/X _10732_/Y _10760_/X _10730_/X vssd1 vssd1 vccd1 vccd1
+ _10761_/X sky130_fd_sc_hd__a311o_1
XANTENNA__12846__S _12867_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12500_ _12568_/A _12500_/B vssd1 vssd1 vccd1 vccd1 _12502_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_82_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10692_ _11709_/A _10692_/B vssd1 vssd1 vccd1 vccd1 _10696_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13480_ hold287/A _13479_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13480_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08625__A _10236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12431_ _12431_/A _12431_/B vssd1 vssd1 vccd1 vccd1 _12432_/B sky130_fd_sc_hd__or2_1
XFILLER_0_81_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12362_ _12362_/A _12362_/B _12362_/C vssd1 vssd1 vccd1 vccd1 _12363_/B sky130_fd_sc_hd__and3_1
XFILLER_0_90_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11313_ _11174_/A _11173_/Y _11172_/A vssd1 vssd1 vccd1 vccd1 _11318_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12293_ _11949_/Y _12293_/B vssd1 vssd1 vccd1 vccd1 _12293_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_50_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11244_ _11125_/X _11129_/B _11242_/X _11243_/Y vssd1 vssd1 vccd1 vccd1 _11244_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13533__B2 _13542_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11175_ fanout50/X fanout29/X fanout27/X fanout51/X vssd1 vssd1 vccd1 vccd1 _11176_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10126_ _10127_/A _10127_/B vssd1 vssd1 vccd1 vccd1 _10128_/A sky130_fd_sc_hd__nor2_1
X_10057_ _10057_/A _10057_/B vssd1 vssd1 vccd1 vccd1 _10058_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12610__A _12666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09268__A2 _12764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08476__B1 _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13747_ instruction[10] vssd1 vssd1 vccd1 vccd1 pred_idx[2] sky130_fd_sc_hd__buf_12
XFILLER_0_70_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10959_ _10959_/A _10959_/B vssd1 vssd1 vccd1 vccd1 _10972_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_58_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13678_ _13684_/CLK hold100/X vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12629_ _12508_/X _12629_/B vssd1 vssd1 vccd1 vccd1 _12629_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_72_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08779__A1 _09671_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11896__A _12372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold105 hold105/A vssd1 vssd1 vccd1 vccd1 hold105/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold116 hold116/A vssd1 vssd1 vccd1 vccd1 hold116/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold127 hold127/A vssd1 vssd1 vccd1 vccd1 hold127/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 hold138/A vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 hold149/A vssd1 vssd1 vccd1 vccd1 hold149/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10338__A1 _12047_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10338__B2 _12759_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09840_ _09442_/X _09448_/X _10004_/S vssd1 vssd1 vccd1 vccd1 _09840_/X sky130_fd_sc_hd__mux2_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ fanout56/X fanout75/X _08704_/B fanout53/X vssd1 vssd1 vccd1 vccd1 _09772_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_95_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06983_ reg1_val[6] _07557_/A vssd1 vssd1 vccd1 vccd1 _10588_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_95_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08722_ _08722_/A _08722_/B vssd1 vssd1 vccd1 vccd1 _08726_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_28_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07614__A _10095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09900__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08653_ _08653_/A _08653_/B vssd1 vssd1 vccd1 vccd1 _08694_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07604_ fanout56/X _10235_/B2 fanout40/X _10235_/A1 vssd1 vssd1 vccd1 vccd1 _07605_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08584_ _09373_/A _08584_/B vssd1 vssd1 vccd1 vccd1 _08588_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12799__C1 _12971_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07535_ _07535_/A _07535_/B vssd1 vssd1 vccd1 vccd1 _07537_/C sky130_fd_sc_hd__nand2_2
XFILLER_0_48_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07466_ _11508_/A _07467_/B vssd1 vssd1 vccd1 vccd1 _07473_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_36_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09205_ _09318_/A _09318_/C vssd1 vssd1 vccd1 vccd1 _09205_/X sky130_fd_sc_hd__or2_1
XFILLER_0_107_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13070__B _13129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07397_ _12485_/A _07401_/B _12551_/A vssd1 vssd1 vccd1 vccd1 _07397_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09136_ fanout83/X fanout74/X fanout70/X fanout79/X vssd1 vssd1 vccd1 vccd1 _09137_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09067_ _09062_/A _09062_/B _09065_/X _11957_/C _11957_/B vssd1 vssd1 vccd1 vccd1
+ _12213_/B sky130_fd_sc_hd__o2111ai_2
XFILLER_0_71_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09719__B1 _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12318__A2 _09520_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08018_ _08018_/A _08018_/B vssd1 vssd1 vccd1 vccd1 _08039_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_8_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10329__B2 _10327_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13687__CLK _13701_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout85_A _07478_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ _09808_/A _09808_/B _09807_/A vssd1 vssd1 vccd1 vccd1 _09979_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_99_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12980_ _12980_/A _12980_/B vssd1 vssd1 vccd1 vccd1 new_PC[27] sky130_fd_sc_hd__xnor2_4
XFILLER_0_99_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11931_ _11931_/A _11931_/B vssd1 vssd1 vccd1 vccd1 _11933_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10501__A1 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10501__B2 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11046__A _11823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11862_ _11862_/A _12163_/C vssd1 vssd1 vccd1 vccd1 _11862_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13601_ _13207_/B _13597_/X hold15/X vssd1 vssd1 vccd1 vccd1 _13601_/Y sky130_fd_sc_hd__o21ai_1
X_10813_ _10813_/A _10813_/B vssd1 vssd1 vccd1 vccd1 _10827_/A sky130_fd_sc_hd__xnor2_1
X_11793_ _11793_/A _11793_/B vssd1 vssd1 vccd1 vccd1 _11793_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10265__B1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13532_ hold257/X _13531_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13532_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_54_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10744_ _10595_/Y _10743_/X _11576_/A vssd1 vssd1 vccd1 vccd1 _10744_/X sky130_fd_sc_hd__mux2_2
XANTENNA__10804__A2 _11423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13463_ hold264/X _13450_/B _13462_/X _13463_/B2 vssd1 vssd1 vccd1 vccd1 hold265/A
+ sky130_fd_sc_hd__a22o_1
X_10675_ _10676_/A _10676_/B vssd1 vssd1 vccd1 vccd1 _10811_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12414_ _12414_/A _12414_/B vssd1 vssd1 vccd1 vccd1 _12431_/A sky130_fd_sc_hd__xor2_1
X_13394_ hold98/X _13416_/A2 _13420_/B1 hold161/X _13383_/A vssd1 vssd1 vccd1 vccd1
+ hold162/A sky130_fd_sc_hd__o221a_1
XFILLER_0_23_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12345_ _12426_/A _12345_/B vssd1 vssd1 vccd1 vccd1 _12346_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08630__B1 _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13506__B2 _13506_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12276_ _12276_/A _12276_/B vssd1 vssd1 vccd1 vccd1 _12278_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11517__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11227_ _11227_/A _11454_/A vssd1 vssd1 vccd1 vccd1 _11227_/Y sky130_fd_sc_hd__nand2_1
X_11158_ _07538_/X fanout6/X _11157_/Y _10507_/A vssd1 vssd1 vccd1 vccd1 _11307_/B
+ sky130_fd_sc_hd__a22o_2
X_10109_ _10109_/A _10109_/B vssd1 vssd1 vccd1 vccd1 _10110_/B sky130_fd_sc_hd__xor2_4
X_11089_ _10939_/A _10939_/B _10938_/A vssd1 vssd1 vccd1 vccd1 _11091_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__12340__A _12666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13155__B _13191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11296__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12994__B _12995_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13442__B1 _13444_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07320_ _13015_/A reg1_val[10] _07320_/C _07320_/D vssd1 vssd1 vccd1 vccd1 _07328_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_0_85_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07251_ _07251_/A _07594_/B vssd1 vssd1 vccd1 vccd1 _07251_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12548__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07182_ _07186_/B _07186_/C vssd1 vssd1 vccd1 vccd1 _07193_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_26_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09823_ _09824_/A _09824_/B vssd1 vssd1 vccd1 vccd1 _09823_/X sky130_fd_sc_hd__or2_1
XANTENNA__09824__A _09824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12720__A2 _12666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09754_ _09752_/Y _09754_/B vssd1 vssd1 vccd1 vccd1 _09755_/B sky130_fd_sc_hd__and2b_1
X_06966_ _06963_/Y _06966_/B vssd1 vssd1 vccd1 vccd1 _10870_/A sky130_fd_sc_hd__nand2b_1
X_08705_ _11072_/A _08742_/A _08742_/B vssd1 vssd1 vccd1 vccd1 _08717_/B sky130_fd_sc_hd__mux2_1
X_09685_ _09483_/X _09485_/X _13145_/A vssd1 vssd1 vccd1 vccd1 _09685_/X sky130_fd_sc_hd__mux2_1
X_06897_ reg2_val[17] _06980_/B _06906_/B1 _06896_/Y vssd1 vssd1 vccd1 vccd1 _11793_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_96_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08636_ _08951_/A _08636_/B vssd1 vssd1 vccd1 vccd1 _08686_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_68_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08567_ _08569_/A _08569_/B vssd1 vssd1 vccd1 vccd1 _08567_/X sky130_fd_sc_hd__or2_1
Xfanout22 fanout23/X vssd1 vssd1 vccd1 vccd1 _08486_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__10247__B1 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07518_ _11281_/A _07524_/A vssd1 vssd1 vccd1 vccd1 _07518_/Y sky130_fd_sc_hd__nor2_1
Xfanout33 _07401_/Y vssd1 vssd1 vccd1 vccd1 _07699_/B sky130_fd_sc_hd__buf_6
XFILLER_0_119_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout44 _07256_/Y vssd1 vssd1 vccd1 vccd1 fanout44/X sky130_fd_sc_hd__buf_4
X_08498_ _08498_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _08521_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout66 _08778_/B vssd1 vssd1 vccd1 vccd1 fanout66/X sky130_fd_sc_hd__buf_6
Xfanout77 _07527_/Y vssd1 vssd1 vccd1 vccd1 _11423_/A sky130_fd_sc_hd__clkbuf_8
X_07449_ _07449_/A _07476_/B vssd1 vssd1 vccd1 vccd1 _07449_/Y sky130_fd_sc_hd__nor2_1
Xfanout88 _11507_/A vssd1 vssd1 vccd1 vccd1 _10263_/A sky130_fd_sc_hd__buf_12
XFILLER_0_9_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout99 _11603_/A vssd1 vssd1 vccd1 vccd1 _10119_/A sky130_fd_sc_hd__buf_12
XFILLER_0_107_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10460_ _10606_/A2 _10604_/B hold237/A vssd1 vssd1 vccd1 vccd1 _10460_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09119_ _09119_/A _09119_/B vssd1 vssd1 vccd1 vccd1 _09121_/B sky130_fd_sc_hd__xnor2_1
X_10391_ _10391_/A _10391_/B vssd1 vssd1 vccd1 vccd1 _10393_/A sky130_fd_sc_hd__nand2_1
X_12130_ _12130_/A _12130_/B vssd1 vssd1 vccd1 vccd1 _12131_/B sky130_fd_sc_hd__and2_1
XFILLER_0_60_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12061_ _07201_/A _12799_/A2 _11688_/B reg1_val[20] vssd1 vssd1 vccd1 vccd1 _12061_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09707__A3 _12314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11012_ _06958_/B _11587_/A2 _09520_/X _06956_/Y _11011_/X vssd1 vssd1 vccd1 vccd1
+ _11012_/X sky130_fd_sc_hd__o221a_1
XANTENNA__12711__A2 _12754_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12963_ _12963_/A _12963_/B _12963_/C _12963_/D vssd1 vssd1 vccd1 vccd1 _12964_/B
+ sky130_fd_sc_hd__and4_2
XFILLER_0_99_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11914_ _11915_/A _11915_/B vssd1 vssd1 vccd1 vccd1 _12016_/B sky130_fd_sc_hd__or2_1
XFILLER_0_87_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12894_ _12900_/B _12894_/B vssd1 vssd1 vccd1 vccd1 new_PC[13] sky130_fd_sc_hd__and2_4
X_11845_ _11845_/A _11845_/B vssd1 vssd1 vccd1 vccd1 _11847_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13424__B1 _13444_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ reg1_val[17] curr_PC[17] vssd1 vssd1 vccd1 vccd1 _11776_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_82_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13515_ hold289/A _13514_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13515_/X sky130_fd_sc_hd__mux2_1
X_10727_ _10727_/A _10727_/B _10727_/C _10727_/D vssd1 vssd1 vccd1 vccd1 _11151_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_0_43_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13446_ _13704_/Q hold13/X fanout2/X vssd1 vssd1 vccd1 vccd1 _13446_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_125_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10658_ _12421_/A _10658_/B vssd1 vssd1 vccd1 vccd1 _10666_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13377_ _13605_/A hold198/X vssd1 vssd1 vccd1 vccd1 hold199/A sky130_fd_sc_hd__and2_1
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10589_ _10589_/A _10589_/B vssd1 vssd1 vccd1 vccd1 _10590_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_51_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12328_ _12406_/B1 _12324_/X _12327_/X vssd1 vssd1 vccd1 vccd1 dest_val[23] sky130_fd_sc_hd__o21ai_4
XFILLER_0_11_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09159__A1 _13129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06989__C_N _13010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12259_ _12336_/A _12259_/B vssd1 vssd1 vccd1 vccd1 _12260_/C sky130_fd_sc_hd__and2_1
XANTENNA__12989__B _12990_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11910__B1 _07891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08382__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06820_ _12647_/A _07062_/B vssd1 vssd1 vccd1 vccd1 _06824_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_92_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06751_ reg1_val[12] vssd1 vssd1 vccd1 vccd1 _07535_/A sky130_fd_sc_hd__inv_2
XANTENNA__08134__A2 _10538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09470_ reg1_val[10] reg1_val[21] _09493_/S vssd1 vssd1 vccd1 vccd1 _09470_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_92_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08421_ _08427_/A _08427_/B vssd1 vssd1 vccd1 vccd1 _08421_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_25_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08352_ _08349_/A _08349_/C _08349_/B vssd1 vssd1 vccd1 vccd1 _08353_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11977__B1 _12793_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07303_ _07572_/S _10750_/A _10750_/B _07301_/X vssd1 vssd1 vccd1 vccd1 _07305_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08283_ _08345_/A _08345_/B _08262_/X vssd1 vssd1 vccd1 vccd1 _08294_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07330__C _07435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout135_A _12056_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07234_ _09950_/A _07235_/B vssd1 vssd1 vccd1 vccd1 _07240_/A sky130_fd_sc_hd__nor2_4
XANTENNA__06999__A3 _13005_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09398__A1 fanout39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09398__B2 _08118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07165_ reg1_val[3] _07572_/S vssd1 vssd1 vccd1 vccd1 _07165_/X sky130_fd_sc_hd__or2_2
XANTENNA__13194__A2 _13194_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07096_ _10449_/A _10311_/A _10165_/A _10026_/A vssd1 vssd1 vccd1 vccd1 _07098_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_0_41_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout201 _07166_/Y vssd1 vssd1 vccd1 vccd1 _08951_/A sky130_fd_sc_hd__buf_12
XFILLER_0_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout212 _07028_/Y vssd1 vssd1 vccd1 vccd1 _09381_/A sky130_fd_sc_hd__buf_4
Xfanout223 _06989_/X vssd1 vssd1 vccd1 vccd1 _12648_/A sky130_fd_sc_hd__buf_4
Xfanout234 _09506_/X vssd1 vssd1 vccd1 vccd1 _12047_/C1 sky130_fd_sc_hd__clkbuf_8
Xfanout245 _06988_/X vssd1 vssd1 vccd1 vccd1 _12782_/B sky130_fd_sc_hd__buf_4
Xfanout256 _12754_/C vssd1 vssd1 vccd1 vccd1 _12235_/C sky130_fd_sc_hd__buf_4
XFILLER_0_5_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09806_ _09806_/A _09806_/B vssd1 vssd1 vccd1 vccd1 _09807_/B sky130_fd_sc_hd__nor2_1
Xfanout267 _06920_/B vssd1 vssd1 vccd1 vccd1 _06980_/B sky130_fd_sc_hd__clkbuf_8
Xfanout278 _13430_/C1 vssd1 vssd1 vccd1 vccd1 _13383_/A sky130_fd_sc_hd__buf_4
X_07998_ _08093_/A _08093_/B _07995_/X vssd1 vssd1 vccd1 vccd1 _08018_/B sky130_fd_sc_hd__o21ai_2
Xfanout289 reg1_val[1] vssd1 vssd1 vccd1 vccd1 _09694_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__07581__B1 _07544_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09737_ _09568_/A _09568_/B _09566_/Y vssd1 vssd1 vccd1 vccd1 _09738_/B sky130_fd_sc_hd__a21oi_4
X_06949_ _11126_/A _07472_/A vssd1 vssd1 vccd1 vccd1 _06950_/B sky130_fd_sc_hd__nand2_1
X_09668_ _09666_/X _09667_/X _10005_/S vssd1 vssd1 vccd1 vccd1 _09668_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09873__A2 _11793_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07802__A _10078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08619_ _08980_/A _08980_/B vssd1 vssd1 vccd1 vccd1 _08981_/B sky130_fd_sc_hd__nand2_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ _09599_/A _09599_/B vssd1 vssd1 vccd1 vccd1 _09600_/C sky130_fd_sc_hd__xnor2_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _11631_/A _11631_/B vssd1 vssd1 vccd1 vccd1 _11743_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_126_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11561_ _11561_/A _11561_/B vssd1 vssd1 vccd1 vccd1 _11561_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_80_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13300_ _13527_/A _13527_/B _13247_/A vssd1 vssd1 vccd1 vccd1 _13531_/B sky130_fd_sc_hd__a21oi_1
X_10512_ _10380_/A _10380_/B _10378_/X vssd1 vssd1 vccd1 vccd1 _10513_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08633__A _09659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11492_ _11348_/B _11600_/B _11457_/Y _11864_/A vssd1 vssd1 vccd1 vccd1 _11561_/A
+ sky130_fd_sc_hd__o31ai_1
XFILLER_0_80_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13231_ hold48/X hold266/X vssd1 vssd1 vccd1 vccd1 _13233_/A sky130_fd_sc_hd__and2b_1
X_10443_ _12130_/A _10344_/X _10441_/X _11955_/A vssd1 vssd1 vccd1 vccd1 _10443_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_0_33_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08061__A1 _12982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13162_ _07494_/X _13194_/A2 hold69/X _13547_/A vssd1 vssd1 vccd1 vccd1 _13617_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08061__B2 _07198_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10374_ _10637_/A fanout9/X fanout4/X _10374_/B2 vssd1 vssd1 vccd1 vccd1 _10375_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10943__A1 _12557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10943__B2 _07597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12113_ _12114_/A _12114_/B vssd1 vssd1 vccd1 vccd1 _12203_/A sky130_fd_sc_hd__nand2_1
X_13093_ _13093_/A _13093_/B vssd1 vssd1 vccd1 vccd1 _13102_/C sky130_fd_sc_hd__nand2_2
XFILLER_0_20_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12044_ _11961_/A _11959_/X _06884_/B vssd1 vssd1 vccd1 vccd1 _12044_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10403__A _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06914__A3 _06928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12946_ reg1_val[22] curr_PC[22] _12978_/S vssd1 vssd1 vccd1 vccd1 _12948_/B sky130_fd_sc_hd__mux2_1
X_12877_ _12886_/A _12877_/B vssd1 vssd1 vccd1 vccd1 _12879_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11828_ _11829_/A _11829_/B vssd1 vssd1 vccd1 vccd1 _11828_/Y sky130_fd_sc_hd__nand2_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07150__C _12578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11759_ _11757_/Y _11759_/B vssd1 vssd1 vccd1 vccd1 _11948_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_71_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08543__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13429_ _12253_/A _13598_/C hold71/X vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__o21a_1
XANTENNA__13176__A2 _13194_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08970_ _08970_/A _08970_/B vssd1 vssd1 vccd1 vccd1 _09019_/B sky130_fd_sc_hd__xor2_1
X_07921_ _07921_/A _07921_/B vssd1 vssd1 vccd1 vccd1 _07922_/B sky130_fd_sc_hd__or2_1
XANTENNA__09552__A1 _07833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11409__A _11709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09552__B2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07852_ _07963_/A _07963_/B _07787_/X vssd1 vssd1 vccd1 vccd1 _07962_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06803_ instruction[40] _12981_/C vssd1 vssd1 vccd1 vccd1 _13059_/B sky130_fd_sc_hd__and2_4
X_07783_ _07783_/A _07783_/B vssd1 vssd1 vccd1 vccd1 _07784_/B sky130_fd_sc_hd__xor2_1
X_09522_ instruction[3] _09524_/B vssd1 vssd1 vccd1 vccd1 _09522_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07622__A _12421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09453_ reg1_val[14] reg1_val[17] _09463_/S vssd1 vssd1 vccd1 vccd1 _09453_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11662__A2 _11550_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout252_A _13141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08404_ _08403_/A _08403_/B _08403_/C vssd1 vssd1 vccd1 vccd1 _08405_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09384_ _10522_/B _09384_/B vssd1 vssd1 vccd1 vccd1 _09386_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08335_ _13149_/A fanout24/X _08486_/B _08923_/B1 vssd1 vssd1 vccd1 vccd1 _08336_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09549__A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08266_ _10236_/A _08266_/B vssd1 vssd1 vccd1 vccd1 _08309_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11798__B _12163_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07217_ _07217_/A _07217_/B vssd1 vssd1 vccd1 vccd1 _07217_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08197_ _08197_/A _08197_/B _08197_/C vssd1 vssd1 vccd1 vccd1 _08199_/B sky130_fd_sc_hd__or3_1
XFILLER_0_116_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07148_ _12971_/S _07148_/B vssd1 vssd1 vccd1 vccd1 dest_mask[1] sky130_fd_sc_hd__nand2_8
XANTENNA__09240__B1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09791__A1 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09791__B2 _08246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07079_ _07079_/A _07079_/B vssd1 vssd1 vccd1 vccd1 _07079_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09284__A _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10090_ _10091_/A _10091_/B vssd1 vssd1 vccd1 vccd1 _10222_/A sky130_fd_sc_hd__and2_1
XFILLER_0_100_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09543__A1 _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07554__B1 _07471_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12800_ _09501_/A curr_PC[0] _12867_/S vssd1 vssd1 vccd1 vccd1 _12802_/B sky130_fd_sc_hd__mux2_1
X_10992_ _10992_/A _10992_/B vssd1 vssd1 vccd1 vccd1 _10992_/Y sky130_fd_sc_hd__nand2_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12731_ _12731_/A _12731_/B _12731_/C vssd1 vssd1 vccd1 vccd1 _12732_/B sky130_fd_sc_hd__or3_1
XANTENNA__07857__A1 _10049_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07857__B2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10861__B1 _10900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07251__B _07594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12662_ _10866_/B _12644_/X _12645_/Y _12661_/X vssd1 vssd1 vccd1 vccd1 _12662_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07609__A1 _11922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _11913_/A _11613_/B vssd1 vssd1 vccd1 vccd1 _11617_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08806__B1 _08806_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07609__B2 _11997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12602__A1 _09839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12593_ _12374_/A _12650_/B _13668_/Q vssd1 vssd1 vccd1 vccd1 _12593_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11544_ _11544_/A _11544_/B vssd1 vssd1 vccd1 vccd1 _11546_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13158__A2 _13196_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11475_ hold289/A _11579_/C _12058_/A vssd1 vssd1 vccd1 vccd1 _11476_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__08082__B _08088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13214_ _13313_/A _13214_/B vssd1 vssd1 vccd1 vccd1 _13579_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_122_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10426_ _10426_/A _10426_/B vssd1 vssd1 vccd1 vccd1 _10428_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09231__B1 _10536_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08585__A2 _13172_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09782__A1 _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13145_ _13145_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13145_/Y sky130_fd_sc_hd__nand2_1
X_10357_ _11281_/A _10357_/B vssd1 vssd1 vccd1 vccd1 _10359_/B sky130_fd_sc_hd__xnor2_2
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_max_cap148_A _07420_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _13081_/C _13076_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[18] sky130_fd_sc_hd__xnor2_4
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10288_ _10288_/A _10288_/B vssd1 vssd1 vccd1 vccd1 _10290_/B sky130_fd_sc_hd__xnor2_2
X_12027_ _12027_/A _12027_/B vssd1 vssd1 vccd1 vccd1 _12029_/C sky130_fd_sc_hd__xor2_1
XANTENNA__13330__A2 _13506_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11229__A _11452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08538__A _08746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10787__B _10787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12929_ _12956_/A _12929_/B vssd1 vssd1 vccd1 vccd1 _12930_/B sky130_fd_sc_hd__or2_1
XANTENNA__13163__B _13191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07161__B _07572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11899__A _12417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09429__D_N _13744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08120_ _10239_/A _08120_/B vssd1 vssd1 vccd1 vccd1 _08125_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08273__A1 _08272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08051_ _07307_/Y fanout82/X fanout76/X _08833_/B vssd1 vssd1 vccd1 vccd1 _08052_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07002_ reg1_val[4] _10603_/S vssd1 vssd1 vccd1 vccd1 _07003_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_24_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07379__A3 _07634_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08953_ _08954_/A _08953_/B vssd1 vssd1 vccd1 vccd1 _08953_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__08328__A2 _11732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07904_ _09575_/A _07904_/B vssd1 vssd1 vccd1 vccd1 _07908_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08884_ _08861_/A _08861_/B _08861_/C vssd1 vssd1 vccd1 vccd1 _08973_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07835_ _07835_/A vssd1 vssd1 vccd1 vccd1 _08027_/A sky130_fd_sc_hd__inv_2
XFILLER_0_79_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07766_ _07970_/A _07970_/B _07766_/C vssd1 vssd1 vccd1 vccd1 _07770_/A sky130_fd_sc_hd__and3_1
XFILLER_0_78_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09505_ _10734_/A _09505_/B vssd1 vssd1 vccd1 vccd1 _09860_/A sky130_fd_sc_hd__or2_4
XANTENNA__13073__B _13129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11635__A2 fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07697_ _07347_/X _08118_/B _13151_/A fanout39/X vssd1 vssd1 vccd1 vccd1 _07698_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09436_ _09694_/A _13129_/A _09463_/S vssd1 vssd1 vccd1 vccd1 _09436_/X sky130_fd_sc_hd__mux2_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ _09367_/A _09367_/B vssd1 vssd1 vccd1 vccd1 _09368_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_81_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08318_ _08746_/A _08318_/B vssd1 vssd1 vccd1 vccd1 _08322_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08183__A _10266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09298_ _09186_/A _09186_/B _09185_/A vssd1 vssd1 vccd1 vccd1 _09308_/A sky130_fd_sc_hd__a21o_2
XANTENNA_50 reg2_val[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_61 reg2_val[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_72 _13036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08249_ _13147_/A fanout28/X _08395_/B _13149_/A vssd1 vssd1 vccd1 vccd1 _08250_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_83 reg1_val[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11260_ _11249_/X _11250_/Y _11259_/X _12710_/B2 _11258_/X vssd1 vssd1 vccd1 vccd1
+ _11260_/X sky130_fd_sc_hd__a221o_1
X_10211_ _10212_/A _10212_/B vssd1 vssd1 vccd1 vccd1 _10213_/A sky130_fd_sc_hd__and2_1
XFILLER_0_120_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11191_ _11191_/A _11191_/B vssd1 vssd1 vccd1 vccd1 _11193_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10374__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10142_ _10142_/A _10142_/B vssd1 vssd1 vccd1 vccd1 _10144_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08319__A2 _07545_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10073_ _11076_/A _10073_/B vssd1 vssd1 vccd1 vccd1 _10074_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11991__B fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10975_ _10976_/A _10976_/B _10976_/C vssd1 vssd1 vccd1 vccd1 _10977_/A sky130_fd_sc_hd__a21o_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12714_ _12714_/A _12714_/B _12714_/C _12701_/X vssd1 vssd1 vccd1 vccd1 _12714_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_85_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13694_ _13700_/CLK hold61/X vssd1 vssd1 vccd1 vccd1 _13694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12645_ _12695_/A _09090_/Y _09097_/A _09095_/Y vssd1 vssd1 vccd1 vccd1 _12645_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_127_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_360 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11512__A _11512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12576_ _12635_/C _12575_/X _09429_/X vssd1 vssd1 vccd1 vccd1 _12576_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11231__B _12372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11527_ _11527_/A _11802_/B vssd1 vssd1 vccd1 vccd1 _11528_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12339__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11458_ _11458_/A _11458_/B vssd1 vssd1 vccd1 vccd1 _11458_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11011__B1 _12657_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10409_ _10410_/A _10409_/B vssd1 vssd1 vccd1 vccd1 _10515_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_68_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11389_ _11288_/A _11288_/C _11288_/B vssd1 vssd1 vccd1 vccd1 _11391_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _13128_/A _13128_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[29] sky130_fd_sc_hd__xnor2_4
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ reg1_val[15] _13059_/B vssd1 vssd1 vccd1 vccd1 _13061_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_84_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07620_ _07620_/A _07620_/B vssd1 vssd1 vccd1 vccd1 _07633_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07172__A _08203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07551_ _07552_/A _07552_/B vssd1 vssd1 vccd1 vccd1 _07911_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_124_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07482_ _07349_/X _07481_/X _07637_/B vssd1 vssd1 vccd1 vccd1 _07486_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_75_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09221_ _09221_/A _09221_/B vssd1 vssd1 vccd1 vccd1 _09223_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11422__A _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09152_ _09153_/A _09153_/B vssd1 vssd1 vccd1 vccd1 _09152_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09443__A0 _13015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08103_ _08101_/A _08101_/B _08102_/Y vssd1 vssd1 vccd1 vccd1 _08997_/A sky130_fd_sc_hd__a21bo_2
XFILLER_0_44_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11250__B1 _12533_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09083_ _08993_/A _08365_/B _08236_/X vssd1 vssd1 vccd1 vccd1 _09086_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout215_A _10456_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08034_ _08104_/A _08104_/B _07967_/X vssd1 vssd1 vccd1 vccd1 _08999_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_24_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11002__B1 _12525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13542__A2 _13555_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12253__A _12253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10356__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09985_ _09985_/A _09985_/B vssd1 vssd1 vccd1 vccd1 _10577_/A sky130_fd_sc_hd__xnor2_4
X_08936_ _08938_/A _08938_/C _08938_/B vssd1 vssd1 vccd1 vccd1 _08964_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__07509__B1 _07572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08867_ _09371_/A _08867_/B vssd1 vssd1 vccd1 vccd1 _08901_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08182__B1 _08246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07818_ _07817_/B _07817_/C _07817_/A vssd1 vssd1 vccd1 vccd1 _07838_/B sky130_fd_sc_hd__o21ba_1
X_08798_ _08799_/A _08799_/B vssd1 vssd1 vccd1 vccd1 _08798_/Y sky130_fd_sc_hd__nand2_1
X_07749_ _07749_/A _07749_/B vssd1 vssd1 vccd1 vccd1 _07772_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_67_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10816__B1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10760_ _12760_/A1 _10745_/X _10759_/X _10737_/X vssd1 vssd1 vccd1 vccd1 _10760_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout30_A _07421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09419_ _09419_/A _09419_/B vssd1 vssd1 vccd1 vccd1 _09421_/B sky130_fd_sc_hd__xnor2_2
X_10691_ _12268_/A fanout25/X fanout23/X fanout46/X vssd1 vssd1 vccd1 vccd1 _10692_/B
+ sky130_fd_sc_hd__o22a_1
X_12430_ _12431_/A _12431_/B vssd1 vssd1 vccd1 vccd1 _12505_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12361_ _12363_/A vssd1 vssd1 vccd1 vccd1 _12361_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11312_ _11311_/A _11311_/B _11311_/C vssd1 vssd1 vccd1 vccd1 _11319_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12292_ _12122_/Y _12290_/B _12442_/B vssd1 vssd1 vccd1 vccd1 _12292_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11243_ reg1_val[12] curr_PC[12] vssd1 vssd1 vccd1 vccd1 _11243_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13533__A2 _13555_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12163__A _12163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11174_ _11174_/A _11174_/B vssd1 vssd1 vccd1 vccd1 _11195_/A sky130_fd_sc_hd__xor2_1
X_10125_ _10125_/A _10125_/B vssd1 vssd1 vccd1 vccd1 _10127_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10056_ _10057_/A _10057_/B vssd1 vssd1 vccd1 vccd1 _10056_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_89_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11507__A _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08088__A _08088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13746_ instruction[9] vssd1 vssd1 vccd1 vccd1 pred_idx[1] sky130_fd_sc_hd__buf_12
XANTENNA__08476__A1 _08806_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10958_ _10958_/A _10958_/B vssd1 vssd1 vccd1 vccd1 _10959_/B sky130_fd_sc_hd__xor2_1
XANTENNA__08476__B2 _08806_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11480__B1 _12657_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13677_ _13684_/CLK _13677_/D vssd1 vssd1 vccd1 vccd1 hold128/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10889_ _10889_/A _10889_/B vssd1 vssd1 vccd1 vccd1 _10889_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12338__A _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12628_ _12506_/A _12567_/X _12569_/B vssd1 vssd1 vccd1 vccd1 _12628_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10035__A1 _10457_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08779__A2 _08778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12559_ _12666_/A _12559_/B vssd1 vssd1 vccd1 vccd1 _12560_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06770__S _07135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold106 hold106/A vssd1 vssd1 vccd1 vccd1 hold106/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 hold117/A vssd1 vssd1 vccd1 vccd1 hold117/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold128 hold128/A vssd1 vssd1 vccd1 vccd1 hold128/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 hold139/A vssd1 vssd1 vccd1 vccd1 hold139/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07739__B1 _10814_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ _09940_/A _09770_/B vssd1 vssd1 vccd1 vccd1 _09774_/A sky130_fd_sc_hd__xnor2_1
X_06982_ _07556_/A vssd1 vssd1 vccd1 vccd1 _07557_/A sky130_fd_sc_hd__inv_2
XANTENNA__12801__A _12982_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ _08700_/A _08700_/B _08720_/Y vssd1 vssd1 vccd1 vccd1 _08726_/A sky130_fd_sc_hd__o21ai_4
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09900__A1 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08652_ _08650_/A _08650_/B _08651_/X vssd1 vssd1 vccd1 vccd1 _08694_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__09900__B2 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07603_ _07603_/A _07603_/B vssd1 vssd1 vccd1 vccd1 _07620_/A sky130_fd_sc_hd__xnor2_2
X_08583_ _08821_/B2 _10049_/A2 _09173_/B2 _08821_/A1 vssd1 vssd1 vccd1 vccd1 _08584_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout165_A _13207_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07534_ _07321_/X _07533_/X _07535_/B vssd1 vssd1 vccd1 vccd1 _07537_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_119_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07465_ _11508_/A _07467_/B vssd1 vssd1 vccd1 vccd1 _07474_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_119_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09204_ _07961_/X _08998_/B _07960_/X vssd1 vssd1 vccd1 vccd1 _09204_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07396_ _12417_/A _07401_/B vssd1 vssd1 vccd1 vccd1 _07396_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_56_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09135_ _09135_/A _09135_/B vssd1 vssd1 vccd1 vccd1 _09139_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_72_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09066_ _12130_/B _12131_/A vssd1 vssd1 vccd1 vccd1 _09066_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_4_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08017_ _08015_/Y _08095_/B _08009_/X vssd1 vssd1 vccd1 vccd1 _08039_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10329__A2 _11793_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09968_ _09968_/A _09968_/B vssd1 vssd1 vccd1 vccd1 _09981_/A sky130_fd_sc_hd__xor2_4
XANTENNA__07805__A _10095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08919_ _09948_/A _08919_/B vssd1 vssd1 vccd1 vccd1 _08920_/C sky130_fd_sc_hd__xnor2_1
X_09899_ _09736_/A _09735_/Y _09733_/Y vssd1 vssd1 vccd1 vccd1 _09914_/A sky130_fd_sc_hd__a21bo_1
X_11930_ _11929_/A _11929_/B _11931_/A vssd1 vssd1 vccd1 vccd1 _12014_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__10231__A _11825_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10501__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11861_ _12035_/A _11861_/B vssd1 vssd1 vccd1 vccd1 _12163_/C sky130_fd_sc_hd__xor2_4
X_13600_ hold170/X _13599_/X _13605_/A vssd1 vssd1 vccd1 vccd1 hold171/A sky130_fd_sc_hd__o21a_1
X_10812_ _10813_/A _10813_/B vssd1 vssd1 vccd1 vccd1 _10812_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_79_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11792_ _11768_/Y _11791_/X _07152_/X vssd1 vssd1 vccd1 vccd1 _11792_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__08636__A _08951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10265__A1 _11732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13531_ _13531_/A _13531_/B vssd1 vssd1 vccd1 vccd1 _13531_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__10265__B2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10743_ _09466_/X _09481_/X _11472_/S vssd1 vssd1 vccd1 vccd1 _10743_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_55_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13462_ hold285/A _13461_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13462_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10674_ _11072_/A _10674_/B vssd1 vssd1 vccd1 vccd1 _10676_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12413_ _12413_/A _12764_/B vssd1 vssd1 vccd1 vccd1 _12414_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11997__A _11997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13393_ _10239_/A _13419_/A2 hold99/X vssd1 vssd1 vccd1 vccd1 hold100/A sky130_fd_sc_hd__o21a_1
XFILLER_0_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12344_ _12344_/A _12344_/B vssd1 vssd1 vccd1 vccd1 _12345_/B sky130_fd_sc_hd__or2_1
XANTENNA__08630__A1 _08933_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08630__B2 _07175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13506__A2 _13506_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12275_ _12276_/A _12276_/B vssd1 vssd1 vccd1 vccd1 _12358_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__11517__A1 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11517__B2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11226_ _10978_/Y _11454_/A _11224_/Y vssd1 vssd1 vccd1 vccd1 _11226_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_120_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11157_ _11157_/A fanout6/X vssd1 vssd1 vccd1 vccd1 _11157_/Y sky130_fd_sc_hd__nand2_1
X_10108_ _10109_/A _10109_/B vssd1 vssd1 vccd1 vccd1 _10108_/X sky130_fd_sc_hd__and2_1
X_11088_ _10931_/A _10931_/B _10928_/Y vssd1 vssd1 vccd1 vccd1 _11091_/A sky130_fd_sc_hd__o21bai_1
XANTENNA__08146__B1 _08868_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10039_ _11866_/A _09996_/Y _10023_/X _10038_/X vssd1 vssd1 vccd1 vccd1 _10039_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13452__A fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13171__B _13191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13729_ _13731_/CLK _13729_/D vssd1 vssd1 vccd1 vccd1 hold269/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07250_ _10239_/A _07250_/B vssd1 vssd1 vccd1 vccd1 _07261_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06880__B1 _06906_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07181_ _07186_/B _07186_/C vssd1 vssd1 vccd1 vccd1 _07192_/A sky130_fd_sc_hd__and2_1
XFILLER_0_6_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09822_ _09822_/A _09822_/B vssd1 vssd1 vccd1 vccd1 _09824_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__09824__B _09824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09753_ _09753_/A _09753_/B _09753_/C vssd1 vssd1 vccd1 vccd1 _09754_/B sky130_fd_sc_hd__nand3_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06965_ _06963_/Y _06966_/B vssd1 vssd1 vccd1 vccd1 _07095_/A sky130_fd_sc_hd__and2b_1
XANTENNA__12469__C1 _12795_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08704_ _09674_/S _08704_/B vssd1 vssd1 vccd1 vccd1 _08742_/B sky130_fd_sc_hd__nor2_1
X_09684_ _09680_/X _09683_/X _10176_/A vssd1 vssd1 vccd1 vccd1 _09684_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09885__B1 _09885_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06896_ _06936_/B _12990_/B vssd1 vssd1 vccd1 vccd1 _06896_/Y sky130_fd_sc_hd__nor2_1
X_08635_ _08866_/B2 _09173_/B2 _11047_/A _08950_/B vssd1 vssd1 vccd1 vccd1 _08636_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ _08571_/A _08571_/B vssd1 vssd1 vccd1 vccd1 _08566_/X sky130_fd_sc_hd__or2_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13433__A1 _12421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10247__A1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout12 fanout13/X vssd1 vssd1 vccd1 vccd1 fanout12/X sky130_fd_sc_hd__buf_6
XANTENNA__10247__B2 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07517_ _07517_/A _07517_/B _07517_/C _07517_/D vssd1 vssd1 vccd1 vccd1 _07524_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_0_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout23 _07474_/Y vssd1 vssd1 vccd1 vccd1 fanout23/X sky130_fd_sc_hd__clkbuf_8
X_08497_ _08495_/A _08495_/B _08557_/A vssd1 vssd1 vccd1 vccd1 _08521_/A sky130_fd_sc_hd__a21bo_1
Xfanout34 fanout35/X vssd1 vssd1 vccd1 vccd1 fanout34/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_49_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout45 _07242_/X vssd1 vssd1 vccd1 vccd1 fanout45/X sky130_fd_sc_hd__buf_6
XFILLER_0_92_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout56 _07197_/X vssd1 vssd1 vccd1 vccd1 fanout56/X sky130_fd_sc_hd__buf_6
Xfanout67 _07577_/X vssd1 vssd1 vccd1 vccd1 _08778_/B sky130_fd_sc_hd__buf_6
X_07448_ _07186_/B _07186_/C _07476_/B vssd1 vssd1 vccd1 vccd1 _07448_/Y sky130_fd_sc_hd__a21oi_1
Xfanout89 _11507_/A vssd1 vssd1 vccd1 vccd1 _11913_/A sky130_fd_sc_hd__buf_8
XFILLER_0_17_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07379_ reg1_val[26] _07634_/B _07634_/C _07378_/D reg1_val[27] vssd1 vssd1 vccd1
+ vccd1 _12598_/B sky130_fd_sc_hd__o41a_1
X_09118_ _07900_/A _07899_/B _07899_/A vssd1 vssd1 vccd1 vccd1 _09119_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_44_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08191__A _09591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10390_ _10390_/A _10390_/B vssd1 vssd1 vccd1 vccd1 _10391_/B sky130_fd_sc_hd__or2_1
X_09049_ _09049_/A _09049_/B vssd1 vssd1 vccd1 vccd1 _09049_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12060_ hold275/A _12058_/X _12059_/Y vssd1 vssd1 vccd1 vccd1 _12060_/Y sky130_fd_sc_hd__a21oi_1
X_11011_ _07456_/A _11793_/B _12657_/B1 reg1_val[10] vssd1 vssd1 vccd1 vccd1 _11011_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11057__A _11709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12962_ _12948_/B _12956_/B _12956_/A vssd1 vssd1 vccd1 vccd1 _12963_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__09750__A _10522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11913_ _11913_/A _11913_/B vssd1 vssd1 vccd1 vccd1 _11915_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_59_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12893_ _12893_/A _12893_/B _12893_/C vssd1 vssd1 vccd1 vccd1 _12894_/B sky130_fd_sc_hd__nand3_1
X_11844_ _11845_/B _11845_/A vssd1 vssd1 vccd1 vccd1 _11844_/X sky130_fd_sc_hd__and2b_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _11682_/A _11679_/Y _11681_/B vssd1 vssd1 vccd1 vccd1 _11779_/A sky130_fd_sc_hd__o21a_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10726_ _10726_/A _10726_/B _10726_/C _09656_/C vssd1 vssd1 vccd1 vccd1 _10727_/D
+ sky130_fd_sc_hd__or4b_1
X_13514_ _13514_/A _13514_/B vssd1 vssd1 vccd1 vccd1 _13514_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13445_ _12764_/B _13445_/A2 hold124/X vssd1 vssd1 vccd1 vccd1 hold125/A sky130_fd_sc_hd__o21a_1
X_10657_ fanout15/X _11527_/A _11638_/A fanout31/X vssd1 vssd1 vccd1 vccd1 _10658_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13376_ hold219/A _13599_/D _13584_/B hold197/X vssd1 vssd1 vccd1 vccd1 hold198/A
+ sky130_fd_sc_hd__a22o_1
X_10588_ _10734_/A _10588_/B _10588_/C vssd1 vssd1 vccd1 vccd1 _10588_/X sky130_fd_sc_hd__and3_1
XFILLER_0_23_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12327_ _12327_/A _12477_/C _12327_/C vssd1 vssd1 vccd1 vccd1 _12327_/X sky130_fd_sc_hd__or3_1
XFILLER_0_23_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12258_ _12258_/A _12258_/B vssd1 vssd1 vccd1 vccd1 _12259_/B sky130_fd_sc_hd__nand2_1
X_11209_ _11209_/A _11209_/B _11209_/C vssd1 vssd1 vccd1 vccd1 _11210_/B sky130_fd_sc_hd__and3_1
XANTENNA__13360__B1 _13450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12189_ _12189_/A _12764_/B vssd1 vssd1 vccd1 vccd1 _12190_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11910__A1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11910__B2 _08118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08119__B1 _11638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06750_ _11126_/A vssd1 vssd1 vccd1 vccd1 _07531_/A sky130_fd_sc_hd__inv_2
XANTENNA__11123__C1 _12047_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09867__B1 _09507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10477__A1 _12047_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08420_ _09940_/A _08420_/B vssd1 vssd1 vccd1 vccd1 _08427_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08276__A _08951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08351_ _08351_/A _08351_/B vssd1 vssd1 vccd1 vccd1 _08353_/B sky130_fd_sc_hd__or2_1
XFILLER_0_86_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07302_ _13015_/A _07320_/C reg1_val[8] vssd1 vssd1 vccd1 vccd1 _10750_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08282_ _08282_/A _08282_/B vssd1 vssd1 vccd1 vccd1 _08345_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_34_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07233_ reg1_val[2] _07535_/B _07232_/X vssd1 vssd1 vccd1 vccd1 _07235_/B sky130_fd_sc_hd__a21o_1
XANTENNA__10745__S _12648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09398__A2 _07451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07164_ reg1_val[3] _09871_/A vssd1 vssd1 vccd1 vccd1 _07164_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07095_ _07095_/A _10592_/A _07095_/C _07094_/X vssd1 vssd1 vccd1 vccd1 _07098_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_112_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12154__A1 _12759_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout202 _07166_/Y vssd1 vssd1 vccd1 vccd1 _09951_/A sky130_fd_sc_hd__buf_6
XANTENNA__12154__B2 _12537_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout213 _10007_/S vssd1 vssd1 vccd1 vccd1 _10005_/S sky130_fd_sc_hd__clkbuf_8
Xfanout224 _06989_/X vssd1 vssd1 vccd1 vccd1 _12225_/A sky130_fd_sc_hd__buf_2
Xfanout235 _09429_/X vssd1 vssd1 vccd1 vccd1 _11955_/A sky130_fd_sc_hd__buf_4
XFILLER_0_5_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout246 _06928_/B vssd1 vssd1 vccd1 vccd1 _06936_/B sky130_fd_sc_hd__buf_8
X_09805_ _09806_/A _09806_/B vssd1 vssd1 vccd1 vccd1 _09807_/A sky130_fd_sc_hd__and2_1
Xfanout257 _09511_/X vssd1 vssd1 vccd1 vccd1 _12754_/C sky130_fd_sc_hd__buf_4
Xfanout268 _07110_/A vssd1 vssd1 vccd1 vccd1 _06873_/B1 sky130_fd_sc_hd__buf_4
X_07997_ _07997_/A _07997_/B vssd1 vssd1 vccd1 vccd1 _08093_/B sky130_fd_sc_hd__xnor2_2
Xfanout279 _13444_/C1 vssd1 vssd1 vccd1 vccd1 _13430_/C1 sky130_fd_sc_hd__buf_2
XANTENNA__07581__A1 _13174_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07581__B2 _07545_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13103__B1 _13129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09736_ _09736_/A _09736_/B vssd1 vssd1 vccd1 vccd1 _09738_/A sky130_fd_sc_hd__xor2_4
X_06948_ _07531_/A _07471_/A vssd1 vssd1 vccd1 vccd1 _11138_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09570__A _10078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09667_ _09444_/X _09446_/X _09674_/S vssd1 vssd1 vccd1 vccd1 _09667_/X sky130_fd_sc_hd__mux2_1
X_06879_ _06886_/A _13000_/B vssd1 vssd1 vccd1 vccd1 _06879_/Y sky130_fd_sc_hd__nor2_1
X_08618_ _08980_/A _08980_/B vssd1 vssd1 vccd1 vccd1 _08981_/A sky130_fd_sc_hd__or2_1
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11605__A _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _09598_/A _09598_/B vssd1 vssd1 vccd1 vccd1 _09599_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_49_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07090__A _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08549_ _08577_/A _08547_/Y _08536_/Y vssd1 vssd1 vccd1 vccd1 _08560_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11560_ _11561_/A _11561_/B vssd1 vssd1 vccd1 vccd1 _11560_/X sky130_fd_sc_hd__and2_1
XFILLER_0_80_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10511_ _10511_/A _10511_/B vssd1 vssd1 vccd1 vccd1 _10513_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11491_ _12867_/S _11487_/X _11488_/X _11490_/Y vssd1 vssd1 vccd1 vccd1 dest_val[14]
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_80_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13230_ hold255/X hold103/X vssd1 vssd1 vccd1 vccd1 _13552_/B sky130_fd_sc_hd__nand2b_1
X_10442_ _12130_/A _10344_/X _10441_/X vssd1 vssd1 vccd1 vccd1 _10442_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13161_ hold68/X _13193_/B vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__or2_1
XANTENNA__13590__B1 _13584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08061__A2 _07203_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10373_ _11731_/A _10373_/B vssd1 vssd1 vccd1 vccd1 _10380_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10943__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12112_ _12112_/A _12112_/B vssd1 vssd1 vccd1 vccd1 _12114_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_20_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13092_ reg1_val[22] _13129_/B vssd1 vssd1 vccd1 vccd1 _13093_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_20_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13342__B1 _13506_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12043_ _12043_/A _12043_/B vssd1 vssd1 vccd1 vccd1 _12043_/Y sky130_fd_sc_hd__xnor2_1
X_12945_ _12951_/B _12945_/B vssd1 vssd1 vccd1 vccd1 new_PC[21] sky130_fd_sc_hd__xnor2_4
XFILLER_0_62_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12876_ _13036_/B _12876_/B vssd1 vssd1 vccd1 vccd1 _12877_/B sky130_fd_sc_hd__or2_1
XFILLER_0_56_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11408__B1 _09146_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11827_ _12417_/A _11827_/B vssd1 vssd1 vccd1 vccd1 _11829_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _11758_/A _11758_/B _11758_/C vssd1 vssd1 vccd1 vccd1 _11759_/B sky130_fd_sc_hd__nand3_1
XANTENNA__08824__A _09659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10709_ _10710_/A _10710_/B vssd1 vssd1 vccd1 vccd1 _10709_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_70_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11689_ _06912_/B _09515_/Y _11586_/B _06910_/A _11688_/Y vssd1 vssd1 vccd1 vccd1
+ _11689_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_71_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13428_ hold146/A _06744_/Y _13444_/B1 hold70/X _13430_/C1 vssd1 vssd1 vccd1 vccd1
+ hold71/A sky130_fd_sc_hd__o221a_1
XFILLER_0_24_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13359_ _13359_/A hold178/X vssd1 vssd1 vccd1 vccd1 hold179/A sky130_fd_sc_hd__and2_1
XFILLER_0_11_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07920_ _07921_/A _07921_/B vssd1 vssd1 vccd1 vccd1 _09179_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09552__A2 wire122/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07851_ _07851_/A _07851_/B vssd1 vssd1 vccd1 vccd1 _07963_/B sky130_fd_sc_hd__xor2_4
X_06802_ _06802_/A _06802_/B vssd1 vssd1 vccd1 vccd1 _12581_/A sky130_fd_sc_hd__nor2_2
X_07782_ _07782_/A _07782_/B vssd1 vssd1 vccd1 vccd1 _07783_/B sky130_fd_sc_hd__xnor2_2
X_09521_ _09524_/A _09523_/B vssd1 vssd1 vccd1 vccd1 _09521_/Y sky130_fd_sc_hd__nor2_4
X_09452_ reg1_val[15] reg1_val[16] _09463_/S vssd1 vssd1 vccd1 vccd1 _09452_/X sky130_fd_sc_hd__mux2_1
X_08403_ _08403_/A _08403_/B _08403_/C vssd1 vssd1 vccd1 vccd1 _08405_/A sky130_fd_sc_hd__or3_1
XFILLER_0_93_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09383_ _09910_/A1 fanout9/X fanout4/X _09604_/A vssd1 vssd1 vccd1 vccd1 _09384_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08334_ _08380_/A _08380_/B _08330_/Y vssd1 vssd1 vccd1 vccd1 _08340_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_117_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10622__A1 _12759_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08265_ _08873_/A2 fanout85/X fanout82/X _08891_/B vssd1 vssd1 vccd1 vccd1 _08266_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07216_ _07252_/C _07217_/B vssd1 vssd1 vccd1 vccd1 _12496_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_116_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08196_ _09948_/A _08196_/B vssd1 vssd1 vccd1 vccd1 _08201_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07147_ _12578_/A is_load _06928_/B _07144_/X vssd1 vssd1 vccd1 vccd1 _07148_/B sky130_fd_sc_hd__a22o_2
XANTENNA__09240__A1 _11732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09240__B2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09791__A2 _07522_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07078_ _07077_/A _07077_/B _12452_/A vssd1 vssd1 vccd1 vccd1 _07079_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_100_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13324__B1 _13450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11886__B1 _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07554__A1 _10915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07554__B2 _08486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10153__A3 _10577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09719_ _09658_/X _09662_/X _09718_/X _12327_/A vssd1 vssd1 vccd1 vccd1 _09719_/X
+ sky130_fd_sc_hd__o31a_1
X_10991_ _11463_/A _06962_/Y _07039_/Y _10990_/Y vssd1 vssd1 vccd1 vccd1 _10992_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_96_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _12730_/A _12730_/B _12730_/C vssd1 vssd1 vccd1 vccd1 _12731_/C sky130_fd_sc_hd__nor3_1
XANTENNA__07857__A2 _08246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_6_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13736_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _12660_/X _12661_/B _12661_/C _12661_/D vssd1 vssd1 vccd1 vccd1 _12661_/X
+ sky130_fd_sc_hd__and4b_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ fanout29/X _07891_/X _09146_/Y fanout27/X vssd1 vssd1 vccd1 vccd1 _11613_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08806__A1 _09703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07609__A2 _10536_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12592_ hold166/A _12592_/B vssd1 vssd1 vccd1 vccd1 _12650_/B sky130_fd_sc_hd__or2_1
XANTENNA__08806__B2 _07399_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11543_ _11543_/A _11543_/B vssd1 vssd1 vccd1 vccd1 _11544_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_9_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07490__B1 _07476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11474_ _11471_/X _11473_/X _12225_/A vssd1 vssd1 vccd1 vccd1 _11474_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_80_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13213_ hold247/X hold30/X vssd1 vssd1 vccd1 vccd1 _13214_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_33_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10425_ _10426_/B _10426_/A vssd1 vssd1 vccd1 vccd1 _10425_/X sky130_fd_sc_hd__and2b_1
XANTENNA__09231__A1 _07203_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09231__B2 _07230_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13144_ _12764_/B _13598_/C hold18/X _13605_/A vssd1 vssd1 vccd1 vccd1 _13608_/D
+ sky130_fd_sc_hd__o211a_1
X_10356_ fanout47/X fanout83/X fanout79/X fanout45/X vssd1 vssd1 vccd1 vccd1 _10357_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13075_ _13081_/A _13081_/B _13129_/B _07435_/B vssd1 vssd1 vccd1 vccd1 _13076_/B
+ sky130_fd_sc_hd__a2bb2o_2
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10287_ _10287_/A _10287_/B vssd1 vssd1 vccd1 vccd1 _10288_/B sky130_fd_sc_hd__xor2_2
X_12026_ _12027_/A _12027_/B vssd1 vssd1 vccd1 vccd1 _12120_/A sky130_fd_sc_hd__or2_1
XFILLER_0_88_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10787__C _10787_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12928_ _12956_/A _12929_/B vssd1 vssd1 vccd1 vccd1 _12938_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_87_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12859_ _12865_/B _12859_/B vssd1 vssd1 vccd1 vccd1 new_PC[8] sky130_fd_sc_hd__and2_4
XFILLER_0_29_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12076__A _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_3_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08050_ _08054_/A _08054_/B vssd1 vssd1 vccd1 vccd1 _08050_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07001_ reg1_val[4] _10603_/S vssd1 vssd1 vccd1 vccd1 _07001_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_114_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07379__A4 _07378_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08952_ _08954_/A _08953_/B vssd1 vssd1 vccd1 vccd1 _08960_/A sky130_fd_sc_hd__nand2_1
X_07903_ _10814_/A1 fanout68/X fanout66/X fanout42/X vssd1 vssd1 vccd1 vccd1 _07904_/B
+ sky130_fd_sc_hd__o22a_1
X_08883_ _08861_/A _08861_/B _08861_/C vssd1 vssd1 vccd1 vccd1 _08883_/X sky130_fd_sc_hd__o21a_1
X_07834_ _07994_/A _12421_/A _07994_/B vssd1 vssd1 vccd1 vccd1 _07835_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07765_ _10119_/A _07765_/B vssd1 vssd1 vccd1 vccd1 _07766_/C sky130_fd_sc_hd__xnor2_1
X_09504_ _10734_/A _09505_/B vssd1 vssd1 vccd1 vccd1 _09504_/Y sky130_fd_sc_hd__nor2_2
X_07696_ _07696_/A _07696_/B vssd1 vssd1 vccd1 vccd1 _07707_/A sky130_fd_sc_hd__xor2_1
X_09435_ _12738_/S _09505_/B vssd1 vssd1 vccd1 vccd1 _09435_/X sky130_fd_sc_hd__or2_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09366_ _09367_/A _09367_/B vssd1 vssd1 vccd1 vccd1 _09368_/A sky130_fd_sc_hd__and2_1
XFILLER_0_19_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08317_ _09885_/B1 _10538_/A _08778_/B _10049_/A2 vssd1 vssd1 vccd1 vccd1 _08318_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09297_ _09297_/A _09297_/B vssd1 vssd1 vccd1 vccd1 _09310_/A sky130_fd_sc_hd__xor2_4
XANTENNA_40 reg1_val[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_51 reg2_val[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_62 reg2_val[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08248_ _08251_/A _08251_/B vssd1 vssd1 vccd1 vccd1 _08252_/A sky130_fd_sc_hd__nor2_1
XANTENNA_73 reg1_val[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_84 reg1_val[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08179_ _08178_/B _08178_/C _08178_/A vssd1 vssd1 vccd1 vccd1 _08220_/A sky130_fd_sc_hd__o21bai_2
X_10210_ _12253_/A _10210_/B vssd1 vssd1 vccd1 vccd1 _10212_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11190_ _11191_/A _11191_/B vssd1 vssd1 vccd1 vccd1 _11315_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_30_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10141_ _10142_/B _10142_/A vssd1 vssd1 vccd1 vccd1 _10141_/Y sky130_fd_sc_hd__nand2b_1
X_10072_ fanout49/X fanout68/X fanout66/X fanout51/X vssd1 vssd1 vccd1 vccd1 _10073_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08639__A _10944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07543__A _07544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10974_ _10974_/A _10974_/B vssd1 vssd1 vccd1 vccd1 _10976_/C sky130_fd_sc_hd__xor2_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12713_ _12703_/Y _12704_/X _12712_/X vssd1 vssd1 vccd1 vccd1 _12714_/C sky130_fd_sc_hd__o21ai_1
X_13693_ _13693_/CLK _13693_/D vssd1 vssd1 vccd1 vccd1 hold138/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12644_ _09097_/A _09095_/Y _12695_/A _09090_/Y vssd1 vssd1 vccd1 vccd1 _12644_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12575_ _12733_/A _12635_/A _12635_/B _12735_/A1 vssd1 vssd1 vccd1 vccd1 _12575_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_26_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11231__C _11600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11526_ _11401_/A _11401_/B _11399_/Y vssd1 vssd1 vccd1 vccd1 _11528_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_53_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12339__A1 _12496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12339__B2 _12413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11457_ _11458_/B vssd1 vssd1 vccd1 vccd1 _11457_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_111_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10408_ _10410_/B vssd1 vssd1 vccd1 vccd1 _10409_/B sky130_fd_sc_hd__inv_2
XFILLER_0_68_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07215__B1 _07521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11388_ _11388_/A _11388_/B vssd1 vssd1 vccd1 vccd1 _11391_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_104_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10339_ _11866_/A _10306_/Y _10307_/X _10338_/X _10305_/Y vssd1 vssd1 vccd1 vccd1
+ _10339_/X sky130_fd_sc_hd__a311o_1
X_13127_ _13120_/A _13123_/B _13120_/B vssd1 vssd1 vccd1 vccd1 _13128_/B sky130_fd_sc_hd__a21bo_2
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _13061_/B _13058_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[14] sky130_fd_sc_hd__and2_4
X_12009_ _12010_/A _12010_/B vssd1 vssd1 vccd1 vccd1 _12009_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__06768__S _07135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07550_ _11286_/A _07550_/B vssd1 vssd1 vccd1 vccd1 _07552_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09140__B1 _07597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07481_ _07377_/A _07337_/B _07483_/A vssd1 vssd1 vccd1 vccd1 _07481_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_124_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09220_ _09220_/A _09220_/B vssd1 vssd1 vccd1 vccd1 _09221_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_8_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09151_ _09151_/A _09151_/B vssd1 vssd1 vccd1 vccd1 _09153_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_44_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08102_ _08166_/B _08166_/A vssd1 vssd1 vccd1 vccd1 _08102_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_71_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09082_ _09082_/A _09082_/B _09082_/C vssd1 vssd1 vccd1 vccd1 _09082_/X sky130_fd_sc_hd__or3_1
XANTENNA__07454__B1 _07476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08033_ _08033_/A _08033_/B vssd1 vssd1 vccd1 vccd1 _08104_/B sky130_fd_sc_hd__xor2_4
XANTENNA_fanout110_A _07495_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout208_A _09671_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09984_ _09985_/A _09985_/B vssd1 vssd1 vccd1 vccd1 _09984_/X sky130_fd_sc_hd__and2_1
XFILLER_0_110_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08935_ _08929_/B _08928_/C _08928_/B vssd1 vssd1 vccd1 vccd1 _08938_/C sky130_fd_sc_hd__a21o_1
XANTENNA__13365__A _13543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08866_ _08950_/B _08866_/A2 _08923_/B1 _08866_/B2 vssd1 vssd1 vccd1 vccd1 _08867_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_99_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08182__A1 _09671_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08182__B2 _08873_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07363__A _12515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07817_ _07817_/A _07817_/B _07817_/C vssd1 vssd1 vccd1 vccd1 _08024_/A sky130_fd_sc_hd__or3_1
X_08797_ _09659_/B _08797_/B vssd1 vssd1 vccd1 vccd1 _08799_/B sky130_fd_sc_hd__xnor2_1
X_07748_ _07747_/A _07747_/B _07776_/A vssd1 vssd1 vccd1 vccd1 _07748_/X sky130_fd_sc_hd__o21a_1
XANTENNA__12266__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09131__B1 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10816__A1 _07299_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07679_ _10263_/A _07679_/B vssd1 vssd1 vccd1 vccd1 _07714_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11613__A _11913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09418_ _09304_/A _09304_/B _09302_/Y vssd1 vssd1 vccd1 vccd1 _09419_/B sky130_fd_sc_hd__a21boi_4
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10690_ _10690_/A vssd1 vssd1 vccd1 vccd1 _10699_/A sky130_fd_sc_hd__inv_2
XFILLER_0_125_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09349_ _09559_/B _09349_/B vssd1 vssd1 vccd1 vccd1 _09390_/A sky130_fd_sc_hd__nand2_1
X_12360_ _12362_/A _12362_/B _12362_/C vssd1 vssd1 vccd1 vccd1 _12363_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_7_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08922__A _09371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11311_ _11311_/A _11311_/B _11311_/C vssd1 vssd1 vccd1 vccd1 _11319_/A sky130_fd_sc_hd__or3_1
X_12291_ _12121_/A _12202_/A _12365_/B vssd1 vssd1 vccd1 vccd1 _12442_/B sky130_fd_sc_hd__a21o_1
X_11242_ reg1_val[12] curr_PC[12] vssd1 vssd1 vccd1 vccd1 _11242_/X sky130_fd_sc_hd__or2_1
XFILLER_0_120_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12163__B _12163_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11173_ _11174_/B vssd1 vssd1 vccd1 vccd1 _11173_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10124_ _10125_/A _10125_/B vssd1 vssd1 vccd1 vccd1 _10124_/X sky130_fd_sc_hd__and2_1
XFILLER_0_100_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10055_ _12092_/A _10055_/B vssd1 vssd1 vccd1 vccd1 _10057_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10504__B1 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09370__B1 _10536_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07273__A _09948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09122__B1 _10536_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13745_ instruction[8] vssd1 vssd1 vccd1 vccd1 pred_idx[0] sky130_fd_sc_hd__buf_12
XANTENNA__08476__A2 _07492_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10957_ _10958_/B _10958_/A vssd1 vssd1 vccd1 vccd1 _11087_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_97_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13676_ _13684_/CLK _13676_/D vssd1 vssd1 vccd1 vccd1 hold101/A sky130_fd_sc_hd__dfxtp_1
X_10888_ _10888_/A _10888_/B vssd1 vssd1 vccd1 vccd1 _10893_/D sky130_fd_sc_hd__or2_1
XFILLER_0_66_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12627_ _12627_/A _12681_/A vssd1 vssd1 vccd1 vccd1 _12730_/B sky130_fd_sc_hd__or2_1
XFILLER_0_109_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10035__A2 _11793_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12558_ _12558_/A _12558_/B vssd1 vssd1 vccd1 vccd1 _12559_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08832__A _10542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10440__C1 _10981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11509_ _11510_/A _11510_/B vssd1 vssd1 vccd1 vccd1 _11509_/X sky130_fd_sc_hd__and2_1
Xhold107 hold136/X vssd1 vssd1 vccd1 vccd1 hold107/X sky130_fd_sc_hd__dlygate4sd3_1
X_12489_ _12560_/A _12489_/B vssd1 vssd1 vccd1 vccd1 _12491_/C sky130_fd_sc_hd__nor2_1
Xhold118 hold118/A vssd1 vssd1 vccd1 vccd1 hold118/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 hold129/A vssd1 vssd1 vccd1 vccd1 hold129/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13169__B _13193_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07739__A1 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07739__B2 _10235_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ _06936_/A _06928_/B _13015_/B _06980_/X vssd1 vssd1 vccd1 vccd1 _07556_/A
+ sky130_fd_sc_hd__a31o_4
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08720_ _08727_/A _08727_/B vssd1 vssd1 vccd1 vccd1 _08720_/Y sky130_fd_sc_hd__nand2b_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08279__A _10266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07183__A _10889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08651_ _08660_/B _08660_/A vssd1 vssd1 vccd1 vccd1 _08651_/X sky130_fd_sc_hd__and2b_1
XANTENNA__09900__A2 _11423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07602_ _07603_/A _07603_/B vssd1 vssd1 vccd1 vccd1 _07874_/B sky130_fd_sc_hd__or2_1
X_08582_ _08644_/B _08582_/B vssd1 vssd1 vccd1 vccd1 _08645_/A sky130_fd_sc_hd__and2b_1
XANTENNA__12248__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12799__A1 _07398_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07533_ _07531_/A _07571_/A _07535_/A vssd1 vssd1 vccd1 vccd1 _07533_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_9_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07675__B1 _08246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07464_ _11281_/A _07467_/B vssd1 vssd1 vccd1 vccd1 _07473_/A sky130_fd_sc_hd__and2_1
XFILLER_0_29_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09203_ _09203_/A _09203_/B vssd1 vssd1 vccd1 vccd1 _09825_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_119_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07395_ _07395_/A _07395_/B _07395_/C _07395_/D vssd1 vssd1 vccd1 vccd1 _07401_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_8_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09134_ _11286_/A _09134_/B vssd1 vssd1 vccd1 vccd1 _09135_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09065_ _09068_/A _09065_/B vssd1 vssd1 vccd1 vccd1 _09065_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_32_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08016_ _08016_/A _08016_/B vssd1 vssd1 vccd1 vccd1 _08095_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09573__A _10095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09967_ _09967_/A _09967_/B vssd1 vssd1 vccd1 vccd1 _09968_/B sky130_fd_sc_hd__nor2_2
XANTENNA__06953__A2 _06936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08918_ _09703_/B _07175_/X _08933_/B _07399_/Y vssd1 vssd1 vccd1 vccd1 _08919_/B
+ sky130_fd_sc_hd__a22o_1
X_09898_ _09898_/A _09898_/B vssd1 vssd1 vccd1 vccd1 _09968_/A sky130_fd_sc_hd__xnor2_4
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09352__B1 _10235_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08849_ _08849_/A _08849_/B vssd1 vssd1 vccd1 vccd1 _08881_/A sky130_fd_sc_hd__xor2_1
X_11860_ _10984_/B _11454_/Y _11858_/Y _11859_/Y vssd1 vssd1 vccd1 vccd1 _11861_/B
+ sky130_fd_sc_hd__o31a_2
XANTENNA__13436__C1 _13568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09104__B1 _09885_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10811_ _10811_/A _10811_/B vssd1 vssd1 vccd1 vccd1 _10813_/B sky130_fd_sc_hd__xor2_1
X_11791_ _11769_/Y _11770_/X _11774_/Y _12047_/C1 _11790_/X vssd1 vssd1 vccd1 vccd1
+ _11791_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_95_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10265__A2 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13530_ _13539_/A hold258/X vssd1 vssd1 vccd1 vccd1 _13722_/D sky130_fd_sc_hd__and2_1
X_10742_ _10742_/A _10742_/B vssd1 vssd1 vccd1 vccd1 _10742_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06976__A_N _07492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10673_ _07546_/X _10787_/B _10787_/C _10787_/A _12557_/B vssd1 vssd1 vccd1 vccd1
+ _10674_/B sky130_fd_sc_hd__o32a_1
X_13461_ _13461_/A _13461_/B vssd1 vssd1 vccd1 vccd1 _13461_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07418__B1 _07398_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12412_ _12412_/A _12412_/B vssd1 vssd1 vccd1 vccd1 _12414_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09748__A _09748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11997__B _12666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13392_ hold128/A _13416_/A2 _13420_/B1 hold98/X _13430_/C1 vssd1 vssd1 vccd1 vccd1
+ hold99/A sky130_fd_sc_hd__o221a_1
XFILLER_0_23_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12343_ _12344_/A _12344_/B vssd1 vssd1 vccd1 vccd1 _12426_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08630__A2 wire122/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07268__A _10095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12274_ _12189_/A _12764_/B _12190_/A _12188_/A vssd1 vssd1 vccd1 vccd1 _12276_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08918__B1 _08933_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11517__A2 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11225_ _11225_/A _11342_/A vssd1 vssd1 vccd1 vccd1 _11454_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_120_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11156_ _11281_/A _11156_/B vssd1 vssd1 vccd1 vccd1 _11307_/A sky130_fd_sc_hd__xnor2_2
X_10107_ _10522_/B _10107_/B vssd1 vssd1 vccd1 vccd1 _10109_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11518__A _12253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12478__B1 _07108_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11087_ _11087_/A _11087_/B vssd1 vssd1 vccd1 vccd1 _11092_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08146__A1 _10522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08146__B2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10038_ _12047_/C1 _10026_/Y _10037_/Y _10018_/X vssd1 vssd1 vccd1 vccd1 _10038_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__08827__A _08951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13442__A2 _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11989_ fanout38/X _07891_/X fanout10/X fanout36/X vssd1 vssd1 vccd1 vccd1 _11990_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11453__A1 _11224_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13728_ _13731_/CLK _13728_/D vssd1 vssd1 vccd1 vccd1 hold282/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06898__A2_N _06906_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13659_ _13659_/CLK _13659_/D vssd1 vssd1 vccd1 vccd1 hold203/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07877__S _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09658__A _10730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07180_ _07492_/A _07556_/A _07180_/C _07363_/B vssd1 vssd1 vccd1 vccd1 _07186_/C
+ sky130_fd_sc_hd__and4bb_4
XFILLER_0_54_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07178__A _07544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08909__B1 _09659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12812__A _12990_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09821_ _09821_/A _09821_/B vssd1 vssd1 vccd1 vccd1 _09822_/B sky130_fd_sc_hd__xor2_4
XANTENNA__07906__A _10095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09752_ _09753_/A _09753_/B _09753_/C vssd1 vssd1 vccd1 vccd1 _09752_/Y sky130_fd_sc_hd__a21oi_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06964_ reg1_val[9] _10889_/A vssd1 vssd1 vccd1 vccd1 _06966_/B sky130_fd_sc_hd__nand2_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09334__B1 _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08703_ _08746_/A _08703_/B vssd1 vssd1 vccd1 vccd1 _08742_/A sky130_fd_sc_hd__xnor2_2
X_09683_ _09681_/X _09682_/X _10005_/S vssd1 vssd1 vccd1 vccd1 _09683_/X sky130_fd_sc_hd__mux2_1
X_06895_ instruction[0] instruction[1] instruction[2] instruction[27] pred_val vssd1
+ vssd1 vccd1 vccd1 _06895_/Y sky130_fd_sc_hd__o311ai_2
XANTENNA__09885__A1 _07699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11141__B1 _12796_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09885__B2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout275_A _13444_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08634_ _08637_/A _08637_/B vssd1 vssd1 vccd1 vccd1 _08634_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07896__B1 _09949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08565_ _08565_/A _08565_/B vssd1 vssd1 vccd1 vccd1 _08571_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__13433__A2 _13598_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10247__A2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07516_ _07517_/C _07517_/D vssd1 vssd1 vccd1 vccd1 _07516_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_77_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout13 _07878_/X vssd1 vssd1 vccd1 vccd1 fanout13/X sky130_fd_sc_hd__clkbuf_8
X_08496_ _08556_/A _08556_/B vssd1 vssd1 vccd1 vccd1 _08557_/A sky130_fd_sc_hd__or2_1
Xfanout24 fanout25/X vssd1 vssd1 vccd1 vccd1 fanout24/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout35 _07397_/X vssd1 vssd1 vccd1 vccd1 fanout35/X sky130_fd_sc_hd__buf_8
XFILLER_0_76_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout46 _07242_/X vssd1 vssd1 vccd1 vccd1 fanout46/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout57 _07197_/X vssd1 vssd1 vccd1 vccd1 _12103_/A sky130_fd_sc_hd__buf_4
X_07447_ _07453_/B _11800_/A _11913_/A vssd1 vssd1 vccd1 vccd1 _07447_/X sky130_fd_sc_hd__mux2_4
XFILLER_0_92_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout68 _10538_/A vssd1 vssd1 vccd1 vccd1 fanout68/X sky130_fd_sc_hd__buf_6
XFILLER_0_119_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout79 _08580_/B vssd1 vssd1 vccd1 vccd1 fanout79/X sky130_fd_sc_hd__buf_6
XFILLER_0_45_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07378_ reg1_val[26] _07634_/B _07634_/C _07378_/D vssd1 vssd1 vccd1 vccd1 _12534_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_0_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09117_ _07909_/A _07909_/B _07907_/Y vssd1 vssd1 vccd1 vccd1 _09121_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__10507__A _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09048_ _11562_/B _09048_/B _11672_/A vssd1 vssd1 vccd1 vccd1 _09048_/X sky130_fd_sc_hd__and3_1
XFILLER_0_20_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11010_ _11010_/A _12235_/C vssd1 vssd1 vccd1 vccd1 _11010_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07535__B _07535_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12961_ _12961_/A _12961_/B _12961_/C _12961_/D vssd1 vssd1 vccd1 vccd1 _12963_/C
+ sky130_fd_sc_hd__or4_1
XANTENNA__09876__B2 _09523_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11912_ _11913_/A _11913_/B vssd1 vssd1 vccd1 vccd1 _12016_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__07887__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12892_ _12893_/A _12893_/B _12893_/C vssd1 vssd1 vccd1 vccd1 _12900_/B sky130_fd_sc_hd__a21o_1
X_11843_ _11843_/A _11843_/B vssd1 vssd1 vccd1 vccd1 _11845_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13424__A2 _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11774_ _11774_/A _11774_/B vssd1 vssd1 vccd1 vccd1 _11774_/Y sky130_fd_sc_hd__xnor2_2
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _13253_/X _13513_/B vssd1 vssd1 vccd1 vccd1 _13514_/B sky130_fd_sc_hd__nand2b_1
X_10725_ _10441_/A _10441_/B _09881_/A _10156_/A _10156_/B vssd1 vssd1 vccd1 vccd1
+ _10727_/C sky130_fd_sc_hd__a2111o_1
XFILLER_0_67_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13188__A1 _07198_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13444_ hold123/X _13142_/A _13444_/B1 _13704_/Q _13444_/C1 vssd1 vssd1 vccd1 vccd1
+ hold124/A sky130_fd_sc_hd__o221a_1
X_10656_ _10656_/A _10656_/B vssd1 vssd1 vccd1 vccd1 _10668_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10587_ _11562_/A _09018_/A _09018_/B _11866_/A vssd1 vssd1 vccd1 vccd1 _10587_/X
+ sky130_fd_sc_hd__o31a_1
X_13375_ _13547_/A hold220/X vssd1 vssd1 vccd1 vccd1 hold221/A sky130_fd_sc_hd__and2_1
XFILLER_0_23_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_8_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12326_ curr_PC[22] _12325_/C curr_PC[23] vssd1 vssd1 vccd1 vccd1 _12327_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12257_ _12258_/A _12258_/B vssd1 vssd1 vccd1 vccd1 _12336_/A sky130_fd_sc_hd__or2_1
XFILLER_0_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07726__A _09591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11208_ _11209_/A _11209_/B _11209_/C vssd1 vssd1 vccd1 vccd1 _11210_/A sky130_fd_sc_hd__a21oi_1
X_12188_ _12188_/A _12188_/B vssd1 vssd1 vccd1 vccd1 _12190_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11371__B1 _12748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11910__A2 _07597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11139_ _07471_/A _11793_/B _12657_/B1 _11126_/A _11138_/Y vssd1 vssd1 vccd1 vccd1
+ _11139_/X sky130_fd_sc_hd__o221a_1
XANTENNA__08119__A1 _08933_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08119__B2 _07175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07461__A _11281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08350_ _08350_/A _08350_/B _08350_/C vssd1 vssd1 vccd1 vccd1 _08351_/B sky130_fd_sc_hd__and3_1
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07301_ reg1_val[8] _07535_/B vssd1 vssd1 vccd1 vccd1 _07301_/X sky130_fd_sc_hd__and2_1
XFILLER_0_73_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08281_ _10266_/A _08279_/B _08351_/A vssd1 vssd1 vccd1 vccd1 _08345_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_73_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07232_ _07572_/S _09871_/A _09871_/B vssd1 vssd1 vccd1 vccd1 _07232_/X sky130_fd_sc_hd__and3_1
XFILLER_0_73_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07163_ _07535_/B _07160_/Y _07161_/X vssd1 vssd1 vccd1 vccd1 _07163_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07094_ _07094_/A _07094_/B _07094_/C _07094_/D vssd1 vssd1 vccd1 vccd1 _07094_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07339__C _13082_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout203 _12799_/A2 vssd1 vssd1 vccd1 vccd1 _11793_/B sky130_fd_sc_hd__buf_4
Xfanout214 _07020_/X vssd1 vssd1 vccd1 vccd1 _10007_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout225 _06906_/B1 vssd1 vssd1 vccd1 vccd1 _06872_/B1 sky130_fd_sc_hd__buf_4
Xfanout236 _07219_/Y vssd1 vssd1 vccd1 vccd1 _08907_/A sky130_fd_sc_hd__clkbuf_8
X_09804_ _09804_/A _09804_/B vssd1 vssd1 vccd1 vccd1 _09806_/B sky130_fd_sc_hd__xnor2_1
Xfanout247 _06886_/A vssd1 vssd1 vccd1 vccd1 _06928_/B sky130_fd_sc_hd__buf_6
XFILLER_0_5_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout258 _07535_/B vssd1 vssd1 vccd1 vccd1 _07637_/B sky130_fd_sc_hd__clkbuf_8
Xfanout269 _06920_/B vssd1 vssd1 vccd1 vccd1 _07110_/A sky130_fd_sc_hd__buf_6
X_07996_ _07996_/A _07996_/B vssd1 vssd1 vccd1 vccd1 _08093_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07581__A2 _07541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13103__B2 _07634_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09735_ _09736_/B vssd1 vssd1 vccd1 vccd1 _09735_/Y sky130_fd_sc_hd__inv_2
X_06947_ _11126_/A _07471_/A vssd1 vssd1 vccd1 vccd1 _06947_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10468__A2 _11587_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09666_ _09443_/X _09463_/X _09703_/B vssd1 vssd1 vccd1 vccd1 _09666_/X sky130_fd_sc_hd__mux2_1
X_06878_ instruction[29] _12981_/C vssd1 vssd1 vccd1 vccd1 _13000_/B sky130_fd_sc_hd__and2_4
X_08617_ _08615_/A _08615_/B _08616_/Y vssd1 vssd1 vccd1 vccd1 _08980_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__13092__B _13129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ _09598_/A _09598_/B vssd1 vssd1 vccd1 vccd1 _09597_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_82_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09997__S _10004_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07090__B _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ _08608_/A _08548_/B vssd1 vssd1 vccd1 vccd1 _08577_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08479_ _09948_/A _08479_/B vssd1 vssd1 vccd1 vccd1 _08480_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11621__A _12417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10510_ _10510_/A _10510_/B vssd1 vssd1 vccd1 vccd1 _10511_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_80_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11490_ _12867_/S _11490_/B vssd1 vssd1 vccd1 vccd1 _11490_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10441_ _10441_/A _10441_/B vssd1 vssd1 vccd1 vccd1 _10441_/X sky130_fd_sc_hd__and2_1
XFILLER_0_17_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08046__B1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10372_ _07455_/Y _07643_/B fanout13/X wire122/X vssd1 vssd1 vccd1 vccd1 _10373_/B
+ sky130_fd_sc_hd__a22o_1
X_13160_ _07492_/Y _13196_/A2 hold74/X _13547_/A vssd1 vssd1 vccd1 vccd1 hold75/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12111_ _12111_/A _12111_/B vssd1 vssd1 vccd1 vccd1 _12112_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13091_ reg1_val[22] _13129_/B vssd1 vssd1 vccd1 vccd1 _13093_/A sky130_fd_sc_hd__or2_1
XFILLER_0_103_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12042_ _11957_/B _11957_/C _12742_/A vssd1 vssd1 vccd1 vccd1 _12043_/B sky130_fd_sc_hd__a21oi_1
Xhold290 hold290/A vssd1 vssd1 vccd1 vccd1 hold290/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09761__A _10095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12944_ _12951_/A _12940_/Y _12936_/A vssd1 vssd1 vccd1 vccd1 _12945_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_87_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07281__A _07281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12875_ _13036_/B _12876_/B vssd1 vssd1 vccd1 vccd1 _12886_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11408__A1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11408__B2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11826_ _12268_/A fanout34/X fanout32/X fanout46/X vssd1 vssd1 vccd1 vccd1 _11827_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ _11758_/A _11758_/B _11758_/C vssd1 vssd1 vccd1 vccd1 _11757_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10708_ _10552_/A _10552_/C _10552_/B vssd1 vssd1 vccd1 vccd1 _10710_/B sky130_fd_sc_hd__o21ba_1
X_11688_ reg1_val[16] _11688_/B vssd1 vssd1 vccd1 vccd1 _11688_/Y sky130_fd_sc_hd__nor2_1
X_13427_ _07358_/X _13445_/A2 hold147/X vssd1 vssd1 vccd1 vccd1 hold148/A sky130_fd_sc_hd__o21a_1
XFILLER_0_113_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10639_ _12668_/A _10639_/B vssd1 vssd1 vccd1 vccd1 _10641_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ _13660_/Q _13463_/B2 _13506_/A2 hold177/X vssd1 vssd1 vccd1 vccd1 hold178/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12309_ _12309_/A _12309_/B vssd1 vssd1 vccd1 vccd1 _12309_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13289_ _13473_/B _13474_/A _13269_/X vssd1 vssd1 vccd1 vccd1 _13479_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_121_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13177__B _13191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07850_ _07848_/A _07848_/B _07849_/Y vssd1 vssd1 vccd1 vccd1 _07963_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__11895__A1 _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06801_ reg1_val[27] _07252_/A vssd1 vssd1 vccd1 vccd1 _06801_/Y sky130_fd_sc_hd__nand2_1
X_07781_ _07780_/A _07780_/B _07782_/A vssd1 vssd1 vccd1 vccd1 _07781_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_36_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09520_ _09520_/A _09520_/B vssd1 vssd1 vccd1 vccd1 _09520_/X sky130_fd_sc_hd__or2_4
XANTENNA__07191__A _07281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09451_ _10176_/A _09449_/X _09450_/X _10457_/S vssd1 vssd1 vccd1 vccd1 _09451_/X
+ sky130_fd_sc_hd__o211a_1
X_08402_ _08402_/A _08402_/B vssd1 vssd1 vccd1 vccd1 _08403_/C sky130_fd_sc_hd__or2_1
X_09382_ _09261_/A _09261_/B _09259_/Y vssd1 vssd1 vccd1 vccd1 _09386_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_19_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08333_ _08333_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08380_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12072__A1 _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout238_A _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10083__B1 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08264_ _08857_/A _08264_/B vssd1 vssd1 vccd1 vccd1 _08309_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_74_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07130__S _07135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07215_ _07213_/A _07213_/B _07214_/Y _07521_/A vssd1 vssd1 vccd1 vccd1 _07217_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_0_116_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08195_ _07175_/X _07544_/Y _11638_/A _08933_/B vssd1 vssd1 vccd1 vccd1 _08196_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12971__S _12971_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07146_ _12971_/S _07146_/B vssd1 vssd1 vccd1 vccd1 dest_mask[0] sky130_fd_sc_hd__nand2_8
XFILLER_0_70_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09240__A2 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07077_ _07077_/A _07077_/B vssd1 vssd1 vccd1 vccd1 _07077_/X sky130_fd_sc_hd__and2_1
XFILLER_0_112_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13087__B _13129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08200__B1 _09949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07554__A2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09581__A _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07979_ _08041_/A _08041_/B _07975_/Y vssd1 vssd1 vccd1 vccd1 _07991_/B sky130_fd_sc_hd__o21a_1
X_09718_ _12537_/B2 _09692_/X _09698_/X _09717_/Y vssd1 vssd1 vccd1 vccd1 _09718_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_97_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08197__A _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990_ _11463_/A _10990_/B vssd1 vssd1 vccd1 vccd1 _10990_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09700__B1 _12795_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09649_ _09649_/A _09649_/B vssd1 vssd1 vccd1 vccd1 _09650_/B sky130_fd_sc_hd__xnor2_4
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10310__A1 _10734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _12710_/B2 _10010_/X _12656_/X _12659_/X vssd1 vssd1 vccd1 vccd1 _12660_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _11611_/A _11611_/B vssd1 vssd1 vccd1 vccd1 _11619_/A sky130_fd_sc_hd__or2_1
XFILLER_0_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08806__A2 _08806_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12591_ _12225_/A _10193_/Y _12589_/X _12590_/Y vssd1 vssd1 vccd1 vccd1 _12591_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11542_ _11542_/A _11542_/B _11542_/C vssd1 vssd1 vccd1 vccd1 _11543_/B sky130_fd_sc_hd__and3_1
XFILLER_0_107_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11473_ _09714_/X _11472_/X _11576_/A vssd1 vssd1 vccd1 vccd1 _11473_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09767__B1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13212_ hold30/X hold247/X vssd1 vssd1 vccd1 vccd1 _13313_/A sky130_fd_sc_hd__and2b_1
X_10424_ _10424_/A _10424_/B vssd1 vssd1 vccd1 vccd1 _10426_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09231__A2 _10536_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13143_ hold17/X _13207_/B vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__or2_1
X_10355_ _11076_/A _10355_/B vssd1 vssd1 vccd1 vccd1 _10359_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_20_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09782__A3 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ _13074_/A _13074_/B vssd1 vssd1 vccd1 vccd1 _13081_/C sky130_fd_sc_hd__nand2_2
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _10286_/A _10286_/B vssd1 vssd1 vccd1 vccd1 _10287_/B sky130_fd_sc_hd__xnor2_4
X_12025_ _12025_/A _12025_/B vssd1 vssd1 vccd1 vccd1 _12027_/B sky130_fd_sc_hd__xnor2_1
X_12927_ reg1_val[19] curr_PC[19] _12978_/S vssd1 vssd1 vccd1 vccd1 _12929_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_88_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12858_ _12858_/A _12858_/B _12858_/C vssd1 vssd1 vccd1 vccd1 _12859_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_75_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11809_ _12253_/A _11809_/B vssd1 vssd1 vccd1 vccd1 _11810_/A sky130_fd_sc_hd__xnor2_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12789_ reg1_val[31] _12754_/A _12788_/Y vssd1 vssd1 vccd1 vccd1 _12789_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11801__B2 _11913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07000_ reg1_val[4] _11576_/A vssd1 vssd1 vccd1 vccd1 _07000_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09758__B1 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12762__C1 _12971_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12092__A _12092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08951_ _08951_/A _08954_/B vssd1 vssd1 vccd1 vccd1 _08953_/B sky130_fd_sc_hd__xnor2_1
X_07902_ _10078_/A _07902_/B vssd1 vssd1 vccd1 vccd1 _07909_/A sky130_fd_sc_hd__xor2_2
X_08882_ _08885_/A _08885_/B vssd1 vssd1 vccd1 vccd1 _08882_/X sky130_fd_sc_hd__and2_1
XANTENNA__12820__A _12995_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07914__A _12092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09930__B1 _10542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07833_ _09161_/A _07833_/B vssd1 vssd1 vccd1 vccd1 _07994_/B sky130_fd_sc_hd__nand2_1
XANTENNA_fanout188_A _07118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07764_ fanout39/X _13149_/A _13151_/A _08118_/B vssd1 vssd1 vccd1 vccd1 _07765_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09503_ _12648_/A _09499_/Y _09502_/Y _09529_/B vssd1 vssd1 vccd1 vccd1 _09503_/X
+ sky130_fd_sc_hd__a211o_1
X_07695_ _07713_/A _07713_/B _07688_/Y vssd1 vssd1 vccd1 vccd1 _07709_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_78_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09434_ _12738_/S _09505_/B vssd1 vssd1 vccd1 vccd1 _09434_/Y sky130_fd_sc_hd__nor2_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08249__B1 _08395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09365_ _10507_/A _09365_/B vssd1 vssd1 vccd1 vccd1 _09367_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12267__A _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08316_ _09591_/A _08316_/B vssd1 vssd1 vccd1 vccd1 _08322_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09296_ _09296_/A _09296_/B vssd1 vssd1 vccd1 vccd1 _09297_/B sky130_fd_sc_hd__nor2_2
XANTENNA_30 reg1_val[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_41 reg1_val[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_52 reg2_val[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_63 reg2_val[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08247_ _10266_/A _08247_/B vssd1 vssd1 vccd1 vccd1 _08251_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_74 reg1_val[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_85 reg1_val[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09749__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08178_ _08178_/A _08178_/B _08178_/C vssd1 vssd1 vccd1 vccd1 _08288_/A sky130_fd_sc_hd__or3_1
XFILLER_0_120_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07129_ instruction[16] _07129_/B vssd1 vssd1 vccd1 vccd1 dest_idx[5] sky130_fd_sc_hd__and2_4
XFILLER_0_113_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10140_ _10140_/A _10140_/B vssd1 vssd1 vccd1 vccd1 _10142_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10071_ _10217_/B _10071_/B vssd1 vssd1 vccd1 vccd1 _10113_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_100_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07824__A _10266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08488__B1 _08580_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10973_ _10974_/B _10974_/A vssd1 vssd1 vccd1 vccd1 _11104_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__11780__S _12525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12712_ _12706_/Y _12707_/X _12711_/Y vssd1 vssd1 vccd1 vccd1 _12712_/X sky130_fd_sc_hd__o21a_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13692_ _13701_/CLK hold115/X vssd1 vssd1 vccd1 vccd1 hold113/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12643_ _12642_/A _12642_/B _12642_/Y _09507_/X vssd1 vssd1 vccd1 vccd1 _12643_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12574_ _12681_/A _12574_/B vssd1 vssd1 vccd1 vccd1 _12635_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_53_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11525_ _11525_/A _11525_/B vssd1 vssd1 vccd1 vccd1 _11533_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_80_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13500__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12339__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11456_ _11663_/A _11456_/B vssd1 vssd1 vccd1 vccd1 _11458_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_21_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07215__A1 _07213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10407_ _10407_/A _10407_/B vssd1 vssd1 vccd1 vccd1 _10410_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_max_cap153_A _07399_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11011__A2 _11793_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11387_ _11301_/A _11301_/B _11300_/A vssd1 vssd1 vccd1 vccd1 _11392_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13126_ _13126_/A _13126_/B vssd1 vssd1 vccd1 vccd1 _13128_/A sky130_fd_sc_hd__nand2_2
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10338_ _12047_/C1 _10311_/X _12525_/B _12759_/A1 _10337_/X vssd1 vssd1 vccd1 vccd1
+ _10338_/X sky130_fd_sc_hd__a221o_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _13057_/A _13057_/B _13057_/C vssd1 vssd1 vccd1 vccd1 _13058_/B sky130_fd_sc_hd__nand3_1
X_10269_ _10270_/A _10270_/B vssd1 vssd1 vccd1 vccd1 _10269_/Y sky130_fd_sc_hd__nand2_1
X_12008_ _12092_/A _12008_/B vssd1 vssd1 vccd1 vccd1 _12010_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09140__A1 _07237_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09140__B2 _08950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07480_ _09940_/A _07480_/B vssd1 vssd1 vccd1 vccd1 _07499_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12087__A _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09150_ _09150_/A _09150_/B vssd1 vssd1 vccd1 vccd1 _09151_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_56_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08101_ _08101_/A _08101_/B vssd1 vssd1 vccd1 vccd1 _08166_/B sky130_fd_sc_hd__xnor2_1
X_09081_ _09081_/A _09081_/B vssd1 vssd1 vccd1 vccd1 _09082_/C sky130_fd_sc_hd__xor2_2
XFILLER_0_44_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08032_ _08030_/A _08030_/B _08031_/Y vssd1 vssd1 vccd1 vccd1 _08104_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_4_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout103_A _07299_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09983_ _09985_/A _09985_/B vssd1 vssd1 vccd1 vccd1 _09983_/X sky130_fd_sc_hd__or2_2
XANTENNA__10761__A1 _11866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08934_ _09948_/A _08944_/B _08933_/X vssd1 vssd1 vccd1 vccd1 _08938_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__12550__A _12551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08865_ _08879_/A _08879_/B vssd1 vssd1 vccd1 vccd1 _08865_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08182__A2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07816_ _07813_/A _07813_/C _07813_/B vssd1 vssd1 vccd1 vccd1 _07817_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__07363__B _07363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08796_ _09501_/A wire122/A _10637_/A _08271_/A vssd1 vssd1 vccd1 vccd1 _08797_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07747_ _07747_/A _07747_/B vssd1 vssd1 vccd1 vccd1 _07776_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_79_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12266__A1 _07257_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12266__B2 _12496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09131__A1 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09131__B2 _08486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07678_ fanout28/X _07491_/X _09885_/B1 _08395_/B vssd1 vssd1 vccd1 vccd1 _07679_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07142__B1 _07110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09417_ _09417_/A _09417_/B vssd1 vssd1 vccd1 vccd1 _09419_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_90_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10029__B1 _12533_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09348_ _09347_/B _09348_/B vssd1 vssd1 vccd1 vccd1 _09349_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_75_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout16_A _07643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09279_ _09279_/A _09279_/B vssd1 vssd1 vccd1 vccd1 _09295_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11310_ _11310_/A _11310_/B vssd1 vssd1 vccd1 vccd1 _11311_/C sky130_fd_sc_hd__xnor2_1
X_12290_ _12290_/A _12290_/B vssd1 vssd1 vccd1 vccd1 _12293_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11241_ _10020_/X _11240_/Y _11576_/A vssd1 vssd1 vccd1 vccd1 _11241_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12163__C _12163_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11172_ _11172_/A _11172_/B vssd1 vssd1 vccd1 vccd1 _11174_/B sky130_fd_sc_hd__or2_1
XFILLER_0_101_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10123_ _09955_/A _10518_/A _09961_/B _09959_/X vssd1 vssd1 vccd1 vccd1 _10125_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_101_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10054_ fanout14/X _07472_/Y _07477_/X _07833_/B vssd1 vssd1 vccd1 vccd1 _10055_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10504__A1 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11701__B1 _12825_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10504__B2 _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09370__A1 _07238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11076__A _11076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09370__B2 _07239_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13454__B1 _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09122__A1 _07198_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09122__B2 _07203_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11804__A _11920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13744_ _13744_/A vssd1 vssd1 vccd1 vccd1 loadstore_size[1] sky130_fd_sc_hd__buf_12
XFILLER_0_58_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10956_ _10956_/A _10956_/B vssd1 vssd1 vccd1 vccd1 _10958_/B sky130_fd_sc_hd__xor2_1
XANTENNA__08385__A _08746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11480__A2 _12799_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13675_ _13684_/CLK _13675_/D vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__dfxtp_1
X_10887_ hold253/A _12058_/A _11007_/B _12748_/B1 vssd1 vssd1 vccd1 vccd1 _10888_/B
+ sky130_fd_sc_hd__a31o_1
X_12626_ _12626_/A _12626_/B vssd1 vssd1 vccd1 vccd1 _12728_/A sky130_fd_sc_hd__or2_2
XFILLER_0_81_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12557_ _12557_/A _12557_/B _12666_/A _12557_/D vssd1 vssd1 vccd1 vccd1 _12558_/B
+ sky130_fd_sc_hd__or4_1
XANTENNA__09928__B _12614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07729__A _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11508_ _11508_/A _11508_/B vssd1 vssd1 vccd1 vccd1 _11510_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11783__A3 _12235_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12488_ _12488_/A _12488_/B vssd1 vssd1 vccd1 vccd1 _12489_/B sky130_fd_sc_hd__and2_1
XANTENNA__11896__D _12163_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold108 hold108/A vssd1 vssd1 vccd1 vccd1 hold108/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold119 hold119/A vssd1 vssd1 vccd1 vccd1 hold119/X sky130_fd_sc_hd__dlygate4sd3_1
X_11439_ _11542_/B _11439_/B vssd1 vssd1 vccd1 vccd1 _11441_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_123_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07739__A2 _10235_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ reg1_val[26] _13136_/A vssd1 vssd1 vccd1 vccd1 _13111_/A sky130_fd_sc_hd__or2_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06980_ reg2_val[6] _06980_/B vssd1 vssd1 vccd1 vccd1 _06980_/X sky130_fd_sc_hd__and2_1
XFILLER_0_95_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07464__A _11281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13185__B _13191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08650_ _08650_/A _08650_/B vssd1 vssd1 vccd1 vccd1 _08660_/B sky130_fd_sc_hd__xnor2_2
X_07601_ _07601_/A _07601_/B vssd1 vssd1 vccd1 vccd1 _07603_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12248__A1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08581_ _09591_/A _08581_/B vssd1 vssd1 vccd1 vccd1 _08644_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12248__B2 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07532_ _07572_/S _07531_/Y _07530_/Y vssd1 vssd1 vccd1 vccd1 _07532_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__12799__A2 _12799_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07675__A1 _07366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07463_ reg1_val[16] _07462_/Y _07865_/B vssd1 vssd1 vccd1 vccd1 _07467_/B sky130_fd_sc_hd__mux2_2
XANTENNA__07675__B2 _07557_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09202_ _09203_/A _09203_/B vssd1 vssd1 vccd1 vccd1 _09202_/X sky130_fd_sc_hd__and2_1
XFILLER_0_8_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07394_ _07395_/A _07395_/B _07395_/C _07395_/D vssd1 vssd1 vccd1 vccd1 _12485_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09133_ _07300_/Y _07541_/X _07545_/Y wire101/A vssd1 vssd1 vccd1 vccd1 _09134_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08624__B1 _08868_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout220_A _07363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09064_ _09068_/A _09065_/B vssd1 vssd1 vccd1 vccd1 _12131_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07639__A _12417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12708__C1 _12799_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08015_ _08095_/A vssd1 vssd1 vccd1 vccd1 _08015_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12184__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09966_ _09966_/A _09966_/B vssd1 vssd1 vccd1 vccd1 _09967_/B sky130_fd_sc_hd__nor2_1
X_08917_ _08910_/B _08910_/C _08910_/A vssd1 vssd1 vccd1 vccd1 _08920_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__06953__A3 _13036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09897_ _09897_/A _09897_/B vssd1 vssd1 vccd1 vccd1 _09898_/B sky130_fd_sc_hd__nor2_2
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09352__A1 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09352__B2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08848_ _08849_/A _08849_/B vssd1 vssd1 vccd1 vccd1 _08861_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10004__S _10004_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08779_ _09671_/S _08778_/B _08746_/A vssd1 vssd1 vccd1 vccd1 _08781_/C sky130_fd_sc_hd__o21bai_1
XANTENNA__12239__B2 _12537_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13436__B1 _13444_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09104__A1 fanout39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09104__B2 _08118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10810_ wire122/X _11802_/B vssd1 vssd1 vccd1 vccd1 _10811_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_95_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11624__A _11731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11790_ _12760_/A1 _11780_/X _11784_/X _11789_/X vssd1 vssd1 vccd1 vccd1 _11790_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10741_ _10739_/Y _10741_/B vssd1 vssd1 vccd1 vccd1 _10742_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_67_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13460_ _13277_/X _13460_/B vssd1 vssd1 vccd1 vccd1 _13461_/B sky130_fd_sc_hd__nand2b_1
X_10672_ _11281_/A _10672_/B vssd1 vssd1 vccd1 vccd1 _10676_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08933__A _09161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07418__A1 _10456_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12411_ _12411_/A _12411_/B vssd1 vssd1 vccd1 vccd1 _12412_/B sky130_fd_sc_hd__or2_1
XFILLER_0_35_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09748__B _10518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13391_ _07172_/B _13419_/A2 hold129/X vssd1 vssd1 vccd1 vccd1 _13677_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12342_ _12417_/A _12342_/B vssd1 vssd1 vccd1 vccd1 _12344_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12273_ _12351_/B _12273_/B vssd1 vssd1 vccd1 vccd1 _12276_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12175__B1 _09145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08918__A1 _09703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08918__B2 _07399_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11224_ _10977_/A _11103_/X _11105_/B vssd1 vssd1 vccd1 vccd1 _11224_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_31_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11155_ fanout84/X _07891_/X fanout10/X _07524_/Y vssd1 vssd1 vccd1 vccd1 _11156_/B
+ sky130_fd_sc_hd__o22a_1
X_10106_ _10349_/A1 fanout9/X fanout4/X _10225_/A vssd1 vssd1 vccd1 vccd1 _10107_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11086_ _10959_/A _10959_/B _10940_/Y vssd1 vssd1 vccd1 vccd1 _11097_/A sky130_fd_sc_hd__o21a_1
XANTENNA__08146__A2 _08580_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10037_ _10028_/Y _10029_/X _10036_/X vssd1 vssd1 vccd1 vccd1 _10037_/Y sky130_fd_sc_hd__o21ai_1
X_11988_ _11988_/A _12164_/A vssd1 vssd1 vccd1 vccd1 _11988_/X sky130_fd_sc_hd__or2_1
XANTENNA__11989__B1 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13727_ _13731_/CLK _13727_/D vssd1 vssd1 vccd1 vccd1 hold255/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08854__B1 _08868_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10939_ _10939_/A _10939_/B vssd1 vssd1 vccd1 vccd1 _10941_/B sky130_fd_sc_hd__xor2_2
XANTENNA__10661__B1 _11423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13658_ _13659_/CLK hold202/X vssd1 vssd1 vccd1 vccd1 hold200/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ _09145_/Y fanout8/X fanout3/X _12667_/A vssd1 vssd1 vccd1 vccd1 _12610_/B
+ sky130_fd_sc_hd__a22o_1
X_13589_ hold172/A _13589_/B vssd1 vssd1 vccd1 vccd1 _13589_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09820_ _09821_/A _09821_/B vssd1 vssd1 vccd1 vccd1 _09820_/X sky130_fd_sc_hd__and2_1
XANTENNA__11709__A _11709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07194__A _07201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09751_ _09751_/A vssd1 vssd1 vccd1 vccd1 _09753_/C sky130_fd_sc_hd__inv_2
X_06963_ reg1_val[9] _10889_/A vssd1 vssd1 vccd1 vccd1 _06963_/Y sky130_fd_sc_hd__nor2_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09334__A1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08702_ _08873_/B2 _10538_/A _08778_/B _13149_/A vssd1 vssd1 vccd1 vccd1 _08703_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09334__B2 _07833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09682_ _09475_/X _09477_/X _09688_/S vssd1 vssd1 vccd1 vccd1 _09682_/X sky130_fd_sc_hd__mux2_1
X_06894_ instruction[27] _06894_/B vssd1 vssd1 vccd1 vccd1 _12990_/B sky130_fd_sc_hd__and2_4
XANTENNA__09885__A2 _07451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11141__B2 _11137_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08633_ _09659_/B _08633_/B vssd1 vssd1 vccd1 vccd1 _08637_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__13418__B1 _13444_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout170_A _12759_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout268_A _07110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ _08573_/A _08563_/Y _08519_/Y vssd1 vssd1 vccd1 vccd1 _08571_/A sky130_fd_sc_hd__o21a_2
XANTENNA__07133__S _07135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07515_ reg1_val[14] _07865_/B vssd1 vssd1 vccd1 vccd1 _07517_/D sky130_fd_sc_hd__nor2_1
X_08495_ _08495_/A _08495_/B vssd1 vssd1 vccd1 vccd1 _08556_/B sky130_fd_sc_hd__xnor2_1
Xfanout14 _07417_/X vssd1 vssd1 vccd1 vccd1 fanout14/X sky130_fd_sc_hd__clkbuf_8
Xfanout25 _07468_/X vssd1 vssd1 vccd1 vccd1 fanout25/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout36 _08118_/B vssd1 vssd1 vccd1 vccd1 fanout36/X sky130_fd_sc_hd__clkbuf_8
Xfanout47 _07229_/X vssd1 vssd1 vccd1 vccd1 fanout47/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07446_ _11913_/A _07453_/B vssd1 vssd1 vccd1 vccd1 _07446_/Y sky130_fd_sc_hd__nor2_1
Xfanout58 _10522_/B vssd1 vssd1 vccd1 vccd1 _12666_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout69 _07576_/Y vssd1 vssd1 vccd1 vccd1 _10538_/A sky130_fd_sc_hd__buf_6
XFILLER_0_9_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07377_ _07377_/A _07377_/B _07377_/C vssd1 vssd1 vccd1 vccd1 _07386_/A sky130_fd_sc_hd__and3_1
X_09116_ _09116_/A _09116_/B vssd1 vssd1 vccd1 vccd1 _09186_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__10404__B1 _07526_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09047_ _09047_/A _09047_/B vssd1 vssd1 vccd1 vccd1 _11672_/A sky130_fd_sc_hd__or2_1
XANTENNA__07088__B _13748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_368 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout83_A fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09949_ _09949_/A _09950_/B vssd1 vssd1 vccd1 vccd1 _09949_/Y sky130_fd_sc_hd__nand2_1
X_12960_ _12979_/A _12960_/B vssd1 vssd1 vccd1 vccd1 _12964_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__11132__B2 _12648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07832__A _10119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11911_ _12253_/A _11911_/B vssd1 vssd1 vccd1 vccd1 _11913_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07887__A1 _08821_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07887__B2 _08821_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12891_ _12900_/A _12891_/B vssd1 vssd1 vccd1 vccd1 _12893_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_87_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10891__B1 _12754_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11842_ _11746_/A _11746_/B _11744_/X vssd1 vssd1 vccd1 vccd1 _11843_/B sky130_fd_sc_hd__a21oi_2
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _12515_/S _11771_/X _11772_/X vssd1 vssd1 vccd1 vccd1 _11774_/B sky130_fd_sc_hd__a21oi_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13512_ _13543_/A hold290/X vssd1 vssd1 vccd1 vccd1 _13718_/D sky130_fd_sc_hd__and2_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09759__A _11076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10724_ _10724_/A _10981_/C vssd1 vssd1 vccd1 vccd1 _11151_/A sky130_fd_sc_hd__xor2_4
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13443_ _09160_/B _13445_/A2 hold33/X vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__o21a_1
XANTENNA__13188__A2 _13196_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10655_ _10656_/A _10656_/B vssd1 vssd1 vccd1 vccd1 _10783_/B sky130_fd_sc_hd__and2_1
XANTENNA__12185__A _12764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12396__B1 _12657_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13374_ _13668_/Q _13599_/D _13584_/B hold219/X vssd1 vssd1 vccd1 vccd1 hold220/A
+ sky130_fd_sc_hd__a22o_1
X_10586_ _11562_/A _09018_/A _09018_/B vssd1 vssd1 vccd1 vccd1 _10586_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12325_ curr_PC[22] curr_PC[23] _12325_/C vssd1 vssd1 vccd1 vccd1 _12477_/C sky130_fd_sc_hd__and3_1
XFILLER_0_106_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12256_ _12334_/B _12256_/B vssd1 vssd1 vccd1 vccd1 _12258_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_31_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11207_ _11066_/A _11065_/B _11065_/A vssd1 vssd1 vccd1 vccd1 _11209_/C sky130_fd_sc_hd__o21ba_1
XFILLER_0_76_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13360__A2 _13463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12187_ _12187_/A _12187_/B _12187_/C vssd1 vssd1 vccd1 vccd1 _12188_/B sky130_fd_sc_hd__and3_1
X_11138_ _11138_/A _11586_/B vssd1 vssd1 vccd1 vccd1 _11138_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08119__A2 _07300_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13744__A _13744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11069_ _11069_/A _11069_/B vssd1 vssd1 vccd1 vccd1 _11085_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_25_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07300_ _07300_/A _07300_/B vssd1 vssd1 vccd1 vccd1 _07300_/Y sky130_fd_sc_hd__xnor2_4
X_08280_ _08350_/A _08350_/B _08350_/C vssd1 vssd1 vccd1 vccd1 _08351_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07231_ _12982_/A _09694_/A reg1_val[2] vssd1 vssd1 vccd1 vccd1 _09871_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07162_ _07535_/B _07160_/Y _07161_/X vssd1 vssd1 vccd1 vccd1 _10240_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__09252__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07093_ _07093_/A _07093_/B vssd1 vssd1 vccd1 vccd1 _07095_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_41_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07917__A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout204 _07151_/X vssd1 vssd1 vccd1 vccd1 _12799_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout215 _10456_/S vssd1 vssd1 vccd1 vccd1 _10600_/S sky130_fd_sc_hd__clkbuf_8
Xfanout226 _06789_/Y vssd1 vssd1 vccd1 vccd1 _06906_/B1 sky130_fd_sc_hd__clkbuf_4
X_09803_ _09804_/B _09804_/A vssd1 vssd1 vccd1 vccd1 _09803_/X sky130_fd_sc_hd__and2b_1
Xfanout237 _12867_/S vssd1 vssd1 vccd1 vccd1 _12825_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout248 _13142_/A vssd1 vssd1 vccd1 vccd1 _13416_/A2 sky130_fd_sc_hd__buf_4
X_07995_ _07997_/A _07997_/B vssd1 vssd1 vccd1 vccd1 _07995_/X sky130_fd_sc_hd__or2_1
Xfanout259 _07156_/Y vssd1 vssd1 vccd1 vccd1 _07535_/B sky130_fd_sc_hd__buf_6
X_09734_ _09734_/A _09734_/B vssd1 vssd1 vccd1 vccd1 _09736_/B sky130_fd_sc_hd__xnor2_4
X_06946_ _06928_/A _06936_/B _13042_/B _06944_/X vssd1 vssd1 vccd1 vccd1 _07471_/A
+ sky130_fd_sc_hd__a31oi_4
X_09665_ _09663_/X _09664_/X _10004_/S vssd1 vssd1 vccd1 vccd1 _09665_/X sky130_fd_sc_hd__mux2_1
X_06877_ _12303_/A _12218_/A _12046_/A _12136_/A vssd1 vssd1 vccd1 vccd1 _07099_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_96_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08616_ _08655_/B _08655_/A vssd1 vssd1 vccd1 vccd1 _08616_/Y sky130_fd_sc_hd__nand2b_1
X_09596_ _10507_/A _09596_/B vssd1 vssd1 vccd1 vccd1 _09598_/B sky130_fd_sc_hd__xnor2_2
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ _08608_/A _08548_/B vssd1 vssd1 vccd1 vccd1 _08547_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_77_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08478_ _08933_/B _07478_/A _07478_/B _13168_/A1 _07175_/X vssd1 vssd1 vccd1 vccd1
+ _08479_/B sky130_fd_sc_hd__a32o_1
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12717__B fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07429_ _07429_/A vssd1 vssd1 vccd1 vccd1 _07486_/A sky130_fd_sc_hd__inv_2
XFILLER_0_64_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10518__A _10518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12378__B1 _10866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08046__A1 _10235_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10440_ _09830_/B _10435_/C _10438_/Y _10981_/A vssd1 vssd1 vccd1 vccd1 _10441_/B
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__08046__B2 _10235_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10371_ _10371_/A _10371_/B vssd1 vssd1 vccd1 vccd1 _10382_/A sky130_fd_sc_hd__xnor2_2
X_12110_ _12110_/A _12110_/B _12110_/C vssd1 vssd1 vccd1 vccd1 _12111_/B sky130_fd_sc_hd__or3_1
XANTENNA__07827__A _10263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13090_ _13102_/B _13090_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[21] sky130_fd_sc_hd__xor2_4
XFILLER_0_103_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12041_ _12695_/A _11988_/X _12164_/B _11955_/A vssd1 vssd1 vccd1 vccd1 _12041_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__13342__A2 _13506_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold280 hold280/A vssd1 vssd1 vccd1 vccd1 hold280/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold291 hold291/A vssd1 vssd1 vccd1 vccd1 hold291/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06897__A2_N _06980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07562__A _10263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12943_ _12956_/A _12943_/B vssd1 vssd1 vccd1 vccd1 _12951_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_99_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12874_ _11126_/A curr_PC[11] _12978_/S vssd1 vssd1 vccd1 vccd1 _12876_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_68_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11825_ _11825_/A _11825_/B vssd1 vssd1 vccd1 vccd1 _11829_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12605__A1 _10866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11408__A2 _07891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11812__A _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09482__A0 _09501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _11756_/A _11756_/B vssd1 vssd1 vccd1 vccd1 _11758_/C sky130_fd_sc_hd__xor2_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10707_ _10511_/A _10511_/B _10513_/B _10516_/A vssd1 vssd1 vccd1 vccd1 _10710_/A
+ sky130_fd_sc_hd__a31oi_2
XFILLER_0_71_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11687_ hold292/A _11685_/X _11686_/Y vssd1 vssd1 vccd1 vccd1 _11696_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13426_ _13694_/Q _13142_/A _13444_/B1 hold146/X _13430_/C1 vssd1 vssd1 vccd1 vccd1
+ hold147/A sky130_fd_sc_hd__o221a_1
XFILLER_0_70_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10638_ _07477_/X fanout16/X fanout12/X _07472_/Y vssd1 vssd1 vccd1 vccd1 _10639_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13357_ _13359_/A hold186/X vssd1 vssd1 vccd1 vccd1 hold187/A sky130_fd_sc_hd__and2_1
X_10569_ _10569_/A _10569_/B vssd1 vssd1 vccd1 vccd1 _10571_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_51_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12308_ _12224_/A _12224_/B _12222_/B vssd1 vssd1 vccd1 vccd1 _12309_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_23_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13288_ _13273_/B _13469_/B _13271_/X vssd1 vssd1 vccd1 vccd1 _13474_/A sky130_fd_sc_hd__a21o_1
X_12239_ _12218_/A _12793_/A2 _10895_/Y _12537_/B2 _12238_/Y vssd1 vssd1 vccd1 vccd1
+ _12239_/X sky130_fd_sc_hd__a221o_1
XANTENNA__07012__A2 _06936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06800_ reg1_val[27] _07252_/A vssd1 vssd1 vccd1 vccd1 _06802_/B sky130_fd_sc_hd__and2_1
X_07780_ _07780_/A _07780_/B vssd1 vssd1 vccd1 vccd1 _07782_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_36_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13193__B _13193_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09450_ _10004_/S _09442_/X _09439_/X _10456_/S vssd1 vssd1 vccd1 vccd1 _09450_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08401_ _08401_/A _08401_/B vssd1 vssd1 vccd1 vccd1 _08402_/B sky130_fd_sc_hd__and2_1
X_09381_ _09381_/A _10522_/B vssd1 vssd1 vccd1 vccd1 _09387_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_47_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08332_ _09371_/A _08332_/B vssd1 vssd1 vccd1 vccd1 _08380_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09399__A _10119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10607__B1 _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10083__A1 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08263_ _08806_/A2 _13166_/A1 _13168_/A1 _08806_/B1 vssd1 vssd1 vccd1 vccd1 _08264_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10083__B2 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11280__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07214_ _07252_/B _07252_/D vssd1 vssd1 vccd1 vccd1 _07214_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_116_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08194_ _08255_/A _08255_/B vssd1 vssd1 vccd1 vccd1 _08256_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07145_ instruction[24] _12578_/A is_load _06989_/B _07144_/X vssd1 vssd1 vccd1 vccd1
+ _07146_/B sky130_fd_sc_hd__a32o_2
XANTENNA__13572__A2 _13584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07076_ _07059_/A _07059_/B _12382_/A vssd1 vssd1 vccd1 vccd1 _07077_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_112_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13324__A2 _13463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11169__A _12253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10073__A _11076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07539__B1 _11076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07978_ _07978_/A _07978_/B vssd1 vssd1 vccd1 vccd1 _08041_/B sky130_fd_sc_hd__xnor2_2
X_09717_ _09699_/Y _09700_/X _09716_/A _09839_/A _09711_/X vssd1 vssd1 vccd1 vccd1
+ _09717_/Y sky130_fd_sc_hd__o221ai_1
X_06929_ reg2_val[13] _06980_/B _06928_/X vssd1 vssd1 vccd1 vccd1 _07522_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_69_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09648_ _09648_/A _09648_/B vssd1 vssd1 vccd1 vccd1 _09649_/B sky130_fd_sc_hd__xor2_4
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _09579_/A _09579_/B vssd1 vssd1 vccd1 vccd1 _09602_/A sky130_fd_sc_hd__xnor2_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12599__B1 _09519_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11610_ _11610_/A _11610_/B _11610_/C vssd1 vssd1 vccd1 vccd1 _11611_/B sky130_fd_sc_hd__and3_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12590_ _12589_/A _12589_/B _12225_/A vssd1 vssd1 vccd1 vccd1 _12590_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10893__D _10893_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11541_ _11542_/A _11542_/B _11542_/C vssd1 vssd1 vccd1 vccd1 _11543_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10248__A _11076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09216__B1 _07699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11472_ _10454_/X _10456_/X _11472_/S vssd1 vssd1 vccd1 vccd1 _11472_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_33_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13211_ _13211_/A _13211_/B vssd1 vssd1 vccd1 vccd1 _13585_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09767__A1 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10423_ _10287_/A _10287_/B _10285_/Y vssd1 vssd1 vccd1 vccd1 _10424_/B sky130_fd_sc_hd__a21boi_4
XANTENNA__09767__B2 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13563__A2 _13584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13142_ _13142_/A _13142_/B vssd1 vssd1 vccd1 vccd1 _13142_/Y sky130_fd_sc_hd__nand2_1
X_10354_ _07577_/X _10787_/B _10787_/C _10538_/A fanout44/X vssd1 vssd1 vccd1 vccd1
+ _10355_/B sky130_fd_sc_hd__o32a_2
XFILLER_0_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13073_ reg1_val[18] _13129_/B vssd1 vssd1 vccd1 vccd1 _13074_/B sky130_fd_sc_hd__nand2_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10285_ _10124_/X _10128_/A _10286_/A vssd1 vssd1 vccd1 vccd1 _10285_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09772__A _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12024_ _12024_/A _12024_/B vssd1 vssd1 vccd1 vccd1 _12025_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08388__A _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07292__A _13015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12926_ _12931_/B _12926_/B vssd1 vssd1 vccd1 vccd1 new_PC[18] sky130_fd_sc_hd__and2_4
XANTENNA__07702__B1 _07833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12857_ _12858_/A _12858_/B _12858_/C vssd1 vssd1 vccd1 vccd1 _12865_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_29_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08835__B _08862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11808_ _12557_/B fanout38/X fanout36/X _07597_/X vssd1 vssd1 vccd1 vccd1 _11809_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_29_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12788_ reg1_val[31] _12754_/A _12598_/C vssd1 vssd1 vccd1 vccd1 _12788_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire101_A wire101/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11739_ _11739_/A _11739_/B vssd1 vssd1 vccd1 vccd1 _11753_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11801__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08851__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09758__A1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09758__B2 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13409_ _10507_/A _13419_/A2 hold93/X vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__o21a_1
XFILLER_0_98_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07467__A _11508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07233__A2 _07535_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08950_ _09671_/S _08950_/B vssd1 vssd1 vccd1 vccd1 _08954_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_20_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07901_ fanout40/X _07307_/Y _08833_/B fanout56/X vssd1 vssd1 vccd1 vccd1 _07902_/B
+ sky130_fd_sc_hd__o22a_1
X_08881_ _08881_/A _08881_/B vssd1 vssd1 vccd1 vccd1 _08885_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07832_ _10119_/A _07832_/B vssd1 vssd1 vccd1 vccd1 _07994_/A sky130_fd_sc_hd__xnor2_2
X_07763_ _09779_/A _07763_/B vssd1 vssd1 vccd1 vccd1 _07970_/B sky130_fd_sc_hd__xnor2_1
X_09502_ _09696_/A _09501_/X _12648_/A vssd1 vssd1 vccd1 vccd1 _09502_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07694_ _10050_/A _07694_/B vssd1 vssd1 vccd1 vccd1 _07713_/B sky130_fd_sc_hd__xnor2_2
X_09433_ instruction[3] _13748_/A _09520_/B _07086_/Y vssd1 vssd1 vccd1 vccd1 _09433_/X
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_63_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout250_A _13463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11452__A _11452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09364_ fanout42/X fanout75/X _08704_/B fanout40/X vssd1 vssd1 vccd1 vccd1 _09365_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08249__A1 _13147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08249__B2 _13149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08315_ _08866_/A2 fanout84/X _08580_/B _09216_/B2 vssd1 vssd1 vccd1 vccd1 _08316_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_117_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09295_ _09295_/A _09295_/B vssd1 vssd1 vccd1 vccd1 _09296_/B sky130_fd_sc_hd__nor2_1
XANTENNA_20 instruction[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_31 reg1_val[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_42 reg1_val[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08246_ _09671_/S _08246_/B vssd1 vssd1 vccd1 vccd1 _08247_/B sky130_fd_sc_hd__nor2_1
XANTENNA_53 reg2_val[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_64 reg2_val[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_75 reg1_val[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_86 reg1_val[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09749__A1 _10104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09749__B2 _09955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08177_ _08177_/A _08177_/B vssd1 vssd1 vccd1 vccd1 _08178_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_30_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07128_ instruction[15] _07129_/B vssd1 vssd1 vccd1 vccd1 dest_idx[4] sky130_fd_sc_hd__and2_4
XFILLER_0_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10007__S _10007_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07059_ _07059_/A _07059_/B vssd1 vssd1 vccd1 vccd1 _07059_/X sky130_fd_sc_hd__and2_1
XFILLER_0_112_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10070_ _10070_/A _10070_/B vssd1 vssd1 vccd1 vccd1 _10071_/B sky130_fd_sc_hd__or2_1
XANTENNA__07932__B1 _11638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap11 _09145_/Y vssd1 vssd1 vccd1 vccd1 _10536_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08488__A1 _08873_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10972_ _10972_/A _10972_/B vssd1 vssd1 vccd1 vccd1 _10974_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08488__B2 _13149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap55 _07203_/Y vssd1 vssd1 vccd1 vccd1 _12189_/A sky130_fd_sc_hd__buf_4
XFILLER_0_69_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12711_ _07866_/X _12754_/C _12710_/X vssd1 vssd1 vccd1 vccd1 _12711_/Y sky130_fd_sc_hd__a21oi_1
X_13691_ _13701_/CLK hold153/X vssd1 vssd1 vccd1 vccd1 hold151/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09437__A0 _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12642_ _12642_/A _12642_/B vssd1 vssd1 vccd1 vccd1 _12642_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12177__B fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09988__A1 _09824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12573_ _12295_/B _12440_/C _12682_/C _12572_/X vssd1 vssd1 vccd1 vccd1 _12574_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07999__B1 _08868_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11524_ _11524_/A _11524_/B vssd1 vssd1 vccd1 vccd1 _11525_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_53_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11455_ _10984_/B _11454_/Y _11453_/X vssd1 vssd1 vccd1 vccd1 _11456_/B sky130_fd_sc_hd__o21ba_1
XANTENNA__06903__B _12981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10406_ _10407_/A _10407_/B vssd1 vssd1 vccd1 vccd1 _10515_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_68_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11386_ _11332_/A _11332_/B _11330_/Y vssd1 vssd1 vccd1 vccd1 _11447_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_21_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13125_ reg1_val[29] _13136_/A vssd1 vssd1 vccd1 vccd1 _13126_/B sky130_fd_sc_hd__or2_1
XFILLER_0_21_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10337_ _10320_/X _10321_/X _10323_/Y _09523_/Y _10336_/X vssd1 vssd1 vccd1 vccd1
+ _10337_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_103_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _13057_/A _13057_/B _13057_/C vssd1 vssd1 vccd1 vccd1 _13061_/B sky130_fd_sc_hd__a21o_1
X_10268_ _11709_/A _10268_/B vssd1 vssd1 vccd1 vccd1 _10270_/B sky130_fd_sc_hd__xnor2_1
X_12007_ _07257_/X fanout15/X fanout31/X _12614_/A vssd1 vssd1 vccd1 vccd1 _12008_/B
+ sky130_fd_sc_hd__a22o_1
X_10199_ _10197_/X _10198_/X _10342_/A vssd1 vssd1 vccd1 vccd1 dest_val[4] sky130_fd_sc_hd__mux2_8
XFILLER_0_108_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09140__A2 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12909_ reg1_val[16] curr_PC[16] _12978_/S vssd1 vssd1 vccd1 vccd1 _12910_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11272__A _11514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12087__B _12666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10038__A1 _12047_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08100_ _08098_/A _08098_/B _08099_/Y vssd1 vssd1 vccd1 vccd1 _08166_/A sky130_fd_sc_hd__o21ai_1
X_09080_ _09080_/A _09080_/B _09080_/C vssd1 vssd1 vccd1 vccd1 _09081_/B sky130_fd_sc_hd__and3_1
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08581__A _09591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08031_ _08038_/B _08038_/A vssd1 vssd1 vccd1 vccd1 _08031_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_71_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12534__C _12754_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12735__B1 _09429_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09982_ _09982_/A _09982_/B vssd1 vssd1 vccd1 vccd1 _09985_/B sky130_fd_sc_hd__xnor2_4
X_08933_ _09161_/A _08933_/B _08944_/A vssd1 vssd1 vccd1 vccd1 _08933_/X sky130_fd_sc_hd__and3_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08864_ _08864_/A _08864_/B vssd1 vssd1 vccd1 vccd1 _08879_/B sky130_fd_sc_hd__xor2_2
X_07815_ _07815_/A _07815_/B vssd1 vssd1 vccd1 vccd1 _07817_/B sky130_fd_sc_hd__nand2_1
X_08795_ _09373_/A _08795_/B vssd1 vssd1 vccd1 vccd1 _08799_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07746_ _07843_/A _07843_/B vssd1 vssd1 vccd1 vccd1 _07747_/B sky130_fd_sc_hd__and2b_1
XANTENNA__12266__A2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13463__B2 _13463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09131__A2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07677_ _07680_/A _07680_/B vssd1 vssd1 vccd1 vccd1 _07683_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_66_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09416_ _09416_/A _09416_/B vssd1 vssd1 vccd1 vccd1 _09417_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_75_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09347_ _09348_/B _09347_/B vssd1 vssd1 vccd1 vccd1 _09559_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__11226__B1 _11224_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09278_ _09278_/A _09278_/B vssd1 vssd1 vccd1 vccd1 _09279_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08491__A _08746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08229_ _08229_/A _08229_/B vssd1 vssd1 vccd1 vccd1 _08240_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_90_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12217__S _12578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11240_ _11240_/A vssd1 vssd1 vccd1 vccd1 _11240_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_30_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10737__C1 _12047_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11171_ _11171_/A _11171_/B vssd1 vssd1 vccd1 vccd1 _11172_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_113_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10122_ _10253_/A _10122_/B vssd1 vssd1 vccd1 vccd1 _10125_/A sky130_fd_sc_hd__and2_1
XFILLER_0_101_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10053_ _11731_/A _10053_/B vssd1 vssd1 vccd1 vccd1 _10057_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07905__B1 _10235_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10504__A2 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09370__A2 _12667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08666__A _09659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09122__A2 _10536_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13743_ instruction[5] vssd1 vssd1 vccd1 vccd1 loadstore_size[0] sky130_fd_sc_hd__buf_12
X_10955_ _10956_/A _10956_/B vssd1 vssd1 vccd1 vccd1 _11087_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_58_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13206__A1 _09145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13674_ _13684_/CLK hold2/X vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
X_10886_ _11252_/B _11007_/B hold253/A vssd1 vssd1 vccd1 vccd1 _10888_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12625_ _12625_/A _12625_/B _12625_/C vssd1 vssd1 vccd1 vccd1 _12626_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_26_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12556_ _12557_/A _12557_/D _12557_/B vssd1 vssd1 vccd1 vccd1 _12558_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11507_ _11507_/A _11507_/B vssd1 vssd1 vccd1 vccd1 _11508_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_123_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12487_ _12488_/A _12488_/B vssd1 vssd1 vccd1 vccd1 _12560_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold109 hold109/A vssd1 vssd1 vccd1 vccd1 hold109/X sky130_fd_sc_hd__dlygate4sd3_1
X_11438_ _11438_/A _11438_/B _11438_/C vssd1 vssd1 vccd1 vccd1 _11439_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_21_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11369_ hold271/A _11369_/B vssd1 vssd1 vccd1 vccd1 _11579_/C sky130_fd_sc_hd__or2_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ _13108_/A _13112_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[25] sky130_fd_sc_hd__xnor2_4
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13039_ _13039_/A _13039_/B _13039_/C vssd1 vssd1 vccd1 vccd1 _13040_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07600_ _07601_/A _07601_/B vssd1 vssd1 vccd1 vccd1 _07874_/A sky130_fd_sc_hd__nand2_1
X_08580_ _09674_/S _08580_/B vssd1 vssd1 vccd1 vccd1 _08581_/B sky130_fd_sc_hd__nor2_1
XANTENNA__13445__A1 _12764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12248__A2 _09145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07480__A _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07531_ _07531_/A _07571_/A vssd1 vssd1 vccd1 vccd1 _07531_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_88_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06808__B _12981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07462_ reg1_val[16] _07462_/B vssd1 vssd1 vccd1 vccd1 _07462_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__07675__A2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09201_ _09203_/A _09203_/B vssd1 vssd1 vccd1 vccd1 _09201_/X sky130_fd_sc_hd__or2_1
XFILLER_0_119_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07393_ _07395_/C _07395_/D vssd1 vssd1 vccd1 vccd1 _07393_/X sky130_fd_sc_hd__and2_1
XANTENNA__12826__A _13000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09132_ _09940_/A _09132_/B vssd1 vssd1 vccd1 vccd1 _09135_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08624__A1 _08891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08624__B2 _08873_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09063_ _12043_/A _11957_/B _11957_/C vssd1 vssd1 vccd1 vccd1 _12130_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_72_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout213_A _10007_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08014_ _08040_/A _08040_/B vssd1 vssd1 vccd1 vccd1 _08095_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12708__B1 _11688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12184__A1 _12331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12184__B2 _07230_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09965_ _09966_/A _09966_/B vssd1 vssd1 vccd1 vccd1 _09967_/A sky130_fd_sc_hd__and2_1
X_08916_ _08920_/A _08916_/B vssd1 vssd1 vccd1 vccd1 _08916_/X sky130_fd_sc_hd__xor2_1
X_09896_ _09896_/A _09896_/B _09896_/C vssd1 vssd1 vccd1 vccd1 _09897_/B sky130_fd_sc_hd__and3_1
XANTENNA__09888__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09352__A2 _10235_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08847_ _08863_/A _08847_/B vssd1 vssd1 vccd1 vccd1 _08849_/B sky130_fd_sc_hd__xnor2_1
X_08778_ _09674_/S _08778_/B _08778_/C vssd1 vssd1 vccd1 vccd1 _08818_/A sky130_fd_sc_hd__or3_1
XANTENNA__12239__A2 _12793_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08486__A _09671_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09104__A2 _10522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07729_ _10507_/A _07729_/B vssd1 vssd1 vccd1 vccd1 _07811_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10740_ reg1_val[8] curr_PC[8] vssd1 vssd1 vccd1 vccd1 _10741_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_54_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10671_ fanout50/X fanout84/X _08580_/B fanout51/X vssd1 vssd1 vccd1 vccd1 _10672_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08933__B _08933_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12410_ _12411_/A _12411_/B vssd1 vssd1 vccd1 vccd1 _12412_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07418__A2 _10004_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13390_ hold101/X _13416_/A2 _13420_/B1 hold128/X _13383_/A vssd1 vssd1 vccd1 vccd1
+ hold129/A sky130_fd_sc_hd__o221a_1
XFILLER_0_118_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12341_ fanout35/X _07891_/X fanout10/X _07699_/B vssd1 vssd1 vccd1 vccd1 _12342_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12272_ _12272_/A _12272_/B vssd1 vssd1 vccd1 vccd1 _12273_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12175__A1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08918__A2 _07175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11223_ _11223_/A _11223_/B vssd1 vssd1 vccd1 vccd1 _11452_/A sky130_fd_sc_hd__xor2_4
XANTENNA__13372__B1 _13584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12175__B2 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11154_ _07472_/Y _11802_/B _11048_/A _11051_/A vssd1 vssd1 vccd1 vccd1 _11163_/A
+ sky130_fd_sc_hd__a31o_1
X_10105_ _09951_/A _09951_/B _09949_/Y vssd1 vssd1 vccd1 vccd1 _10109_/A sky130_fd_sc_hd__a21bo_2
X_11085_ _11085_/A _11085_/B vssd1 vssd1 vccd1 vccd1 _11099_/A sky130_fd_sc_hd__xor2_1
XANTENNA__09780__A _09949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10036_ _07010_/B _11587_/A2 _10030_/Y _07008_/Y _10035_/X vssd1 vssd1 vccd1 vccd1
+ _10036_/X sky130_fd_sc_hd__o221a_1
XANTENNA__11686__B1 _09521_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11987_ _10342_/A _11984_/X _11986_/X vssd1 vssd1 vccd1 vccd1 dest_val[19] sky130_fd_sc_hd__o21ai_4
XFILLER_0_105_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11989__A1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11989__B2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13726_ _13731_/CLK _13726_/D vssd1 vssd1 vccd1 vccd1 hold266/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08854__A1 _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10938_ _10938_/A _10938_/B vssd1 vssd1 vccd1 vccd1 _10939_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08854__B2 _08907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10661__A1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10869_ _10734_/A _10868_/X _10867_/X vssd1 vssd1 vccd1 vccd1 _10870_/B sky130_fd_sc_hd__o21a_1
XANTENNA__10661__B2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13657_ _13659_/CLK _13657_/D vssd1 vssd1 vccd1 vccd1 hold231/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12608_ _12555_/A _12555_/B _12552_/A vssd1 vssd1 vccd1 vccd1 _12612_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_26_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13588_ _13584_/X _13587_/X _13568_/A vssd1 vssd1 vccd1 vccd1 _13735_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_5_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12539_ _12532_/Y _12533_/X _12538_/Y _12529_/X vssd1 vssd1 vccd1 vccd1 _12539_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07290__B1 _10235_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09955__A _09955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07593__A1 _07594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07194__B _07521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09750_ _10522_/B _09750_/B vssd1 vssd1 vccd1 vccd1 _09751_/A sky130_fd_sc_hd__xnor2_1
X_06962_ _10889_/A reg1_val[9] vssd1 vssd1 vccd1 vccd1 _06962_/Y sky130_fd_sc_hd__nand2b_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08701_ _08701_/A _08701_/B vssd1 vssd1 vccd1 vccd1 _08717_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09334__A2 _10374_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09681_ _09471_/X _09474_/X _09688_/S vssd1 vssd1 vccd1 vccd1 _09681_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11677__B1 _12047_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06893_ _06893_/A _06893_/B vssd1 vssd1 vccd1 vccd1 _07092_/B sky130_fd_sc_hd__nor2_2
XANTENNA__08542__B1 _07556_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11141__A2 _12598_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08632_ _08271_/A _07477_/X _13172_/A1 _09501_/A vssd1 vssd1 vccd1 vccd1 _08633_/B
+ sky130_fd_sc_hd__a22o_1
X_08563_ _08573_/B vssd1 vssd1 vccd1 vccd1 _08563_/Y sky130_fd_sc_hd__inv_2
X_07514_ _07513_/A _07513_/B _07535_/B vssd1 vssd1 vccd1 vccd1 _07517_/C sky130_fd_sc_hd__a21oi_2
XFILLER_0_76_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08494_ _08494_/A vssd1 vssd1 vccd1 vccd1 _08556_/A sky130_fd_sc_hd__inv_2
Xfanout15 _07417_/X vssd1 vssd1 vccd1 vccd1 fanout15/X sky130_fd_sc_hd__buf_4
Xfanout26 fanout27/X vssd1 vssd1 vccd1 vccd1 _08395_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07445_ _07445_/A _07445_/B _07445_/C _07445_/D vssd1 vssd1 vccd1 vccd1 _07453_/B
+ sky130_fd_sc_hd__nand4_2
Xfanout37 _07368_/Y vssd1 vssd1 vccd1 vccd1 _08118_/B sky130_fd_sc_hd__buf_8
XFILLER_0_91_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout48 _07229_/X vssd1 vssd1 vccd1 vccd1 _12268_/A sky130_fd_sc_hd__buf_4
Xfanout59 _10522_/B vssd1 vssd1 vccd1 vccd1 _11825_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07376_ _07377_/A _07377_/B _07376_/C vssd1 vssd1 vccd1 vccd1 _12598_/A sky130_fd_sc_hd__and3_1
X_09115_ _09116_/A _09116_/B vssd1 vssd1 vccd1 vccd1 _09299_/B sky130_fd_sc_hd__and2b_1
XANTENNA__10404__A1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10404__B2 _07833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10076__A _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09046_ _09046_/A _09046_/B _09046_/C vssd1 vssd1 vccd1 vccd1 _09047_/B sky130_fd_sc_hd__and3_1
XFILLER_0_32_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09865__A _12515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13354__B1 _13450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09948_ _09948_/A _09948_/B vssd1 vssd1 vccd1 vccd1 _09950_/B sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout76_A _11423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09879_ curr_PC[0] curr_PC[1] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _09879_/X sky130_fd_sc_hd__a21o_1
XANTENNA__08533__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11910_ fanout38/X _07597_/X _07891_/X _08118_/B vssd1 vssd1 vccd1 vccd1 _11911_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13409__A1 _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07887__A2 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12890_ _13048_/B _12890_/B vssd1 vssd1 vccd1 vccd1 _12891_/B sky130_fd_sc_hd__or2_1
XFILLER_0_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09105__A _10119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11841_ _11841_/A _11841_/B vssd1 vssd1 vccd1 vccd1 _11843_/A sky130_fd_sc_hd__xnor2_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11045__A1_N _11527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _11958_/A _11772_/B _11772_/C vssd1 vssd1 vccd1 vccd1 _11772_/X sky130_fd_sc_hd__and3_1
XFILLER_0_28_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10723_ _10723_/A _10723_/B vssd1 vssd1 vccd1 vccd1 _10981_/C sky130_fd_sc_hd__xnor2_4
XFILLER_0_83_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13511_ hold289/X _13555_/A2 _13510_/X _13542_/B2 vssd1 vssd1 vccd1 vccd1 hold290/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10654_ _10654_/A _10654_/B vssd1 vssd1 vccd1 vccd1 _10656_/B sky130_fd_sc_hd__xnor2_1
X_13442_ hold32/X _13142_/A _13444_/B1 hold123/A _13444_/C1 vssd1 vssd1 vccd1 vccd1
+ hold33/A sky130_fd_sc_hd__o221a_1
XFILLER_0_36_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07279__B _07476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13373_ _13547_/A hold167/X vssd1 vssd1 vccd1 vccd1 hold168/A sky130_fd_sc_hd__and2_1
X_10585_ _10483_/X _10727_/B _10584_/Y vssd1 vssd1 vccd1 vccd1 _10585_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12324_ _12296_/Y _12297_/X _12299_/X _10866_/B _12323_/Y vssd1 vssd1 vccd1 vccd1
+ _12324_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_11_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12255_ _12255_/A _12255_/B vssd1 vssd1 vccd1 vccd1 _12256_/B sky130_fd_sc_hd__or2_1
XFILLER_0_50_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11206_ _11084_/A _11084_/B _11083_/A vssd1 vssd1 vccd1 vccd1 _11211_/A sky130_fd_sc_hd__o21ai_1
X_12186_ _12187_/A _12187_/B _12187_/C vssd1 vssd1 vccd1 vccd1 _12188_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__10433__B _10577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08772__B1 _08923_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11137_ hold291/A _11137_/B vssd1 vssd1 vccd1 vccd1 _11137_/Y sky130_fd_sc_hd__xnor2_2
X_11068_ _11068_/A _11068_/B vssd1 vssd1 vccd1 vccd1 _11069_/B sky130_fd_sc_hd__or2_1
XANTENNA__08524__B1 _08580_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12320__A1 _12710_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10019_ _10456_/S _09488_/X _10601_/C vssd1 vssd1 vccd1 vccd1 _10019_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_92_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12320__B2 _12537_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07878__A2 _11823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07180__D _07363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13709_ _13736_/CLK _13709_/D vssd1 vssd1 vccd1 vccd1 hold283/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07230_ _07230_/A _07230_/B vssd1 vssd1 vccd1 vccd1 _07230_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_27_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10608__B _11688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07161_ reg1_val[5] _07572_/S vssd1 vssd1 vccd1 vccd1 _07161_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07092_ _11961_/A _07092_/B _11774_/A _07092_/D vssd1 vssd1 vccd1 vccd1 _07098_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_0_2_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13336__B1 _13506_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11898__B1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout205 _07137_/Y vssd1 vssd1 vccd1 vccd1 _12760_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout216 _07013_/X vssd1 vssd1 vccd1 vccd1 _10456_/S sky130_fd_sc_hd__buf_4
XFILLER_0_10_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09802_ _09802_/A _09802_/B vssd1 vssd1 vccd1 vccd1 _09804_/B sky130_fd_sc_hd__xnor2_1
Xfanout227 _11252_/B vssd1 vssd1 vccd1 vccd1 _12058_/A sky130_fd_sc_hd__buf_4
Xfanout238 _12327_/A vssd1 vssd1 vccd1 vccd1 _12867_/S sky130_fd_sc_hd__clkbuf_8
X_07994_ _07994_/A _07994_/B vssd1 vssd1 vccd1 vccd1 _07997_/B sky130_fd_sc_hd__xor2_2
Xfanout249 _06744_/Y vssd1 vssd1 vccd1 vccd1 _13142_/A sky130_fd_sc_hd__buf_4
XFILLER_0_5_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07933__A _11286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09733_ _09734_/A _09734_/B vssd1 vssd1 vccd1 vccd1 _09733_/Y sky130_fd_sc_hd__nand2_1
X_06945_ _06928_/A _06936_/B _13042_/B _06944_/X vssd1 vssd1 vccd1 vccd1 _07472_/A
+ sky130_fd_sc_hd__a31o_2
XFILLER_0_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout280_A _13568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09664_ _09440_/X _09447_/X _09703_/B vssd1 vssd1 vccd1 vccd1 _09664_/X sky130_fd_sc_hd__mux2_1
X_06876_ _06876_/A _06876_/B vssd1 vssd1 vccd1 vccd1 _12136_/A sky130_fd_sc_hd__nor2_2
X_08615_ _08615_/A _08615_/B vssd1 vssd1 vccd1 vccd1 _08655_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09595_ fanout40/X fanout75/X _08704_/B fanout56/X vssd1 vssd1 vccd1 vccd1 _09596_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08546_ _08610_/A _08610_/B _08545_/A vssd1 vssd1 vccd1 vccd1 _08577_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12075__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08477_ _08857_/A _08477_/B vssd1 vssd1 vccd1 vccd1 _08480_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_77_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11822__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07428_ reg1_val[19] _07865_/B vssd1 vssd1 vccd1 vccd1 _07429_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_92_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07359_ _07360_/A _07360_/B _07360_/C _07360_/D vssd1 vssd1 vccd1 vccd1 _12177_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08046__A2 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10370_ _10520_/A _10370_/B vssd1 vssd1 vccd1 vccd1 _10371_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_5_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09029_ _08844_/A _08973_/B _08844_/B vssd1 vssd1 vccd1 vccd1 _09029_/Y sky130_fd_sc_hd__a21boi_1
X_12040_ _12695_/A _11988_/X _12164_/B vssd1 vssd1 vccd1 vccd1 _12040_/Y sky130_fd_sc_hd__a21oi_1
Xhold270 hold270/A vssd1 vssd1 vccd1 vccd1 hold270/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 hold281/A vssd1 vssd1 vccd1 vccd1 hold281/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 hold292/A vssd1 vssd1 vccd1 vccd1 hold292/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_12_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12302__A1 _12515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12942_ reg1_val[21] curr_PC[21] _12978_/S vssd1 vssd1 vccd1 vccd1 _12943_/B sky130_fd_sc_hd__mux2_2
X_12873_ _12879_/B _12873_/B vssd1 vssd1 vccd1 vccd1 new_PC[10] sky130_fd_sc_hd__and2_4
X_11824_ _11997_/A fanout8/X fanout3/X _11922_/A vssd1 vssd1 vccd1 vccd1 _11825_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11813__B1 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _11756_/A _11756_/B vssd1 vssd1 vccd1 vccd1 _11853_/B sky130_fd_sc_hd__nand2b_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10706_ _10500_/A _10500_/B _10498_/Y vssd1 vssd1 vccd1 vccd1 _10711_/A sky130_fd_sc_hd__a21bo_1
X_11686_ hold292/A _11685_/X _09521_/Y vssd1 vssd1 vccd1 vccd1 _11686_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13425_ _12094_/A _13445_/A2 hold60/X vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__o21a_1
X_10637_ _10637_/A _12764_/B vssd1 vssd1 vccd1 vccd1 _10641_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10568_ _10569_/B _10569_/A vssd1 vssd1 vccd1 vccd1 _10719_/B sky130_fd_sc_hd__nand2b_1
X_13356_ hold185/X _13506_/B2 _13506_/A2 _13660_/Q vssd1 vssd1 vccd1 vccd1 hold186/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13318__B1 fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12307_ _12305_/Y _12307_/B vssd1 vssd1 vccd1 vccd1 _12309_/A sky130_fd_sc_hd__and2b_1
XANTENNA__12135__S _12578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10499_ _10499_/A _10499_/B vssd1 vssd1 vccd1 vccd1 _10500_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_87_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13287_ _13276_/B _13465_/B _13274_/X vssd1 vssd1 vccd1 vccd1 _13469_/B sky130_fd_sc_hd__a21o_1
X_12238_ _06863_/A _09516_/X _12237_/X vssd1 vssd1 vccd1 vccd1 _12238_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__08745__B1 _08778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12541__A1 _09429_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12169_ _12496_/A fanout16/X fanout12/X _12413_/A vssd1 vssd1 vccd1 vccd1 _12170_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07012__A3 _12995_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07753__A _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10304__B1 _10730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07191__C _11793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08400_ _08350_/B _08313_/C _08313_/B vssd1 vssd1 vccd1 vccd1 _08403_/B sky130_fd_sc_hd__a21oi_1
X_09380_ _09380_/A _09380_/B vssd1 vssd1 vccd1 vccd1 _09389_/A sky130_fd_sc_hd__xor2_1
XANTENNA__08584__A _09373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08331_ _07238_/X _07544_/Y _11638_/A _07239_/Y vssd1 vssd1 vccd1 vccd1 _08332_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06816__B _12981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08262_ _08282_/A _08282_/B vssd1 vssd1 vccd1 vccd1 _08262_/X sky130_fd_sc_hd__and2_1
XANTENNA__10083__A2 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11280__A1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11280__B2 _08580_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07213_ _07213_/A _07213_/B vssd1 vssd1 vccd1 vccd1 _07213_/Y sky130_fd_sc_hd__nand2_1
X_08193_ _11286_/A _08193_/B vssd1 vssd1 vccd1 vccd1 _08255_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12834__A _13005_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13690__CLK _13701_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07144_ instruction[40] _07110_/B _07142_/X _07143_/Y vssd1 vssd1 vccd1 vccd1 _07144_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07075_ _07075_/A vssd1 vssd1 vccd1 vccd1 _07075_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12045__S _12515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10543__B1 _10542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07663__A _09591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ _10078_/A _07977_/B vssd1 vssd1 vccd1 vccd1 _08041_/A sky130_fd_sc_hd__xnor2_2
X_09716_ _09716_/A vssd1 vssd1 vccd1 vccd1 _09716_/Y sky130_fd_sc_hd__inv_2
X_06928_ _06928_/A _06928_/B _13054_/B vssd1 vssd1 vccd1 vccd1 _06928_/X sky130_fd_sc_hd__and3_1
X_09647_ _09648_/A _09648_/B vssd1 vssd1 vccd1 vccd1 _09647_/X sky130_fd_sc_hd__and2_1
X_06859_ reg2_val[22] _06873_/B1 _06872_/B1 _06858_/Y vssd1 vssd1 vccd1 vccd1 _07212_/B
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_97_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11913__A _11913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ _09578_/A _09578_/B vssd1 vssd1 vccd1 vccd1 _09579_/B sky130_fd_sc_hd__nand2_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ _08907_/A fanout76/X fanout74/X _08197_/A vssd1 vssd1 vccd1 vccd1 _08530_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10529__A _11823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11271__A1 _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11540_ _11540_/A _11540_/B vssd1 vssd1 vccd1 vccd1 _11542_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11271__B2 _12103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout5_A fanout5/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11471_ _11471_/A _11471_/B vssd1 vssd1 vccd1 vccd1 _11471_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_80_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09216__A1 _07347_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09216__B2 _09216_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07490__A3 _07363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12744__A _13129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10422_ _10422_/A _10422_/B vssd1 vssd1 vccd1 vccd1 _10424_/A sky130_fd_sc_hd__xnor2_2
X_13210_ hold268/X hold44/X vssd1 vssd1 vccd1 vccd1 _13211_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__09767__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10353_ _10507_/A _10353_/B vssd1 vssd1 vccd1 vccd1 _10360_/A sky130_fd_sc_hd__xnor2_4
X_13141_ _13141_/A _13141_/B vssd1 vssd1 vccd1 vccd1 _13141_/Y sky130_fd_sc_hd__nor2_1
X_13072_ reg1_val[18] _13129_/B vssd1 vssd1 vccd1 vccd1 _13074_/A sky130_fd_sc_hd__or2_1
X_10284_ _10127_/A _10127_/B _10124_/X vssd1 vssd1 vccd1 vccd1 _10286_/B sky130_fd_sc_hd__o21ba_1
X_12023_ _12014_/A _12014_/B _12024_/B vssd1 vssd1 vccd1 vccd1 _12023_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__08669__A _08951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12925_ _12937_/A _12937_/B _12938_/B vssd1 vssd1 vccd1 vccd1 _12926_/B sky130_fd_sc_hd__nand3_1
XANTENNA__07702__A1 _09604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07702__B2 _09748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11823__A _11823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12856_ _12865_/A _12856_/B vssd1 vssd1 vccd1 vccd1 _12858_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_56_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11807_ _11807_/A _11807_/B vssd1 vssd1 vccd1 vccd1 _11821_/A sky130_fd_sc_hd__xnor2_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ hold140/A _12787_/B vssd1 vssd1 vccd1 vccd1 _12787_/Y sky130_fd_sc_hd__xnor2_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11262__A1 _11866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11738_ _11737_/A _11737_/B _11737_/C vssd1 vssd1 vccd1 vccd1 _11739_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11669_ _11231_/A _11601_/X _12163_/A vssd1 vssd1 vccd1 vccd1 _11669_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13408_ _13685_/Q _13416_/A2 _13420_/B1 hold92/X _13383_/A vssd1 vssd1 vccd1 vccd1
+ hold93/A sky130_fd_sc_hd__o221a_1
XANTENNA__09758__A2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12211__B1 _12372_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12762__A1 _09254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13339_ _13359_/A hold241/X vssd1 vssd1 vccd1 vccd1 hold242/A sky130_fd_sc_hd__and2_1
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10773__B1 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07900_ _07900_/A _07900_/B vssd1 vssd1 vccd1 vccd1 _07912_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_20_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08880_ _08878_/Y _08898_/B _08865_/Y vssd1 vssd1 vccd1 vccd1 _08885_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__08579__A _11286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07831_ fanout39/X _08873_/B2 _13149_/A _08118_/B vssd1 vssd1 vccd1 vccd1 _07832_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07762_ _08907_/A fanout47/X fanout45/X _08328_/B2 vssd1 vssd1 vccd1 vccd1 _07763_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09501_ _09501_/A curr_PC[0] vssd1 vssd1 vccd1 vccd1 _09501_/X sky130_fd_sc_hd__or2_1
X_07693_ _07788_/A _07788_/B vssd1 vssd1 vccd1 vccd1 _07713_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09432_ _09432_/A _09432_/B vssd1 vssd1 vccd1 vccd1 _09432_/X sky130_fd_sc_hd__or2_1
XFILLER_0_63_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10528__A2_N fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11452__B _11554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09363_ _09940_/A _09363_/B vssd1 vssd1 vccd1 vccd1 _09367_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08249__A2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout243_A _07108_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08314_ _08350_/B _08313_/B _08313_/C _08310_/Y vssd1 vssd1 vccd1 vccd1 _08343_/A
+ sky130_fd_sc_hd__a31o_2
XANTENNA__07457__B1 _08395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09294_ _09295_/A _09295_/B vssd1 vssd1 vccd1 vccd1 _09296_/A sky130_fd_sc_hd__and2_1
XFILLER_0_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_10 instruction[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_21 instruction[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_32 reg1_val[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08245_ _11708_/A _08245_/B vssd1 vssd1 vccd1 vccd1 _08251_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_43 reg2_val[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_54 reg2_val[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_65 reg2_val[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_76 reg1_val[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08176_ _08176_/A _08176_/B vssd1 vssd1 vccd1 vccd1 _08177_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09749__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07127_ instruction[14] _07129_/B vssd1 vssd1 vccd1 vccd1 dest_idx[3] sky130_fd_sc_hd__and2_4
XANTENNA__10084__A _11709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07058_ _12303_/A _07057_/X _07052_/Y vssd1 vssd1 vccd1 vccd1 _07059_/B sky130_fd_sc_hd__o21a_1
XANTENNA__08709__B1 _11047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08489__A _09591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07932__A1 _07300_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07932__B2 _07541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08488__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10971_ _10972_/A _10972_/B vssd1 vssd1 vccd1 vccd1 _11104_/A sky130_fd_sc_hd__nand2_1
X_12710_ _09504_/Y _09838_/Y _09853_/X _12710_/B2 _12709_/X vssd1 vssd1 vccd1 vccd1
+ _12710_/X sky130_fd_sc_hd__a221o_1
Xmax_cap78 _07526_/Y vssd1 vssd1 vccd1 vccd1 _13174_/A1 sky130_fd_sc_hd__buf_6
XFILLER_0_57_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13690_ _13701_/CLK hold24/X vssd1 vssd1 vccd1 vccd1 _13690_/Q sky130_fd_sc_hd__dfxtp_1
X_12641_ _07082_/Y _12640_/X _12738_/S vssd1 vssd1 vccd1 vccd1 _12642_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_84_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09437__A1 _13135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07448__B1 _07476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09988__A2 _09824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12572_ _12441_/Y _12682_/C _12571_/X vssd1 vssd1 vccd1 vccd1 _12572_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07999__A1 _08486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07999__B2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11523_ _11524_/A _11524_/B vssd1 vssd1 vccd1 vccd1 _11646_/D sky130_fd_sc_hd__and2b_1
XFILLER_0_108_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11454_ _11454_/A _11665_/A vssd1 vssd1 vccd1 vccd1 _11454_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_123_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08948__B1 _09910_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10405_ _12092_/A _10405_/B vssd1 vssd1 vccd1 vccd1 _10407_/B sky130_fd_sc_hd__xnor2_4
X_11385_ _11348_/B _11600_/B _11864_/A vssd1 vssd1 vccd1 vccd1 _11458_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10755__B1 _10753_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13124_ reg1_val[29] _13136_/A vssd1 vssd1 vccd1 vccd1 _13126_/A sky130_fd_sc_hd__nand2_1
X_10336_ _12525_/A _12760_/A1 _10335_/Y _10330_/Y vssd1 vssd1 vccd1 vccd1 _10336_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ _13055_/A _13061_/A vssd1 vssd1 vccd1 vccd1 _13057_/C sky130_fd_sc_hd__nand2_1
X_10267_ fanout40/X fanout25/X fanout23/X fanout56/X vssd1 vssd1 vccd1 vccd1 _10268_/B
+ sky130_fd_sc_hd__o22a_1
X_12006_ _12668_/A _12006_/B vssd1 vssd1 vccd1 vccd1 _12010_/A sky130_fd_sc_hd__xnor2_1
X_10198_ curr_PC[4] _10340_/C vssd1 vssd1 vccd1 vccd1 _10198_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_108_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11483__A1 _09521_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12908_ _12912_/B _12908_/B vssd1 vssd1 vccd1 vccd1 new_PC[15] sky130_fd_sc_hd__and2_4
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12839_ reg1_val[6] curr_PC[6] _12867_/S vssd1 vssd1 vccd1 vccd1 _12841_/B sky130_fd_sc_hd__mux2_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09958__A _10522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08030_ _08030_/A _08030_/B vssd1 vssd1 vccd1 vccd1 _08038_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13199__B _13207_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08939__B1 _07239_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_5_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13725_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09693__A _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07611__B1 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09981_ _09981_/A _09981_/B vssd1 vssd1 vccd1 vccd1 _09982_/B sky130_fd_sc_hd__xor2_4
X_08932_ _09703_/B _08933_/B vssd1 vssd1 vccd1 vccd1 _08944_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_110_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09364__B1 _08704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13160__A1 _07492_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08863_ _08863_/A _08863_/B vssd1 vssd1 vccd1 vccd1 _08879_/A sky130_fd_sc_hd__nor2_1
XANTENNA_fanout193_A _09519_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07814_ _07814_/A _07814_/B vssd1 vssd1 vccd1 vccd1 _07815_/B sky130_fd_sc_hd__nand2_1
X_08794_ _08821_/B2 _08866_/A2 _09216_/B2 _08821_/A1 vssd1 vssd1 vccd1 vccd1 _08795_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07745_ _07747_/A _07745_/B vssd1 vssd1 vccd1 vccd1 _07843_/B sky130_fd_sc_hd__nor2_1
XANTENNA__13463__A2 _13450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12559__A _12666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07678__B1 _09885_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07676_ _10266_/A _07676_/B vssd1 vssd1 vccd1 vccd1 _07680_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07142__A2 _09529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09415_ _09414_/A _09414_/B _09416_/A vssd1 vssd1 vccd1 vccd1 _09415_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11226__A1 _10978_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09346_ _09346_/A _09346_/B vssd1 vssd1 vccd1 vccd1 _09348_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09277_ _09278_/A _09278_/B vssd1 vssd1 vccd1 vccd1 _09277_/X sky130_fd_sc_hd__or2_1
XFILLER_0_117_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10985__B1 _10984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08228_ _08226_/A _08226_/B _08301_/A vssd1 vssd1 vccd1 vccd1 _08240_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_117_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08159_ _08157_/Y _08159_/B vssd1 vssd1 vccd1 vccd1 _08239_/A sky130_fd_sc_hd__and2b_1
XANTENNA__11151__C_N _10900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11170_ _11171_/A _11171_/B vssd1 vssd1 vccd1 vccd1 _11172_/A sky130_fd_sc_hd__and2_1
X_10121_ _10121_/A _10121_/B vssd1 vssd1 vccd1 vccd1 _10122_/B sky130_fd_sc_hd__or2_1
XFILLER_0_30_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11638__A _11638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10542__A _10542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ _10637_/A _07643_/B fanout13/X _10374_/B2 vssd1 vssd1 vccd1 vccd1 _10053_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07905__A1 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07905__B2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13742_ _13742_/CLK hold160/X vssd1 vssd1 vccd1 vccd1 hold159/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12662__B1 _12661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10954_ _10806_/A _10806_/B _10809_/A vssd1 vssd1 vccd1 vccd1 _10956_/B sky130_fd_sc_hd__a21bo_1
X_13673_ _13684_/CLK _13673_/D vssd1 vssd1 vccd1 vccd1 hold149/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10885_ hold295/A _10885_/B vssd1 vssd1 vccd1 vccd1 _11007_/B sky130_fd_sc_hd__or2_1
XANTENNA__13206__A2 _13598_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09778__A _09948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12624_ _12625_/A _12625_/B _12625_/C vssd1 vssd1 vccd1 vccd1 _12626_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_72_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11768__A2 _12163_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12555_ _12555_/A _12555_/B vssd1 vssd1 vccd1 vccd1 _12562_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11506_ fanout29/X _07597_/X _07891_/X fanout27/X vssd1 vssd1 vccd1 vccd1 _11507_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_81_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12486_ _07396_/Y fanout7/X _12485_/X _12417_/A vssd1 vssd1 vccd1 vccd1 _12488_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11437_ _11438_/A _11438_/B _11438_/C vssd1 vssd1 vccd1 vccd1 _11542_/B sky130_fd_sc_hd__a21o_1
XANTENNA__10728__B1 _11151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11368_ hold297/A _11693_/A2 _11582_/C _12533_/B1 vssd1 vssd1 vccd1 vccd1 _11368_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ reg1_val[25] _13136_/A vssd1 vssd1 vccd1 vccd1 _13112_/B sky130_fd_sc_hd__xnor2_2
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10319_ _09835_/X _10318_/X _10457_/S vssd1 vssd1 vccd1 vccd1 _10319_/X sky130_fd_sc_hd__mux2_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11299_ _11299_/A _11299_/B vssd1 vssd1 vccd1 vccd1 _11300_/B sky130_fd_sc_hd__or2_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _13039_/A _13039_/B _13039_/C vssd1 vssd1 vccd1 vccd1 _13045_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08857__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07761__A _09371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13445__A2 _13445_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07530_ _11126_/A _07572_/S vssd1 vssd1 vccd1 vccd1 _07530_/Y sky130_fd_sc_hd__nor2_1
X_07461_ _11281_/A vssd1 vssd1 vccd1 vccd1 _10944_/A sky130_fd_sc_hd__inv_6
XFILLER_0_119_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09200_ _09200_/A _09200_/B vssd1 vssd1 vccd1 vccd1 _09203_/B sky130_fd_sc_hd__xor2_4
X_07392_ _07392_/A _07535_/B vssd1 vssd1 vccd1 vccd1 _07395_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09131_ fanout24/X fanout82/X fanout76/X _08486_/B vssd1 vssd1 vccd1 vccd1 _09132_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08085__B1 _08395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08624__A2 _10522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09062_ _09062_/A _09062_/B vssd1 vssd1 vccd1 vccd1 _12043_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08013_ _10266_/A _08013_/B vssd1 vssd1 vccd1 vccd1 _08040_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout206_A _09161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12184__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06938__A2 _06980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10195__B2 _09529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09964_ _09964_/A _09964_/B vssd1 vssd1 vccd1 vccd1 _09966_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12053__S _12525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08915_ _08897_/B _08913_/X _08912_/X _08903_/Y vssd1 vssd1 vccd1 vccd1 _09016_/B
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__07374__C _07378_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09895_ _09896_/A _09896_/B _09896_/C vssd1 vssd1 vccd1 vccd1 _09897_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__09888__A1 _10374_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09888__B2 _10349_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _08846_/A _08846_/B vssd1 vssd1 vccd1 vccd1 _08849_/A sky130_fd_sc_hd__or2_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11695__A1 _09493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08777_ _08777_/A _08777_/B vssd1 vssd1 vccd1 vccd1 _08778_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__13436__A2 _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08486__B _08486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07728_ fanout85/X fanout75/X _08704_/B fanout82/X vssd1 vssd1 vccd1 vccd1 _07729_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12644__B1 _12695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07659_ _07659_/A _07659_/B vssd1 vssd1 vccd1 vccd1 _07710_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10670_ _10497_/A _10497_/B _10496_/A vssd1 vssd1 vccd1 vccd1 _10682_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_94_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09329_ _07366_/X fanout35/X _07699_/B _07557_/Y vssd1 vssd1 vccd1 vccd1 _09330_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_63_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07418__A3 _09703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12340_ _12666_/A _12340_/B vssd1 vssd1 vccd1 vccd1 _12344_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07823__B1 _08246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12271_ _12272_/A _12272_/B vssd1 vssd1 vccd1 vccd1 _12351_/B sky130_fd_sc_hd__or2_1
XFILLER_0_120_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12175__A2 _12667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11222_ _11222_/A _11222_/B _11223_/B vssd1 vssd1 vccd1 vccd1 _11222_/X sky130_fd_sc_hd__and3_1
XFILLER_0_120_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06750__A _11126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11383__B1 _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06929__A2 _06980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11153_ _11153_/A _11153_/B vssd1 vssd1 vccd1 vccd1 _11219_/A sky130_fd_sc_hd__nand2_1
X_10104_ _10104_/A _10518_/A vssd1 vssd1 vccd1 vccd1 _10110_/A sky130_fd_sc_hd__nand2_2
X_11084_ _11084_/A _11084_/B vssd1 vssd1 vccd1 vccd1 _11085_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11135__B1 _12533_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10035_ _10457_/S _11793_/B _10032_/Y _10033_/X _10034_/X vssd1 vssd1 vccd1 vccd1
+ _10035_/X sky130_fd_sc_hd__o221a_1
XANTENNA__13427__A2 _13445_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11986_ curr_PC[19] _12070_/C _11985_/Y vssd1 vssd1 vccd1 vccd1 _11986_/X sky130_fd_sc_hd__a21o_1
XANTENNA__11989__A2 _07891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13725_ _13725_/CLK _13725_/D vssd1 vssd1 vccd1 vccd1 hold275/A sky130_fd_sc_hd__dfxtp_1
X_10937_ _10937_/A _10937_/B _11027_/A vssd1 vssd1 vccd1 vccd1 _10938_/B sky130_fd_sc_hd__and3_1
XFILLER_0_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08854__A2 _10522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08955__A1_N _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10661__A2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13656_ _13659_/CLK _13656_/D vssd1 vssd1 vccd1 vccd1 hold195/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10868_ _06971_/Y _10734_/B _06973_/B vssd1 vssd1 vccd1 vccd1 _10868_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07520__S _11281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12607_ _12666_/A _12560_/A _12559_/B _12558_/B vssd1 vssd1 vccd1 vccd1 _12621_/A
+ sky130_fd_sc_hd__o31a_1
XANTENNA__10447__A _10734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13587_ hold268/X fanout2/X _13586_/Y _13599_/D vssd1 vssd1 vccd1 vccd1 _13587_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10799_ _11309_/A fanout16/X fanout12/X _07477_/X vssd1 vssd1 vccd1 vccd1 _10800_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12538_ _12710_/B2 _10320_/X _12534_/X _12537_/X vssd1 vssd1 vccd1 vccd1 _12538_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07290__A1 _10235_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07290__B2 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09955__B _10518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12469_ hold207/A _12374_/A _12530_/B _12468_/Y _12795_/A1 vssd1 vssd1 vccd1 vccd1
+ _12475_/C sky130_fd_sc_hd__a311o_1
XFILLER_0_124_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07756__A _10263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11374__B1 _12657_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06961_ _06936_/A _06936_/B _13029_/B _06960_/X vssd1 vssd1 vccd1 vccd1 _10889_/A
+ sky130_fd_sc_hd__a31o_4
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08700_ _08700_/A _08700_/B vssd1 vssd1 vccd1 vccd1 _08727_/A sky130_fd_sc_hd__xnor2_4
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12874__A0 _11126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09680_ _09678_/X _09679_/X _10005_/S vssd1 vssd1 vccd1 vccd1 _09680_/X sky130_fd_sc_hd__mux2_1
X_06892_ _07442_/A _07309_/A vssd1 vssd1 vccd1 vccd1 _06893_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08542__A1 _08806_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07491__A _07492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08631_ _09948_/A _08631_/B vssd1 vssd1 vccd1 vccd1 _08637_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08542__B2 _08806_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13418__A2 _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08562_ _08562_/A _08562_/B vssd1 vssd1 vccd1 vccd1 _08573_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_77_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07513_ _07513_/A _07513_/B vssd1 vssd1 vccd1 vccd1 _07513_/X sky130_fd_sc_hd__and2_1
X_08493_ _11072_/A _08493_/B vssd1 vssd1 vccd1 vccd1 _08494_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout16 _07643_/B vssd1 vssd1 vccd1 vccd1 fanout16/X sky130_fd_sc_hd__clkbuf_8
Xfanout27 _07453_/Y vssd1 vssd1 vccd1 vccd1 fanout27/X sky130_fd_sc_hd__buf_8
XFILLER_0_119_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07444_ _07445_/A _07445_/B _07445_/C _07445_/D vssd1 vssd1 vccd1 vccd1 _11800_/A
+ sky130_fd_sc_hd__a22o_1
Xfanout38 fanout39/X vssd1 vssd1 vccd1 vccd1 fanout38/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout49 _07223_/Y vssd1 vssd1 vccd1 vccd1 fanout49/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_64_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10357__A _11281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07375_ _07634_/D vssd1 vssd1 vccd1 vccd1 _07376_/C sky130_fd_sc_hd__inv_2
X_09114_ _09299_/A _09114_/B vssd1 vssd1 vccd1 vccd1 _09116_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_115_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10404__A2 _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09045_ _09046_/B _09046_/C _09046_/A vssd1 vssd1 vccd1 vccd1 _09047_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07666__A _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09947_ _07175_/X _10536_/A2 fanout6/X _08933_/B vssd1 vssd1 vccd1 vccd1 _09948_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ curr_PC[0] curr_PC[1] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _10041_/B sky130_fd_sc_hd__nand3_2
XANTENNA__08533__A1 _08866_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08533__B2 _08950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08829_ _08850_/A _08850_/B _08825_/Y vssd1 vssd1 vccd1 vccd1 _08836_/B sky130_fd_sc_hd__o21a_1
X_11840_ _11841_/A _11841_/B vssd1 vssd1 vccd1 vccd1 _11935_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10891__A2 _12793_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11771_ _06910_/A _11674_/B _06912_/B vssd1 vssd1 vccd1 vccd1 _11771_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_95_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13510_ hold271/X _13509_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13510_/X sky130_fd_sc_hd__mux2_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _10723_/A _10723_/B vssd1 vssd1 vccd1 vccd1 _10722_/Y sky130_fd_sc_hd__nor2_1
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13441_ _11823_/A _13598_/C hold82/X vssd1 vssd1 vccd1 vccd1 _13702_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10653_ _10544_/B _10546_/B _10654_/B vssd1 vssd1 vccd1 vccd1 _10783_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12396__A2 _12799_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13372_ hold166/X _13542_/B2 _13584_/B _13668_/Q vssd1 vssd1 vccd1 vccd1 hold167/A
+ sky130_fd_sc_hd__a22o_1
X_10584_ _10483_/X _10727_/B _10730_/B vssd1 vssd1 vccd1 vccd1 _10584_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07272__A1 _07535_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12323_ _07137_/Y _12310_/X _12322_/X _12304_/X vssd1 vssd1 vccd1 vccd1 _12323_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_121_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12254_ _12255_/A _12255_/B vssd1 vssd1 vccd1 vccd1 _12334_/B sky130_fd_sc_hd__nand2_1
X_11205_ _11085_/A _11085_/B _11069_/A vssd1 vssd1 vccd1 vccd1 _11215_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12185_ _12764_/B _12185_/B vssd1 vssd1 vccd1 vccd1 _12187_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__08772__A1 _08891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10433__C _10631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08772__B2 _08873_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11136_ hold280/A _11251_/C _11252_/B vssd1 vssd1 vccd1 vccd1 _11137_/B sky130_fd_sc_hd__o21a_1
XANTENNA_max_cap121_A _07455_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11067_ _11068_/A _11068_/B vssd1 vssd1 vccd1 vccd1 _11069_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08524__A1 _09674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08524__B2 _08873_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10018_ _12525_/A _10010_/X _10017_/X _12760_/A1 vssd1 vssd1 vccd1 vccd1 _10018_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11969_ hold259/A _11969_/B vssd1 vssd1 vccd1 vccd1 _12057_/B sky130_fd_sc_hd__or2_1
X_13708_ _13708_/CLK _13708_/D vssd1 vssd1 vccd1 vccd1 hold264/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13639_ _13739_/CLK _13639_/D vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07160_ reg1_val[5] _07160_/B vssd1 vssd1 vccd1 vccd1 _07160_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__09252__A2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07091_ _09659_/A _07091_/B vssd1 vssd1 vccd1 vccd1 _07091_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10905__A _12420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08212__B1 _07477_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13000__B _13000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11898__A1 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11898__B2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout206 _09161_/A vssd1 vssd1 vccd1 vccd1 _09703_/B sky130_fd_sc_hd__buf_6
X_09801_ _09604_/A _10518_/A _09610_/B _09608_/X vssd1 vssd1 vccd1 vccd1 _09802_/B
+ sky130_fd_sc_hd__a31o_1
Xfanout217 _09496_/S vssd1 vssd1 vccd1 vccd1 _10176_/A sky130_fd_sc_hd__clkbuf_8
Xfanout228 _09705_/X vssd1 vssd1 vccd1 vccd1 _11252_/B sky130_fd_sc_hd__buf_2
X_07993_ _07993_/A _07993_/B vssd1 vssd1 vccd1 vccd1 _07997_/A sky130_fd_sc_hd__xnor2_2
Xfanout239 _12971_/S vssd1 vssd1 vccd1 vccd1 _12978_/S sky130_fd_sc_hd__clkbuf_8
X_09732_ _12092_/A _09732_/B vssd1 vssd1 vccd1 vccd1 _09734_/B sky130_fd_sc_hd__xnor2_4
X_06944_ reg2_val[11] _06980_/B vssd1 vssd1 vccd1 vccd1 _06944_/X sky130_fd_sc_hd__and2_1
X_09663_ _09436_/X _09441_/X _09703_/B vssd1 vssd1 vccd1 vccd1 _09663_/X sky130_fd_sc_hd__mux2_1
X_06875_ reg1_val[21] _06875_/B vssd1 vssd1 vccd1 vccd1 _06876_/B sky130_fd_sc_hd__nor2_1
XANTENNA_fanout273_A _13444_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08614_ _08622_/A _08622_/B _08605_/Y vssd1 vssd1 vccd1 vccd1 _08655_/A sky130_fd_sc_hd__a21bo_1
X_09594_ _09940_/A _09594_/B vssd1 vssd1 vccd1 vccd1 _09598_/A sky130_fd_sc_hd__xnor2_2
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08545_ _08545_/A _08545_/B vssd1 vssd1 vccd1 vccd1 _08610_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12075__A1 _12413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12075__B2 _12331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10086__B1 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11822__A1 _12189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08476_ _08806_/A2 _07492_/Y _10637_/A _08806_/B1 vssd1 vssd1 vccd1 vccd1 _08477_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11822__B2 _07198_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07427_ _07652_/A _07652_/B vssd1 vssd1 vccd1 vccd1 _07653_/A sky130_fd_sc_hd__or2_1
XANTENNA__10087__A _11913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07358_ _07360_/C _07360_/D vssd1 vssd1 vccd1 vccd1 _07358_/X sky130_fd_sc_hd__and2_1
XFILLER_0_32_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07289_ _08197_/B _08197_/C vssd1 vssd1 vccd1 vccd1 _07289_/X sky130_fd_sc_hd__or2_1
XANTENNA__10815__A _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09028_ _09028_/A _09028_/B vssd1 vssd1 vccd1 vccd1 _11118_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07396__A _12417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold260 hold260/A vssd1 vssd1 vccd1 vccd1 hold260/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 hold271/A vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 hold282/A vssd1 vssd1 vccd1 vccd1 hold282/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 hold293/A vssd1 vssd1 vccd1 vccd1 hold293/X sky130_fd_sc_hd__dlygate4sd3_1
X_12941_ _12951_/A _12941_/B vssd1 vssd1 vccd1 vccd1 new_PC[20] sky130_fd_sc_hd__xnor2_4
XFILLER_0_87_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12872_ _12872_/A _12872_/B _12872_/C vssd1 vssd1 vccd1 vccd1 _12873_/B sky130_fd_sc_hd__nand3_1
XANTENNA__12066__A1 _09523_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11823_ _11823_/A _11823_/B vssd1 vssd1 vccd1 vccd1 _11830_/A sky130_fd_sc_hd__xnor2_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _11650_/A _11650_/B _11651_/Y vssd1 vssd1 vccd1 vccd1 _11756_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__11813__A1 _12413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11813__B2 _12496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _10557_/A _10556_/B _10556_/A vssd1 vssd1 vccd1 vccd1 _10715_/A sky130_fd_sc_hd__o21ba_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11685_ hold296/A _11881_/D _12058_/A vssd1 vssd1 vccd1 vccd1 _11685_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_102_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13424_ hold59/X _13142_/A _13444_/B1 _13694_/Q _13430_/C1 vssd1 vssd1 vccd1 vccd1
+ hold60/A sky130_fd_sc_hd__o221a_1
X_10636_ _11825_/A _10636_/B vssd1 vssd1 vccd1 vccd1 _10643_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08442__B1 _08580_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13355_ _13359_/A hold204/X vssd1 vssd1 vccd1 vccd1 _13659_/D sky130_fd_sc_hd__and2_1
X_10567_ _10567_/A _10567_/B vssd1 vssd1 vccd1 vccd1 _10569_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13318__B2 _13463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12306_ reg1_val[23] curr_PC[23] vssd1 vssd1 vccd1 vccd1 _12307_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_23_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13286_ _13460_/B _13461_/A _13277_/X vssd1 vssd1 vccd1 vccd1 _13465_/B sky130_fd_sc_hd__a21o_1
X_10498_ _10499_/A _10499_/B vssd1 vssd1 vccd1 vccd1 _10498_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12526__C1 _09529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12237_ _07212_/B _12799_/A2 _11688_/B reg1_val[22] _12236_/X vssd1 vssd1 vccd1 vccd1
+ _12237_/X sky130_fd_sc_hd__o221a_1
XANTENNA__08745__A1 _09674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08745__B2 _08873_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12168_ _12417_/A _12168_/B vssd1 vssd1 vccd1 vccd1 _12260_/A sky130_fd_sc_hd__xnor2_2
X_11119_ _07093_/B _10990_/B _06958_/B vssd1 vssd1 vccd1 vccd1 _11120_/B sky130_fd_sc_hd__o21a_1
X_12099_ _12099_/A _12099_/B vssd1 vssd1 vccd1 vccd1 _12100_/B sky130_fd_sc_hd__and2_1
X_08330_ _08333_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08330_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_47_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10607__A2 _12793_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08261_ _08260_/B _08260_/C _08260_/A vssd1 vssd1 vccd1 vccd1 _08282_/B sky130_fd_sc_hd__o21bai_2
XFILLER_0_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11280__A2 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07212_ _07230_/A _07212_/B _07212_/C vssd1 vssd1 vccd1 vccd1 _07254_/B sky130_fd_sc_hd__nand3_2
X_08192_ _07492_/Y _07541_/X _07545_/Y _10637_/A vssd1 vssd1 vccd1 vccd1 _08193_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11568__B1 _12047_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07143_ is_load _09514_/B vssd1 vssd1 vccd1 vccd1 _07143_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__06832__B _12981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout119_A _07456_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07074_ _12778_/A _07072_/X _07073_/X _06794_/A vssd1 vssd1 vccd1 vccd1 _07075_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12517__C1 _09507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07976_ _08806_/A2 _13174_/A1 _07544_/Y _08806_/B1 vssd1 vssd1 vccd1 vccd1 _07977_/B
+ sky130_fd_sc_hd__a22o_1
X_09715_ _10458_/S _09714_/X _09537_/B vssd1 vssd1 vccd1 vccd1 _09716_/A sky130_fd_sc_hd__o21ai_2
X_06927_ _06927_/A _06927_/B vssd1 vssd1 vccd1 vccd1 _07094_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_97_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09646_ _09646_/A _09646_/B vssd1 vssd1 vccd1 vccd1 _09648_/B sky130_fd_sc_hd__xnor2_2
X_06858_ _06928_/B _13015_/B vssd1 vssd1 vccd1 vccd1 _06858_/Y sky130_fd_sc_hd__nor2_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _09577_/A _09577_/B vssd1 vssd1 vccd1 vccd1 _09578_/B sky130_fd_sc_hd__or2_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06789_ _06936_/A _06789_/B vssd1 vssd1 vccd1 vccd1 _06789_/Y sky130_fd_sc_hd__nand2_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08528_ _09373_/A _08528_/B vssd1 vssd1 vccd1 vccd1 _08532_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07475__A1 _07476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08672__B1 _08778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08459_ _08456_/A _08456_/B _08517_/A vssd1 vssd1 vccd1 vccd1 _08473_/A sky130_fd_sc_hd__o21ba_2
XFILLER_0_107_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11470_ _11362_/A _11362_/B _11360_/B vssd1 vssd1 vccd1 vccd1 _11471_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_18_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09216__A2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10421_ _10421_/A _10421_/B vssd1 vssd1 vccd1 vccd1 _10422_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08424__B1 _11638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11023__A2 _10984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13140_ rst _13584_/B _13140_/C vssd1 vssd1 vccd1 vccd1 _13607_/D sky130_fd_sc_hd__nor3_1
X_10352_ fanout49/X fanout75/X _07546_/X fanout51/X vssd1 vssd1 vccd1 vccd1 _10353_/B
+ sky130_fd_sc_hd__o22a_2
X_13071_ _13071_/A _13081_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[17] sky130_fd_sc_hd__xnor2_4
X_10283_ _10113_/A _10113_/B _10111_/Y vssd1 vssd1 vccd1 vccd1 _10286_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__09924__B1 _10536_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12022_ _12110_/B _12022_/B vssd1 vssd1 vccd1 vccd1 _12024_/B sky130_fd_sc_hd__or2_1
X_12924_ _12937_/B _12938_/B _12937_/A vssd1 vssd1 vccd1 vccd1 _12931_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07702__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12855_ _13020_/B _12855_/B vssd1 vssd1 vccd1 vccd1 _12856_/B sky130_fd_sc_hd__or2_1
XANTENNA__06917__B _07544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11806_ _11710_/A _11710_/B _11708_/Y vssd1 vssd1 vccd1 vccd1 _11807_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_28_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12786_ hold233/A _12746_/X _12786_/B1 vssd1 vssd1 vccd1 vccd1 _12787_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_83_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _11737_/A _11737_/B _11737_/C vssd1 vssd1 vccd1 vccd1 _11739_/A sky130_fd_sc_hd__and3_1
XANTENNA__08663__B1 _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11668_ _11856_/A _11668_/B vssd1 vssd1 vccd1 vccd1 _12163_/A sky130_fd_sc_hd__xnor2_4
X_13407_ _07536_/X _13419_/A2 hold121/X vssd1 vssd1 vccd1 vccd1 hold122/A sky130_fd_sc_hd__o21a_1
XFILLER_0_114_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10619_ _10617_/Y _10619_/B vssd1 vssd1 vccd1 vccd1 _10620_/B sky130_fd_sc_hd__and2b_1
XANTENNA__12211__A1 _12695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11599_ _11794_/C _11598_/Y _12867_/S _11596_/X vssd1 vssd1 vccd1 vccd1 dest_val[15]
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_98_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13338_ hold240/X _13506_/B2 _13506_/A2 _13651_/Q vssd1 vssd1 vccd1 vccd1 hold241/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12762__A2 _12799_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10773__A1 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10773__B2 _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13269_ hold35/X hold294/A vssd1 vssd1 vccd1 vccd1 _13269_/X sky130_fd_sc_hd__and2b_1
XANTENNA__13172__C1 _13543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11286__A _11286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07830_ _07830_/A _07830_/B _07836_/B vssd1 vssd1 vccd1 vccd1 _07968_/A sky130_fd_sc_hd__or3b_1
X_07761_ _09371_/A _07761_/B vssd1 vssd1 vccd1 vccd1 _07970_/A sky130_fd_sc_hd__xnor2_2
X_09500_ _09501_/A curr_PC[0] vssd1 vssd1 vccd1 vccd1 _09696_/A sky130_fd_sc_hd__nand2_1
X_07692_ _09950_/A _07692_/B vssd1 vssd1 vccd1 vccd1 _07788_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09431_ _12695_/A _09881_/A _10726_/A _11955_/A vssd1 vssd1 vccd1 vccd1 _09432_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09362_ fanout25/X fanout74/X fanout70/X fanout23/X vssd1 vssd1 vccd1 vccd1 _09363_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11238__C1 _12047_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08313_ _08350_/B _08313_/B _08313_/C vssd1 vssd1 vccd1 vccd1 _08403_/A sky130_fd_sc_hd__and3_1
XFILLER_0_19_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07457__A1 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09293_ _09293_/A _09293_/B vssd1 vssd1 vccd1 vccd1 _09295_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07457__B2 _10915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_11 instruction[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 reg1_val[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08244_ _08923_/B1 fanout24/X _08486_/B _08866_/A2 vssd1 vssd1 vccd1 vccd1 _08245_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_33 reg1_val[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10461__B1 _12533_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_44 reg2_val[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_55 reg2_val[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_66 reg2_val[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07209__A1 _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_77 reg1_val[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08175_ _08174_/A _08174_/B _08174_/C vssd1 vssd1 vccd1 vccd1 _08178_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07126_ instruction[13] _07129_/B vssd1 vssd1 vccd1 vccd1 dest_idx[2] sky130_fd_sc_hd__and2_4
XFILLER_0_70_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07057_ _12218_/A _07056_/X _07053_/Y vssd1 vssd1 vccd1 vccd1 _07057_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_30_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08709__A1 _08907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08709__B2 _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07674__A _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07932__A2 _07545_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07959_ _07959_/A _07959_/B vssd1 vssd1 vccd1 vccd1 _07962_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_97_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10970_ _10970_/A _10970_/B vssd1 vssd1 vccd1 vccd1 _10972_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09629_ _09630_/A _09630_/B vssd1 vssd1 vccd1 vccd1 _09629_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11492__A2 _11600_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12640_ _06802_/A _06802_/B _12516_/A _12514_/Y _12639_/X vssd1 vssd1 vccd1 vccd1
+ _12640_/X sky130_fd_sc_hd__o41a_1
XFILLER_0_65_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12571_ _12436_/Y _12506_/A _12506_/B vssd1 vssd1 vccd1 vccd1 _12571_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_38_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07999__A2 _10522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11522_ _11522_/A _11522_/B vssd1 vssd1 vccd1 vccd1 _11524_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_80_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11453_ _11224_/Y _11665_/A _11451_/Y vssd1 vssd1 vccd1 vccd1 _11453_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_33_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08948__A1 _08271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10404_ fanout14/X _11309_/A _07526_/Y _07833_/B vssd1 vssd1 vccd1 vccd1 _10405_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08948__B2 _09501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11384_ _11597_/C _11383_/Y _12867_/S _11381_/X vssd1 vssd1 vccd1 vccd1 dest_val[13]
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_21_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10755__B2 _10754_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13123_ _13123_/A _13123_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[28] sky130_fd_sc_hd__xnor2_4
XANTENNA__13586__A fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10335_ _10335_/A _10335_/B vssd1 vssd1 vccd1 vccd1 _10335_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ reg1_val[14] _13054_/B vssd1 vssd1 vccd1 vccd1 _13061_/A sky130_fd_sc_hd__nand2_1
X_10266_ _10266_/A _10266_/B vssd1 vssd1 vccd1 vccd1 _10270_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11704__B1 fanout5/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12005_ _12331_/A fanout16/X fanout12/X _07230_/Y vssd1 vssd1 vccd1 vccd1 _12006_/B
+ sky130_fd_sc_hd__a22o_1
X_10197_ _11866_/A _10159_/Y _10160_/X _10196_/X _10158_/Y vssd1 vssd1 vccd1 vccd1
+ _10197_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_17_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12907_ _12907_/A _12907_/B _12907_/C vssd1 vssd1 vccd1 vccd1 _12908_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_76_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10691__B1 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12838_ _12844_/B _12838_/B vssd1 vssd1 vccd1 vccd1 new_PC[5] sky130_fd_sc_hd__and2_4
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12769_ _12723_/A _12722_/Y _12769_/S vssd1 vssd1 vccd1 vccd1 _12773_/B sky130_fd_sc_hd__mux2_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08862__B _08862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10443__B1 _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08939__A1 _09161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08939__B2 _07399_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07611__A1 _11732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09980_ _09981_/A _09981_/B vssd1 vssd1 vccd1 vccd1 _09980_/X sky130_fd_sc_hd__and2_1
XFILLER_0_122_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07611__B2 _10814_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10913__A _11825_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08931_ _08931_/A _08931_/B vssd1 vssd1 vccd1 vccd1 _08944_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_110_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09364__A1 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09364__B2 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13160__A2 _13196_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08862_ _08862_/A _08862_/B vssd1 vssd1 vccd1 vccd1 _08863_/B sky130_fd_sc_hd__and2_1
X_07813_ _07813_/A _07813_/B _07813_/C vssd1 vssd1 vccd1 vccd1 _07817_/A sky130_fd_sc_hd__and3_1
X_08793_ _08793_/A _08793_/B vssd1 vssd1 vccd1 vccd1 _08815_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13448__B1 _13450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07744_ _07744_/A _07744_/B _07744_/C vssd1 vssd1 vccd1 vccd1 _07745_/B sky130_fd_sc_hd__and3_1
XFILLER_0_74_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07678__A1 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07678__B2 _08395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07675_ _07366_/X fanout21/X _08246_/B _07557_/Y vssd1 vssd1 vccd1 vccd1 _07676_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09414_ _09414_/A _09414_/B vssd1 vssd1 vccd1 vccd1 _09416_/B sky130_fd_sc_hd__nor2_2
X_09345_ _09346_/A _09346_/B vssd1 vssd1 vccd1 vccd1 _09559_/A sky130_fd_sc_hd__or2_1
XFILLER_0_90_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09276_ _09276_/A _09276_/B vssd1 vssd1 vccd1 vccd1 _09278_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_118_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08227_ _08300_/A _08300_/B vssd1 vssd1 vccd1 vccd1 _08301_/A sky130_fd_sc_hd__or2_1
XANTENNA__10095__A _10095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08158_ _08158_/A _08158_/B vssd1 vssd1 vccd1 vccd1 _08159_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07109_ reg1_idx[0] reg1_idx[1] reg1_idx[4] _07109_/D vssd1 vssd1 vccd1 vccd1 int_return
+ sky130_fd_sc_hd__and4_4
XANTENNA__11919__A _11920_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08089_ _08112_/A _08112_/B _08160_/B _08082_/X vssd1 vssd1 vccd1 vccd1 _08111_/A
+ sky130_fd_sc_hd__a31o_1
X_10120_ _10121_/A _10121_/B vssd1 vssd1 vccd1 vccd1 _10253_/A sky130_fd_sc_hd__nand2_2
XANTENNA_fanout99_A _11603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11638__B _11802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10051_ _10051_/A vssd1 vssd1 vccd1 vccd1 _10058_/A sky130_fd_sc_hd__inv_2
XFILLER_0_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07905__A2 _10235_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06748__A _12982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11373__B _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13741_ _13742_/CLK hold145/X vssd1 vssd1 vccd1 vccd1 hold143/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12662__A1 _10866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10953_ _11029_/B _10953_/B vssd1 vssd1 vccd1 vccd1 _10956_/A sky130_fd_sc_hd__or2_1
XANTENNA__08866__B1 _08923_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13672_ _13735_/CLK hold156/X vssd1 vssd1 vccd1 vccd1 hold154/A sky130_fd_sc_hd__dfxtp_1
X_10884_ hold240/A _11693_/A2 _11004_/B _10883_/Y _12533_/B1 vssd1 vssd1 vccd1 vccd1
+ _10893_/C sky130_fd_sc_hd__a311o_1
XFILLER_0_85_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12623_ _12677_/B _12623_/B vssd1 vssd1 vccd1 vccd1 _12625_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07579__A _09575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12554_ _12668_/A _12554_/B vssd1 vssd1 vccd1 vccd1 _12555_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11505_ _11709_/A _11505_/B vssd1 vssd1 vccd1 vccd1 _11510_/A sky130_fd_sc_hd__xnor2_2
X_12485_ _12485_/A fanout5/X vssd1 vssd1 vccd1 vccd1 _12485_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09794__A _10263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11436_ _11436_/A _11436_/B vssd1 vssd1 vccd1 vccd1 _11438_/C sky130_fd_sc_hd__xnor2_1
X_11367_ _11693_/A2 _11582_/C hold297/A vssd1 vssd1 vccd1 vccd1 _11367_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13106_ _13106_/A _13112_/A vssd1 vssd1 vccd1 vccd1 _13108_/A sky130_fd_sc_hd__nand2_2
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10318_ _09680_/X _09689_/X _10600_/S vssd1 vssd1 vccd1 vccd1 _10318_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08203__A _08203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ _11299_/A _11299_/B vssd1 vssd1 vccd1 vccd1 _11300_/A sky130_fd_sc_hd__nand2_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ _13037_/A _13045_/A vssd1 vssd1 vccd1 vccd1 _13039_/C sky130_fd_sc_hd__nand2_1
X_10249_ _10250_/A _10250_/B vssd1 vssd1 vccd1 vccd1 _10249_/X sky130_fd_sc_hd__and2_1
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11283__B _12667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07460_ reg1_val[15] _11585_/A _07572_/S vssd1 vssd1 vccd1 vccd1 _07460_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_69_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07391_ _12534_/A _12534_/B _07156_/Y vssd1 vssd1 vccd1 vccd1 _07395_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_91_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09130_ _09130_/A _09130_/B vssd1 vssd1 vccd1 vccd1 _09154_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08085__A1 _13151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08085__B2 _08866_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09061_ _09060_/B _09060_/C _09068_/B vssd1 vssd1 vccd1 vccd1 _09062_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12169__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08012_ _13149_/A fanout21/X _08246_/B _08923_/B1 vssd1 vssd1 vccd1 vccd1 _08013_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07001__B _10603_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12708__A2 _09520_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11458__B _11458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09963_ _09963_/A _09963_/B vssd1 vssd1 vccd1 vccd1 _09964_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08914_ _08903_/Y _08912_/X _08913_/X _08897_/B vssd1 vssd1 vccd1 vccd1 _09016_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09894_ _09894_/A _09894_/B vssd1 vssd1 vccd1 vccd1 _09896_/C sky130_fd_sc_hd__xnor2_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11144__A1 _12537_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09888__A2 _07643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11144__B2 _12710_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12341__B1 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _08845_/A _08845_/B vssd1 vssd1 vccd1 vccd1 _08846_/B sky130_fd_sc_hd__nor2_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08776_ _08776_/A _08776_/B vssd1 vssd1 vccd1 vccd1 _08791_/A sky130_fd_sc_hd__xnor2_1
X_07727_ _07731_/A _07731_/B vssd1 vssd1 vccd1 vccd1 _07744_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_95_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07658_ _07658_/A _07658_/B vssd1 vssd1 vccd1 vccd1 _07659_/B sky130_fd_sc_hd__xor2_1
X_07589_ fanout49/X _08866_/B2 _08950_/B fanout51/X vssd1 vssd1 vccd1 vccd1 _07590_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09328_ _09249_/A _09249_/B _09262_/B _09263_/X vssd1 vssd1 vccd1 vccd1 _09342_/A
+ sky130_fd_sc_hd__a31o_2
XANTENNA__07399__A _10007_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout14_A _07417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_562 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07823__A1 _08923_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09259_ _09260_/A _09260_/B vssd1 vssd1 vccd1 vccd1 _09259_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07823__B2 _07347_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12270_ _12270_/A _12270_/B vssd1 vssd1 vccd1 vccd1 _12272_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11221_ _11222_/A _11222_/B _11223_/B vssd1 vssd1 vccd1 vccd1 _11221_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_31_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13372__A2 _13542_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11152_ _11222_/A _11222_/B vssd1 vssd1 vccd1 vccd1 _11223_/A sky130_fd_sc_hd__nand2_2
X_10103_ _10103_/A _10103_/B vssd1 vssd1 vccd1 vccd1 _10112_/A sky130_fd_sc_hd__and2_2
X_11083_ _11083_/A _11083_/B vssd1 vssd1 vccd1 vccd1 _11084_/B sky130_fd_sc_hd__nand2_1
X_10034_ _07164_/X _12235_/C _12657_/B1 reg1_val[3] vssd1 vssd1 vccd1 vccd1 _10034_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_98_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11985_ curr_PC[19] _12070_/C _10342_/A vssd1 vssd1 vccd1 vccd1 _11985_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10936_ _10937_/A _10937_/B _11027_/A vssd1 vssd1 vccd1 vccd1 _10938_/A sky130_fd_sc_hd__a21oi_1
X_13724_ _13725_/CLK _13724_/D vssd1 vssd1 vccd1 vccd1 hold298/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10867_ _12515_/S _10867_/B _10867_/C vssd1 vssd1 vccd1 vccd1 _10867_/X sky130_fd_sc_hd__or3_1
X_13655_ _13659_/CLK _13655_/D vssd1 vssd1 vccd1 vccd1 hold193/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12606_ _12577_/X _12582_/X _12605_/Y _12547_/X _12546_/Y vssd1 vssd1 vccd1 vccd1
+ dest_val[27] sky130_fd_sc_hd__o32a_4
XFILLER_0_26_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13586_ fanout2/X _13586_/B vssd1 vssd1 vccd1 vccd1 _13586_/Y sky130_fd_sc_hd__nand2_1
X_10798_ _10798_/A _10798_/B _10798_/C vssd1 vssd1 vccd1 vccd1 _10830_/B sky130_fd_sc_hd__and3_1
XFILLER_0_30_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11071__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12537_ _06849_/C _12793_/A2 _12525_/B _12537_/B2 _12536_/X vssd1 vssd1 vccd1 vccd1
+ _12537_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_54_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07290__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12468_ _12374_/A _12530_/B hold207/A vssd1 vssd1 vccd1 vccd1 _12468_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11419_ _11638_/A fanout9/X fanout3/X _11527_/A vssd1 vssd1 vccd1 vccd1 _11420_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10466__A2_N _12235_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12399_ _07384_/X _07408_/X _12235_/C _12398_/X vssd1 vssd1 vccd1 vccd1 _12399_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_22_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07578__B1 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06960_ reg2_val[9] _06980_/B vssd1 vssd1 vccd1 vccd1 _06960_/X sky130_fd_sc_hd__and2_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06891_ _07442_/A _07309_/A vssd1 vssd1 vccd1 vccd1 _06891_/Y sky130_fd_sc_hd__nand2_1
X_08630_ _08933_/B wire122/A _10637_/A _07175_/X vssd1 vssd1 vccd1 vccd1 _08631_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08542__A2 _07492_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07750__B1 _08246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08561_ _08576_/B _08576_/A vssd1 vssd1 vccd1 vccd1 _08562_/B sky130_fd_sc_hd__nand2b_1
X_07512_ _07531_/A _07571_/A _07324_/C _06923_/A vssd1 vssd1 vccd1 vccd1 _07513_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08492_ _08923_/B1 fanout75/X _08704_/B _08866_/A2 vssd1 vssd1 vccd1 vccd1 _08493_/B
+ sky130_fd_sc_hd__o22a_1
Xfanout17 _07642_/X vssd1 vssd1 vccd1 vccd1 _07643_/B sky130_fd_sc_hd__buf_8
XFILLER_0_71_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07443_ _07445_/C _07445_/D vssd1 vssd1 vccd1 vccd1 _07443_/X sky130_fd_sc_hd__and2_1
Xfanout28 _07447_/X vssd1 vssd1 vccd1 vccd1 fanout28/X sky130_fd_sc_hd__clkbuf_8
Xfanout39 _07362_/X vssd1 vssd1 vccd1 vccd1 fanout39/X sky130_fd_sc_hd__buf_8
XFILLER_0_92_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout149_A _13151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07374_ reg1_val[26] reg1_val[27] _07378_/D vssd1 vssd1 vccd1 vccd1 _07634_/D sky130_fd_sc_hd__or3_4
XFILLER_0_45_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09113_ _09113_/A _09113_/B _09113_/C vssd1 vssd1 vccd1 vccd1 _09114_/B sky130_fd_sc_hd__and3_1
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09044_ _09044_/A _09044_/B _09044_/C _09044_/D vssd1 vssd1 vccd1 vccd1 _09046_/C
+ sky130_fd_sc_hd__nand4_4
XFILLER_0_103_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13354__A2 _13506_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10373__A _11731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09946_ _09946_/A _09946_/B vssd1 vssd1 vccd1 vccd1 _09953_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08778__A _09674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _09832_/X _09834_/X _09839_/Y _09876_/X _12327_/A vssd1 vssd1 vccd1 vccd1
+ _09877_/X sky130_fd_sc_hd__o41a_2
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08533__A2 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08828_ _08828_/A _08828_/B vssd1 vssd1 vccd1 vccd1 _08850_/B sky130_fd_sc_hd__xnor2_2
X_08759_ _08784_/A _08784_/B _08731_/X vssd1 vssd1 vccd1 vccd1 _08786_/B sky130_fd_sc_hd__a21oi_2
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _11562_/A _09048_/X _09049_/Y _11866_/A vssd1 vssd1 vccd1 vccd1 _11770_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _10723_/A _10723_/B vssd1 vssd1 vccd1 vccd1 _10721_/Y sky130_fd_sc_hd__nand2_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13440_ hold81/X _13142_/A _13444_/B1 hold32/X _13568_/A vssd1 vssd1 vccd1 vccd1
+ hold82/A sky130_fd_sc_hd__o221a_1
X_10652_ _10652_/A _10652_/B vssd1 vssd1 vccd1 vccd1 _10654_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_35_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13371_ _13547_/A hold208/X vssd1 vssd1 vccd1 vccd1 _13667_/D sky130_fd_sc_hd__and2_1
XFILLER_0_106_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10583_ _10981_/B _10583_/B vssd1 vssd1 vccd1 vccd1 _10727_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_51_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12322_ _09523_/Y _12312_/Y _12316_/Y _12321_/X vssd1 vssd1 vccd1 vccd1 _12322_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_121_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12253_ _12253_/A _12253_/B vssd1 vssd1 vccd1 vccd1 _12255_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11204_ _11204_/A _11204_/B vssd1 vssd1 vccd1 vccd1 _11217_/A sky130_fd_sc_hd__xor2_1
XANTENNA__12553__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12184_ _12331_/A fanout8/X fanout3/X _07230_/Y vssd1 vssd1 vccd1 vccd1 _12185_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08772__A2 _08866_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10433__D _10857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11135_ hold209/A _11693_/A2 _11133_/X _12533_/B1 vssd1 vssd1 vccd1 vccd1 _11135_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07592__A _10239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11066_ _11066_/A _11066_/B vssd1 vssd1 vccd1 vccd1 _11068_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10730__B _10730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08524__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10017_ _12648_/A _10017_/B _10017_/C vssd1 vssd1 vccd1 vccd1 _10017_/X sky130_fd_sc_hd__or3_1
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_max_cap114_A _07472_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12003__A _12417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06936__A _06936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11968_ _11259_/X _11967_/X _12525_/A vssd1 vssd1 vccd1 vccd1 _11968_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11561__B _11561_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13707_ _13708_/CLK _13707_/D vssd1 vssd1 vccd1 vccd1 hold285/A sky130_fd_sc_hd__dfxtp_2
XANTENNA__11292__B1 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10919_ _11512_/A _10919_/B vssd1 vssd1 vccd1 vccd1 _10927_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11899_ _12417_/A _11899_/B vssd1 vssd1 vccd1 vccd1 _11907_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_73_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13638_ _13742_/CLK _13638_/D vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13569_ _13218_/X _13569_/B vssd1 vssd1 vccd1 vccd1 _13570_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07799__B1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11595__A1 _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07090_ _08197_/A _13145_/A vssd1 vssd1 vccd1 vccd1 _07091_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_124_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13336__A2 _13506_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08212__A1 _08806_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08212__B2 _08806_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11898__A2 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout207 _07029_/X vssd1 vssd1 vccd1 vccd1 _09161_/A sky130_fd_sc_hd__buf_4
X_09800_ _09800_/A _09800_/B vssd1 vssd1 vccd1 vccd1 _09802_/A sky130_fd_sc_hd__xnor2_1
Xfanout218 _11472_/S vssd1 vssd1 vccd1 vccd1 _11575_/S sky130_fd_sc_hd__buf_4
X_07992_ _08092_/A _08092_/B _07980_/X vssd1 vssd1 vccd1 vccd1 _08018_/A sky130_fd_sc_hd__a21o_1
XANTENNA__10921__A _12253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout229 _12314_/A vssd1 vssd1 vccd1 vccd1 _12786_/B1 sky130_fd_sc_hd__buf_4
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07971__B1 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09731_ fanout14/X wire122/X _07455_/Y _07833_/B vssd1 vssd1 vccd1 vccd1 _09732_/B
+ sky130_fd_sc_hd__a22o_1
X_06943_ _06943_/A _06943_/B vssd1 vssd1 vccd1 vccd1 _07094_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09662_ _09659_/A _11562_/A _09660_/Y _09661_/Y _11866_/A vssd1 vssd1 vccd1 vccd1
+ _09662_/X sky130_fd_sc_hd__o311a_1
X_06874_ _07348_/A _07201_/B vssd1 vssd1 vccd1 vccd1 _06876_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07723__B1 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08613_ _08613_/A _08613_/B vssd1 vssd1 vccd1 vccd1 _08622_/B sky130_fd_sc_hd__xnor2_1
X_09593_ _11732_/A fanout23/X fanout70/X fanout25/X vssd1 vssd1 vccd1 vccd1 _09594_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12848__A _13015_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08544_ _08544_/A _08544_/B vssd1 vssd1 vccd1 vccd1 _08545_/B sky130_fd_sc_hd__or2_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12075__A2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10086__A1 _11732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10086__B2 _07310_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08475_ _08475_/A _08475_/B vssd1 vssd1 vccd1 vccd1 _08565_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_37_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11822__A2 _07643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07426_ _07504_/A _07426_/B vssd1 vssd1 vccd1 vccd1 _07652_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_9_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11035__B1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07357_ _07357_/A _07535_/B vssd1 vssd1 vccd1 vccd1 _07360_/D sky130_fd_sc_hd__nand2_1
XANTENNA__12583__A _12695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07288_ _08197_/B _08197_/C vssd1 vssd1 vccd1 vccd1 _11997_/A sky130_fd_sc_hd__nor2_8
XFILLER_0_115_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09027_ _09028_/A _09028_/B vssd1 vssd1 vccd1 vccd1 _09034_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07006__A2 _06936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold250 hold250/A vssd1 vssd1 vccd1 vccd1 hold250/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold261 hold298/X vssd1 vssd1 vccd1 vccd1 hold261/X sky130_fd_sc_hd__buf_1
Xhold272 hold272/A vssd1 vssd1 vccd1 vccd1 hold272/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 hold283/A vssd1 vssd1 vccd1 vccd1 hold283/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 hold294/A vssd1 vssd1 vccd1 vccd1 hold294/X sky130_fd_sc_hd__dlygate4sd3_1
X_09929_ _09929_/A _12667_/A vssd1 vssd1 vccd1 vccd1 _09931_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_99_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12940_ _12941_/B vssd1 vssd1 vccd1 vccd1 _12940_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_87_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12871_ _12872_/A _12872_/B _12872_/C vssd1 vssd1 vccd1 vccd1 _12879_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_68_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11822_ _12189_/A _07643_/B fanout12/X _07198_/Y vssd1 vssd1 vccd1 vccd1 _11823_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09132__A _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10077__B2 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11753_ _11753_/A _11753_/B vssd1 vssd1 vccd1 vccd1 _11756_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11813__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _10704_/A _10704_/B vssd1 vssd1 vccd1 vccd1 _10717_/A sky130_fd_sc_hd__xor2_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ _12225_/A _11682_/Y _11683_/X _12760_/A1 vssd1 vssd1 vccd1 vccd1 _11696_/A
+ sky130_fd_sc_hd__o211a_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10635_ _07455_/Y fanout8/X fanout3/X wire122/X vssd1 vssd1 vccd1 vccd1 _10636_/B
+ sky130_fd_sc_hd__a22o_1
X_13423_ _07484_/X _13445_/A2 hold139/X vssd1 vssd1 vccd1 vccd1 _13693_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_125_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13354_ hold200/X _13506_/B2 _13450_/B hold185/X vssd1 vssd1 vccd1 vccd1 hold204/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08442__A1 _13149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10566_ _10567_/A _10567_/B vssd1 vssd1 vccd1 vccd1 _10719_/A sky130_fd_sc_hd__or2_1
XANTENNA__08442__B2 _08923_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12305_ reg1_val[23] curr_PC[23] vssd1 vssd1 vccd1 vccd1 _12305_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13318__A2 _13450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13285_ _13455_/B _13456_/A _13279_/X vssd1 vssd1 vccd1 vccd1 _13461_/A sky130_fd_sc_hd__a21o_1
X_10497_ _10497_/A _10497_/B vssd1 vssd1 vccd1 vccd1 _10499_/B sky130_fd_sc_hd__xor2_4
X_12236_ _07357_/A _07212_/B _09520_/X vssd1 vssd1 vccd1 vccd1 _12236_/X sky130_fd_sc_hd__a21o_1
XANTENNA__08745__A2 _10538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13528__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12167_ _12557_/B fanout35/X _07699_/B _07597_/X vssd1 vssd1 vccd1 vccd1 _12168_/B
+ sky130_fd_sc_hd__o22a_1
X_11118_ _11118_/A _11118_/B vssd1 vssd1 vccd1 vccd1 _11118_/Y sky130_fd_sc_hd__xnor2_1
X_12098_ _12099_/A _12099_/B vssd1 vssd1 vccd1 vccd1 _12100_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_36_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11049_ _11050_/A _11050_/B vssd1 vssd1 vccd1 vccd1 _11051_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_127_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10304__A2 _10727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12668__A _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08260_ _08260_/A _08260_/B _08260_/C vssd1 vssd1 vccd1 vccd1 _08349_/A sky130_fd_sc_hd__or3_1
X_07211_ _07230_/A _07212_/B _07212_/C vssd1 vssd1 vccd1 vccd1 _07213_/B sky130_fd_sc_hd__and3_1
XFILLER_0_6_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08191_ _09591_/A _08191_/B vssd1 vssd1 vccd1 vccd1 _08255_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07497__A _10266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07142_ instruction[17] _09529_/B _09505_/B _07110_/A vssd1 vssd1 vccd1 vccd1 _07142_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07073_ _07099_/A _07059_/X instruction[6] vssd1 vssd1 vccd1 vccd1 _07073_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_2_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09217__A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07975_ _07978_/A _07978_/B vssd1 vssd1 vccd1 vccd1 _07975_/Y sky130_fd_sc_hd__nand2_1
X_09714_ _11472_/S _09713_/X _09534_/C vssd1 vssd1 vccd1 vccd1 _09714_/X sky130_fd_sc_hd__o21a_1
X_06926_ _06927_/A _06927_/B vssd1 vssd1 vccd1 vccd1 _11465_/A sky130_fd_sc_hd__and2_1
XFILLER_0_93_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09645_ _09646_/B _09646_/A vssd1 vssd1 vccd1 vccd1 _09645_/Y sky130_fd_sc_hd__nand2b_1
X_06857_ instruction[32] _12981_/C vssd1 vssd1 vccd1 vccd1 _13015_/B sky130_fd_sc_hd__and2_4
XANTENNA__12578__A _12578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09576_ _09577_/A _09577_/B vssd1 vssd1 vccd1 vccd1 _09578_/A sky130_fd_sc_hd__nand2_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06788_ instruction[24] _13082_/A _06781_/X instruction[41] _06784_/X vssd1 vssd1
+ vccd1 vccd1 _06789_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_38_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _08821_/B2 _09173_/B2 _11047_/A _08821_/A1 vssd1 vssd1 vccd1 vccd1 _08528_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11256__B1 _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08121__B1 _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08458_ _08516_/B _08458_/B vssd1 vssd1 vccd1 vccd1 _08517_/A sky130_fd_sc_hd__and2b_1
XANTENNA__08672__A1 _13149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08672__B2 _08923_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07409_ _07384_/X _07408_/X _07637_/B vssd1 vssd1 vccd1 vccd1 _07414_/C sky130_fd_sc_hd__a21o_1
X_08389_ _08389_/A _08389_/B vssd1 vssd1 vccd1 vccd1 _08454_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10420_ _10421_/A _10421_/B vssd1 vssd1 vccd1 vccd1 _10420_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_73_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12756__B1 _12799_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08424__A1 _08271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08424__B2 _09501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10351_ _10351_/A _10351_/B vssd1 vssd1 vccd1 vccd1 _10383_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_20_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13070_ reg1_val[17] _13129_/B vssd1 vssd1 vccd1 vccd1 _13081_/B sky130_fd_sc_hd__xnor2_4
X_10282_ _10282_/A _10282_/B vssd1 vssd1 vccd1 vccd1 _10287_/A sky130_fd_sc_hd__or2_2
X_12021_ _12021_/A _12021_/B vssd1 vssd1 vccd1 vccd1 _12022_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09924__A1 _12496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09924__B2 _07257_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09127__A _10095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12923_ _12910_/B _12915_/B _12956_/A vssd1 vssd1 vccd1 vccd1 _12938_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__11495__B1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07163__A1 _07535_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12854_ _13020_/B _12855_/B vssd1 vssd1 vccd1 vccd1 _12865_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_96_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11247__B1 _12648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11805_ _11805_/A _11805_/B vssd1 vssd1 vccd1 vccd1 _11807_/A sky130_fd_sc_hd__nor2_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ hold154/A _12785_/B vssd1 vssd1 vccd1 vccd1 _12785_/Y sky130_fd_sc_hd__xnor2_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08663__A1 _07175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11736_ _11736_/A _11736_/B vssd1 vssd1 vccd1 vccd1 _11737_/C sky130_fd_sc_hd__nor2_1
XANTENNA__08663__B2 _08933_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11667_ _10724_/A _11227_/Y _11665_/Y _11666_/Y vssd1 vssd1 vccd1 vccd1 _11668_/B
+ sky130_fd_sc_hd__o31ai_4
XFILLER_0_36_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13406_ hold120/X _13416_/A2 _13420_/B1 _13685_/Q _13383_/A vssd1 vssd1 vccd1 vccd1
+ hold121/A sky130_fd_sc_hd__o221a_1
X_10618_ _13015_/A curr_PC[7] vssd1 vssd1 vccd1 vccd1 _10619_/B sky130_fd_sc_hd__nand2_1
X_11598_ curr_PC[15] _11490_/B _10342_/A vssd1 vssd1 vccd1 vccd1 _11598_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07110__A _07110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10549_ _10686_/A _10548_/C _10391_/A vssd1 vssd1 vccd1 vccd1 _10550_/C sky130_fd_sc_hd__a21bo_1
X_13337_ _13359_/A hold164/X vssd1 vssd1 vccd1 vccd1 hold165/A sky130_fd_sc_hd__and2_1
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10773__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13268_ hold287/X hold73/X vssd1 vssd1 vccd1 vccd1 _13478_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_121_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12219_ _12218_/A _12218_/B _09506_/X vssd1 vssd1 vccd1 vccd1 _12219_/X sky130_fd_sc_hd__o21a_1
X_13199_ hold42/X _13207_/B vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__or2_1
X_07760_ fanout56/X _08866_/B2 _08950_/B fanout53/X vssd1 vssd1 vccd1 vccd1 _07761_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09471__S _09493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07691_ _08328_/B2 fanout49/X fanout45/X _08907_/A vssd1 vssd1 vccd1 vccd1 _07692_/B
+ sky130_fd_sc_hd__o22a_1
X_09430_ _12695_/A _09881_/A _10726_/A vssd1 vssd1 vccd1 vccd1 _09432_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09361_ _09591_/A _09361_/B vssd1 vssd1 vccd1 vccd1 _09369_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11789__A1 _09521_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08312_ _08350_/A _08278_/C _08278_/B vssd1 vssd1 vccd1 vccd1 _08313_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_74_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11789__B2 _09523_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09292_ _09293_/A _09293_/B vssd1 vssd1 vccd1 vccd1 _09414_/B sky130_fd_sc_hd__and2b_1
XANTENNA__07457__A2 _10049_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07004__B _07110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_12 instruction[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ _08243_/A _08243_/B vssd1 vssd1 vccd1 vccd1 _08294_/A sky130_fd_sc_hd__xnor2_2
XANTENNA_23 reg1_val[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09500__A _09501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_34 reg1_val[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout131_A _07285_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_45 reg2_val[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_56 reg2_val[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout229_A _12314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_67 rst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08174_ _08174_/A _08174_/B _08174_/C vssd1 vssd1 vccd1 vccd1 _08178_/A sky130_fd_sc_hd__and3_1
XANTENNA__07209__A2 _07572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_78 reg1_val[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07125_ instruction[12] _07129_/B vssd1 vssd1 vccd1 vccd1 dest_idx[1] sky130_fd_sc_hd__and2_4
XANTENNA__12861__A _13025_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07056_ _12136_/A _07055_/Y _07054_/Y vssd1 vssd1 vccd1 vccd1 _07056_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_2_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08709__A2 _09173_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12800__S _12867_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07958_ _07958_/A _07958_/B vssd1 vssd1 vccd1 vccd1 _07959_/B sky130_fd_sc_hd__xor2_4
XANTENNA__07690__A _08951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06909_ reg1_val[16] _06911_/B vssd1 vssd1 vccd1 vccd1 _06910_/A sky130_fd_sc_hd__or2_1
X_07889_ _07062_/B _07595_/A _07476_/B _09254_/B vssd1 vssd1 vccd1 vccd1 _07892_/A
+ sky130_fd_sc_hd__a211o_4
XFILLER_0_97_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09628_ _09387_/A _09387_/B _09385_/X vssd1 vssd1 vccd1 vccd1 _09630_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_97_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09559_ _09559_/A _09559_/B _09559_/C vssd1 vssd1 vccd1 vccd1 _09560_/B sky130_fd_sc_hd__and3_1
XFILLER_0_78_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10437__D1 _10857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12570_ _12570_/A _12627_/A vssd1 vssd1 vccd1 vccd1 _12682_/C sky130_fd_sc_hd__nor2_1
X_11521_ _11521_/A _11521_/B _11522_/B vssd1 vssd1 vccd1 vccd1 _11646_/C sky130_fd_sc_hd__and3_1
XFILLER_0_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11452_ _11452_/A _11554_/A vssd1 vssd1 vccd1 vccd1 _11665_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_61_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10403_ _12094_/A _10403_/B vssd1 vssd1 vccd1 vccd1 _10407_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08948__A2 _07399_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11383_ curr_PC[13] _11266_/B _10342_/A vssd1 vssd1 vccd1 vccd1 _11383_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_104_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10755__A2 _11587_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13122_ _13112_/X _13121_/X _13136_/A _07634_/D vssd1 vssd1 vccd1 vccd1 _13123_/B
+ sky130_fd_sc_hd__a2bb2o_2
X_10334_ _10332_/Y _10334_/B vssd1 vssd1 vccd1 vccd1 _10335_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_104_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13053_ reg1_val[14] _13054_/B vssd1 vssd1 vccd1 vccd1 _13055_/A sky130_fd_sc_hd__or2_1
X_10265_ _11732_/A fanout18/X fanout70/X fanout20/X vssd1 vssd1 vccd1 vccd1 _10266_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11704__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10189__A2_N _12235_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11704__B2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12004_ _12004_/A vssd1 vssd1 vccd1 vccd1 _12011_/A sky130_fd_sc_hd__inv_2
X_10196_ _12047_/C1 _10164_/Y _10165_/X _10195_/Y vssd1 vssd1 vccd1 vccd1 _10196_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06928__B _06928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12906_ _12907_/A _12907_/B _12907_/C vssd1 vssd1 vccd1 vccd1 _12912_/B sky130_fd_sc_hd__a21o_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10691__A1 _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10691__B2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12837_ _12837_/A _12837_/B _12837_/C vssd1 vssd1 vccd1 vccd1 _12838_/B sky130_fd_sc_hd__nand3_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13541__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12768_ _12768_/A _12768_/B vssd1 vssd1 vccd1 vccd1 _12773_/A sky130_fd_sc_hd__xnor2_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11719_ _11719_/A _11719_/B vssd1 vssd1 vccd1 vccd1 _11722_/A sky130_fd_sc_hd__xnor2_1
X_12699_ reg1_val[28] _12698_/C reg1_val[29] vssd1 vssd1 vccd1 vccd1 _12699_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08939__A2 _07238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07611__A2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11297__A _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08930_ _08929_/B _08938_/A _08916_/X vssd1 vssd1 vccd1 vccd1 _08967_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09364__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08861_ _08861_/A _08861_/B _08861_/C vssd1 vssd1 vccd1 vccd1 _08974_/A sky130_fd_sc_hd__or3_1
X_07812_ _07770_/A _07770_/C _07770_/B vssd1 vssd1 vccd1 vccd1 _07813_/C sky130_fd_sc_hd__o21ai_1
X_08792_ _08793_/A _08793_/B vssd1 vssd1 vccd1 vccd1 _08814_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07180__A_N _07492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13448__A1 _13463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07743_ _07741_/A _07741_/B _07830_/A vssd1 vssd1 vccd1 vccd1 _07843_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__11459__B1 _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout179_A _09373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07674_ _09940_/A _07674_/B vssd1 vssd1 vccd1 vccd1 _07680_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07678__A2 _07491_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09413_ _09279_/A _09279_/B _09277_/X vssd1 vssd1 vccd1 vccd1 _09416_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_47_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09344_ _09239_/A _09239_/B _09237_/Y vssd1 vssd1 vccd1 vccd1 _09346_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09275_ _09275_/A _09275_/B vssd1 vssd1 vccd1 vccd1 _09276_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_90_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08226_ _08226_/A _08226_/B vssd1 vssd1 vccd1 vccd1 _08300_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13384__B1 _09950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08157_ _08158_/A _08158_/B vssd1 vssd1 vccd1 vccd1 _08157_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_43_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07108_ reg1_idx[5] reg1_idx[2] reg1_idx[3] _07108_/D vssd1 vssd1 vccd1 vccd1 _07109_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_0_30_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08088_ _08088_/A _08088_/B vssd1 vssd1 vccd1 vccd1 _08160_/B sky130_fd_sc_hd__xnor2_2
X_07039_ _10867_/B _10867_/C _10870_/A vssd1 vssd1 vccd1 vccd1 _07039_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10050_ _10050_/A _10050_/B vssd1 vssd1 vccd1 vccd1 _10051_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11698__B1 _11672_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08315__B1 _08580_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13740_ _13742_/CLK hold16/X vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08866__A1 _08950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10952_ _10952_/A _10952_/B vssd1 vssd1 vccd1 vccd1 _10953_/B sky130_fd_sc_hd__and2_1
XANTENNA__08866__B2 _08866_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10673__A1 _07546_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11870__B1 _12047_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10673__B2 _12557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13671_ _13735_/CLK _13671_/D vssd1 vssd1 vccd1 vccd1 hold224/A sky130_fd_sc_hd__dfxtp_1
X_10883_ _11693_/A2 _11004_/B hold240/A vssd1 vssd1 vccd1 vccd1 _10883_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12622_ _12677_/A _12621_/C _12621_/A vssd1 vssd1 vccd1 vccd1 _12623_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_66_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12485__B fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12553_ fanout12/X _09145_/Y fanout7/X fanout16/X vssd1 vssd1 vccd1 vccd1 _12554_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11504_ fanout25/X _09146_/Y fanout5/A fanout23/X vssd1 vssd1 vccd1 vccd1 _11505_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_124_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12484_ _12668_/A _12484_/B vssd1 vssd1 vccd1 vccd1 _12488_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12178__B2 _12253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11435_ _11436_/A _11436_/B vssd1 vssd1 vccd1 vccd1 _11542_/A sky130_fd_sc_hd__or2_1
XFILLER_0_124_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10189__B1 _12657_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11366_ hold214/A _11366_/B vssd1 vssd1 vccd1 vccd1 _11582_/C sky130_fd_sc_hd__or2_1
XFILLER_0_104_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13105_ _13105_/A _13105_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[24] sky130_fd_sc_hd__xnor2_4
X_10317_ _10315_/X _10316_/X _11575_/S vssd1 vssd1 vccd1 vccd1 _10317_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11297_ _11507_/A _11297_/B vssd1 vssd1 vccd1 vccd1 _11299_/B sky130_fd_sc_hd__xnor2_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12006__A _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13036_ reg1_val[11] _13036_/B vssd1 vssd1 vccd1 vccd1 _13045_/A sky130_fd_sc_hd__nand2_1
X_10248_ _11076_/A _10248_/B vssd1 vssd1 vccd1 vccd1 _10250_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11689__B1 _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10179_ _10019_/X _10178_/Y _10457_/S vssd1 vssd1 vccd1 vccd1 _10179_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08306__B1 _13166_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09503__C1 _09529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07390_ _07377_/A _07377_/B _07377_/C _07392_/A vssd1 vssd1 vccd1 vccd1 _12534_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09267__D1 _13135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08085__A2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09060_ _09068_/B _09060_/B _09060_/C vssd1 vssd1 vccd1 vccd1 _09062_/A sky130_fd_sc_hd__and3_1
XFILLER_0_4_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12169__A1 _12496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08011_ _10263_/A _08011_/B vssd1 vssd1 vccd1 vccd1 _08040_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12169__B2 _12413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09962_ _09963_/A _09963_/B vssd1 vssd1 vccd1 vccd1 _09962_/Y sky130_fd_sc_hd__nand2_1
X_08913_ _08897_/A _08896_/B _08896_/C _08896_/D vssd1 vssd1 vccd1 vccd1 _08913_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09893_ _09893_/A _09893_/B vssd1 vssd1 vccd1 vccd1 _09894_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12341__A1 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12341__B2 _07699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08844_ _08844_/A _08844_/B vssd1 vssd1 vccd1 vccd1 _09028_/A sky130_fd_sc_hd__and2_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10352__B1 _07546_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08775_ _08804_/A _08804_/B _08771_/X vssd1 vssd1 vccd1 vccd1 _08776_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_79_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07726_ _09591_/A _07726_/B vssd1 vssd1 vccd1 vccd1 _07731_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07657_ _07658_/A _07658_/B vssd1 vssd1 vccd1 vccd1 _07657_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_67_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11490__A _12867_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07588_ _07588_/A _07588_/B vssd1 vssd1 vccd1 vccd1 _07649_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_48_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09327_ _09306_/A _09306_/B _09307_/Y vssd1 vssd1 vccd1 vccd1 _09424_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_48_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11604__B1 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09258_ _09949_/A _09258_/B vssd1 vssd1 vccd1 vccd1 _09260_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__07823__A2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08209_ _10049_/A2 _10538_/A _08778_/B _09173_/B2 vssd1 vssd1 vccd1 vccd1 _08210_/B
+ sky130_fd_sc_hd__o22a_1
X_09189_ _07929_/A _07929_/B _07926_/Y vssd1 vssd1 vccd1 vccd1 _09192_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_16_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11220_ _11340_/B _11220_/B vssd1 vssd1 vccd1 vccd1 _11223_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_120_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11151_ _11151_/A _11151_/B _10900_/B _11150_/X vssd1 vssd1 vccd1 vccd1 _12372_/A
+ sky130_fd_sc_hd__or4bb_4
X_10102_ _10102_/A _10102_/B vssd1 vssd1 vccd1 vccd1 _10103_/B sky130_fd_sc_hd__nand2_1
X_11082_ _11082_/A _11082_/B vssd1 vssd1 vccd1 vccd1 _11083_/B sky130_fd_sc_hd__nand2_1
X_10033_ hold264/A _12314_/A _10031_/X _12796_/A1 vssd1 vssd1 vccd1 vccd1 _10033_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10343__B1 _12825_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11984_ _07281_/A _11793_/B _07152_/X _11983_/X vssd1 vssd1 vccd1 vccd1 _11984_/X
+ sky130_fd_sc_hd__o22a_1
X_13723_ _13725_/CLK _13723_/D vssd1 vssd1 vccd1 vccd1 hold259/A sky130_fd_sc_hd__dfxtp_1
X_10935_ _07575_/X fanout6/X _10934_/Y _11076_/A vssd1 vssd1 vccd1 vccd1 _11027_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12496__A _12496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13654_ _13659_/CLK _13654_/D vssd1 vssd1 vccd1 vccd1 hold297/A sky130_fd_sc_hd__dfxtp_1
X_10866_ _10866_/A _10866_/B _10864_/X vssd1 vssd1 vccd1 vccd1 _10866_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_85_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12605_ _10866_/B _12584_/Y _12604_/X vssd1 vssd1 vccd1 vccd1 _12605_/Y sky130_fd_sc_hd__o21ai_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13585_ _13585_/A _13585_/B vssd1 vssd1 vccd1 vccd1 _13586_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10797_ _10798_/A _10798_/B _10798_/C vssd1 vssd1 vccd1 vccd1 _10830_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07102__B _13748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11071__B2 _07546_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12536_ _06837_/Y _09515_/Y _09519_/Y _06840_/B _12535_/X vssd1 vssd1 vccd1 vccd1
+ _12536_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_109_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13348__B1 _13506_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12467_ hold216/A _12467_/B vssd1 vssd1 vccd1 vccd1 _12530_/B sky130_fd_sc_hd__or2_1
XFILLER_0_34_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11418_ _11538_/B _11418_/B vssd1 vssd1 vccd1 vccd1 _11428_/A sky130_fd_sc_hd__or2_1
XANTENNA__07578__A1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12398_ _12382_/A _12709_/A2 _09515_/Y _06847_/B _12397_/Y vssd1 vssd1 vccd1 vccd1
+ _12398_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11374__A2 _11793_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07578__B2 _11732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11349_ _11864_/A _11348_/B _11600_/B vssd1 vssd1 vccd1 vccd1 _11349_/X sky130_fd_sc_hd__a21o_1
XANTENNA__08527__B1 _11047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13019_ reg1_val[8] _13020_/B vssd1 vssd1 vccd1 vccd1 _13019_/Y sky130_fd_sc_hd__nor2_1
X_06890_ reg1_val[18] _07310_/A vssd1 vssd1 vccd1 vccd1 _06893_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07750__A1 _08866_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07750__B2 _07366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08560_ _08560_/A _08560_/B vssd1 vssd1 vccd1 vccd1 _08576_/B sky130_fd_sc_hd__xor2_1
X_07511_ _10507_/A vssd1 vssd1 vccd1 vccd1 _11286_/A sky130_fd_sc_hd__inv_8
X_08491_ _08746_/A _08491_/B vssd1 vssd1 vccd1 vccd1 _08495_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10919__A _11512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07442_ _07442_/A _07637_/B vssd1 vssd1 vccd1 vccd1 _07445_/D sky130_fd_sc_hd__nand2_1
Xfanout18 _07493_/Y vssd1 vssd1 vccd1 vccd1 fanout18/X sky130_fd_sc_hd__clkbuf_8
Xfanout29 _07447_/X vssd1 vssd1 vccd1 vccd1 fanout29/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_29_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13014__B _13015_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07373_ reg1_val[24] reg1_val[25] vssd1 vssd1 vccd1 vccd1 _07378_/D sky130_fd_sc_hd__or2_2
XFILLER_0_84_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09112_ _09113_/A _09113_/B _09113_/C vssd1 vssd1 vccd1 vccd1 _09299_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09043_ _08726_/A _08726_/B _09042_/X vssd1 vssd1 vccd1 vccd1 _09046_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__09007__A1 _08951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout211_A _09381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06851__B _12981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap173 _07462_/B vssd1 vssd1 vccd1 vccd1 _07377_/A sky130_fd_sc_hd__buf_2
XFILLER_0_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09945_ _09945_/A _09945_/B vssd1 vssd1 vccd1 vccd1 _09946_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08778__B _08778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _09853_/X _09860_/Y _09862_/Y _09523_/Y _09875_/Y vssd1 vssd1 vccd1 vccd1
+ _09876_/X sky130_fd_sc_hd__a221o_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _08951_/A _08827_/B vssd1 vssd1 vccd1 vccd1 _08850_/A sky130_fd_sc_hd__xnor2_2
X_08758_ _08758_/A _08758_/B vssd1 vssd1 vccd1 vccd1 _08784_/B sky130_fd_sc_hd__xor2_4
X_07709_ _07709_/A _07709_/B vssd1 vssd1 vccd1 vccd1 _07964_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ _08687_/A _08687_/B _08729_/A vssd1 vssd1 vccd1 vccd1 _08699_/A sky130_fd_sc_hd__o21bai_4
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ _10852_/B _10720_/B vssd1 vssd1 vccd1 vccd1 _10723_/B sky130_fd_sc_hd__and2_2
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10651_ _10652_/A _10652_/B vssd1 vssd1 vccd1 vccd1 _10813_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_36_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10582_ _09991_/B _10579_/C _10581_/Y vssd1 vssd1 vccd1 vccd1 _10583_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13370_ hold207/X _13563_/B2 _13584_/B hold166/X vssd1 vssd1 vccd1 vccd1 hold208/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12250__B1 _07891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12321_ _07336_/Y _07340_/X _12235_/C _12320_/X vssd1 vssd1 vccd1 vccd1 _12321_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12002__B1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12252_ _12252_/A _12253_/B vssd1 vssd1 vccd1 vccd1 _12334_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12553__A1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11203_ _11203_/A _11203_/B vssd1 vssd1 vccd1 vccd1 _11204_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12553__B2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12183_ _12173_/B _12086_/B _12088_/B _12100_/A vssd1 vssd1 vccd1 vccd1 _12195_/A
+ sky130_fd_sc_hd__a31o_1
X_11134_ _11693_/A2 _11133_/X hold209/A vssd1 vssd1 vccd1 vccd1 _11134_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11065_ _11065_/A _11065_/B vssd1 vssd1 vccd1 vccd1 _11066_/B sky130_fd_sc_hd__nor2_1
X_10016_ _10016_/A _10016_/B _10016_/C vssd1 vssd1 vccd1 vccd1 _10017_/C sky130_fd_sc_hd__and3_1
XFILLER_0_116_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_max_cap107_A _07556_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11967_ _11967_/A _11967_/B vssd1 vssd1 vccd1 vccd1 _11967_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_59_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06936__B _06936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13706_ _13708_/CLK hold263/X vssd1 vssd1 vccd1 vccd1 hold262/A sky130_fd_sc_hd__dfxtp_2
XANTENNA__11292__A1 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07496__B1 _08246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10918_ fanout56/X fanout20/X _08246_/B fanout53/X vssd1 vssd1 vccd1 vccd1 _10919_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_128_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11292__B2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11898_ fanout46/X fanout34/X fanout32/X fanout50/X vssd1 vssd1 vccd1 vccd1 _11899_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_41_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07113__A _13748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13637_ _13739_/CLK _13637_/D vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__dfxtp_1
X_10849_ _10849_/A _10849_/B vssd1 vssd1 vccd1 vccd1 _10852_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_27_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13568_ _13568_/A hold274/X vssd1 vssd1 vccd1 vccd1 _13731_/D sky130_fd_sc_hd__and2_1
XANTENNA__07799__A1 _08821_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07799__B2 _08821_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12519_ _12130_/A _09082_/X _09087_/X _10866_/B vssd1 vssd1 vccd1 vccd1 _12519_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_81_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13499_ _13499_/A _13499_/B vssd1 vssd1 vccd1 vccd1 _13499_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08748__B1 _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08212__A2 _13168_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09474__S _09493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout208 _09671_/S vssd1 vssd1 vccd1 vccd1 _09674_/S sky130_fd_sc_hd__clkbuf_8
Xfanout219 _07419_/A vssd1 vssd1 vccd1 vccd1 _11472_/S sky130_fd_sc_hd__buf_4
X_07991_ _07991_/A _07991_/B vssd1 vssd1 vccd1 vccd1 _08092_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07971__A1 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09730_ _11731_/A _09730_/B vssd1 vssd1 vccd1 vccd1 _09734_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__07971__B2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06942_ _06943_/A _06943_/B vssd1 vssd1 vccd1 vccd1 _11237_/A sky130_fd_sc_hd__and2_1
XANTENNA__09173__B1 _08246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13009__B _13010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09661_ _09659_/A _12742_/A _09660_/Y vssd1 vssd1 vccd1 vccd1 _09661_/Y sky130_fd_sc_hd__o21ai_1
X_06873_ _06871_/Y _06906_/B1 _06873_/B1 reg2_val[21] vssd1 vssd1 vccd1 vccd1 _06875_/B
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07723__A1 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07723__B2 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08612_ _08609_/A _08609_/B _08659_/A vssd1 vssd1 vccd1 vccd1 _08622_/A sky130_fd_sc_hd__o21bai_1
XANTENNA__07007__B _10457_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09592_ _09599_/A vssd1 vssd1 vccd1 vccd1 _09592_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08543_ _08857_/A _08543_/B vssd1 vssd1 vccd1 vccd1 _08610_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout161_A _13598_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10086__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08474_ _08475_/A _08475_/B vssd1 vssd1 vccd1 vccd1 _08474_/X sky130_fd_sc_hd__and2_1
XFILLER_0_9_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07425_ _07425_/A _07425_/B vssd1 vssd1 vccd1 vccd1 _07426_/B sky130_fd_sc_hd__or2_1
XFILLER_0_17_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11035__A1 _07299_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07356_ _12235_/A _12235_/B _07637_/B vssd1 vssd1 vccd1 vccd1 _07360_/C sky130_fd_sc_hd__a21o_1
XANTENNA__11035__B2 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07287_ _07287_/A _07287_/B vssd1 vssd1 vccd1 vccd1 _08197_/C sky130_fd_sc_hd__and2_2
XFILLER_0_17_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07169__S _07572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09026_ _09025_/A _09025_/B _10864_/B _10864_/C vssd1 vssd1 vccd1 vccd1 _11117_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12535__B2 _10889_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold240 hold240/A vssd1 vssd1 vccd1 vccd1 hold240/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07006__A3 _13000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold251 hold300/X vssd1 vssd1 vccd1 vccd1 hold251/X sky130_fd_sc_hd__buf_1
XFILLER_0_40_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold262 hold262/A vssd1 vssd1 vccd1 vccd1 hold262/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 hold273/A vssd1 vssd1 vccd1 vccd1 hold273/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 hold284/A vssd1 vssd1 vccd1 vccd1 hold284/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 hold295/A vssd1 vssd1 vccd1 vccd1 hold295/X sky130_fd_sc_hd__dlygate4sd3_1
X_09928_ _09928_/A _12614_/A vssd1 vssd1 vccd1 vccd1 _09931_/B sky130_fd_sc_hd__nand2_1
XANTENNA_fanout74_A _07543_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09859_ _12525_/A _09858_/Y _09529_/B vssd1 vssd1 vccd1 vccd1 _09860_/B sky130_fd_sc_hd__a21o_1
X_12870_ _12879_/A _12870_/B vssd1 vssd1 vccd1 vccd1 _12872_/C sky130_fd_sc_hd__nand2_1
X_11821_ _11821_/A _11821_/B vssd1 vssd1 vccd1 vccd1 _11832_/A sky130_fd_sc_hd__xnor2_1
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10077__A2 _10787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12471__B1 _12657_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _11753_/A _11753_/B vssd1 vssd1 vccd1 vccd1 _11853_/A sky130_fd_sc_hd__nand2_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _10703_/A _10703_/B vssd1 vssd1 vccd1 vccd1 _10704_/B sky130_fd_sc_hd__xnor2_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_606 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _12525_/A _11683_/B vssd1 vssd1 vccd1 vccd1 _11683_/X sky130_fd_sc_hd__or2_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13422_ hold113/X _13142_/A _13444_/B1 hold59/X _13430_/C1 vssd1 vssd1 vccd1 vccd1
+ hold139/A sky130_fd_sc_hd__o221a_1
X_10634_ _10572_/A _10572_/B _10570_/X vssd1 vssd1 vccd1 vccd1 _10723_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13353_ _13359_/A hold201/X vssd1 vssd1 vccd1 vccd1 hold202/A sky130_fd_sc_hd__and2_1
XANTENNA__08442__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10565_ _10565_/A _10565_/B vssd1 vssd1 vccd1 vccd1 _10567_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10785__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12304_ _12303_/A _12303_/B _12303_/Y _09506_/X vssd1 vssd1 vccd1 vccd1 _12304_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13284_ _13451_/A _13451_/B _13281_/Y vssd1 vssd1 vccd1 vccd1 _13456_/A sky130_fd_sc_hd__o21ai_1
X_10496_ _10496_/A _10496_/B vssd1 vssd1 vccd1 vccd1 _10497_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_32_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12526__A1 _12525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12235_ _12235_/A _12235_/B _12235_/C vssd1 vssd1 vccd1 vccd1 _12235_/X sky130_fd_sc_hd__and3_1
XANTENNA__07402__B1 _08873_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12166_ _12112_/A _12112_/B _12111_/A vssd1 vssd1 vccd1 vccd1 _12200_/A sky130_fd_sc_hd__o21ai_1
X_11117_ _11562_/A _11117_/B vssd1 vssd1 vccd1 vccd1 _11118_/B sky130_fd_sc_hd__nor2_1
X_12097_ _12187_/B _12097_/B vssd1 vssd1 vccd1 vccd1 _12099_/B sky130_fd_sc_hd__nand2_1
X_11048_ _11048_/A _11048_/B vssd1 vssd1 vccd1 vccd1 _11050_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06947__A _11126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08779__B1_N _08746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12999_ reg1_val[4] _13000_/B vssd1 vssd1 vccd1 vccd1 _12999_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_52_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07210_ _09694_/A _07572_/S _07208_/X vssd1 vssd1 vccd1 vccd1 _07210_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_0_55_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08190_ _09216_/B2 fanout84/X _08580_/B _08868_/B1 vssd1 vssd1 vccd1 vccd1 _08191_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07141_ _09507_/C _09520_/A vssd1 vssd1 vccd1 vccd1 _09505_/B sky130_fd_sc_hd__or2_2
XFILLER_0_6_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07072_ _12740_/A _07071_/X _07060_/Y vssd1 vssd1 vccd1 vccd1 _07072_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10528__B1 _07877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13190__A1 _12189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07974_ _10095_/A _07974_/B vssd1 vssd1 vccd1 vccd1 _07978_/B sky130_fd_sc_hd__xnor2_2
X_09713_ _10600_/S _09712_/X _10601_/C vssd1 vssd1 vccd1 vccd1 _09713_/X sky130_fd_sc_hd__o21a_1
X_06925_ reg1_val[14] _07527_/A vssd1 vssd1 vccd1 vccd1 _06927_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_93_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09644_ _09644_/A _09644_/B vssd1 vssd1 vccd1 vccd1 _09646_/B sky130_fd_sc_hd__xnor2_2
X_06856_ _06856_/A _06856_/B vssd1 vssd1 vccd1 vccd1 _12303_/A sky130_fd_sc_hd__nor2_2
X_09575_ _09575_/A _09575_/B vssd1 vssd1 vccd1 vccd1 _09577_/B sky130_fd_sc_hd__xnor2_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06787_ instruction[41] _06781_/X _06784_/X vssd1 vssd1 vccd1 vccd1 _06886_/A sky130_fd_sc_hd__a21oi_4
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08526_ _08607_/A _08607_/B vssd1 vssd1 vccd1 vccd1 _08608_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_38_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08457_ _08457_/A _08457_/B vssd1 vssd1 vccd1 vccd1 _08516_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08672__A2 _10538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07688__A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07408_ _07377_/A _07377_/B _07410_/A vssd1 vssd1 vccd1 vccd1 _07408_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_108_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08388_ _11072_/A _08388_/B vssd1 vssd1 vccd1 vccd1 _08454_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12756__A1 _13129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07339_ reg1_val[22] _07634_/B _13082_/B _07339_/D vssd1 vssd1 vccd1 vccd1 _12235_/A
+ sky130_fd_sc_hd__or4_1
XANTENNA__08424__A2 _07544_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10350_ _10348_/X _10350_/B vssd1 vssd1 vccd1 vccd1 _10351_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_60_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09009_ _09994_/B _09994_/C vssd1 vssd1 vccd1 vccd1 _10160_/B sky130_fd_sc_hd__nor2_1
X_10281_ _10138_/A _10138_/B _10136_/X vssd1 vssd1 vccd1 vccd1 _10288_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12020_ _12021_/A _12021_/B vssd1 vssd1 vccd1 vccd1 _12110_/B sky130_fd_sc_hd__and2_1
XANTENNA__09924__A2 _10536_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12922_ _12922_/A _12922_/B vssd1 vssd1 vccd1 vccd1 _12937_/B sky130_fd_sc_hd__or2_1
XANTENNA__11495__A1 _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11495__B2 _12103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07362__S _12252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09143__A _10239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12853_ reg1_val[8] curr_PC[8] _12867_/S vssd1 vssd1 vccd1 vccd1 _12855_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_96_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11804_ _11920_/A _11804_/B vssd1 vssd1 vccd1 vccd1 _11805_/B sky130_fd_sc_hd__nor2_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12784_ hold224/A _12750_/X _12374_/A vssd1 vssd1 vccd1 vccd1 _12785_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_29_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _11735_/A _11735_/B vssd1 vssd1 vccd1 vccd1 _11736_/B sky130_fd_sc_hd__and2_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08663__A2 _07492_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11666_ _11226_/X _11665_/A _11857_/A _11664_/X vssd1 vssd1 vccd1 vccd1 _11666_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_0_24_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13405_ _11076_/A _13445_/A2 hold158/X vssd1 vssd1 vccd1 vccd1 _13684_/D sky130_fd_sc_hd__o21a_1
X_10617_ _13015_/A curr_PC[7] vssd1 vssd1 vccd1 vccd1 _10617_/Y sky130_fd_sc_hd__nor2_1
X_11597_ curr_PC[14] curr_PC[15] _11597_/C vssd1 vssd1 vccd1 vccd1 _11794_/C sky130_fd_sc_hd__and3_2
XFILLER_0_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07623__B1 _07699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13336_ hold163/X _13506_/B2 _13506_/A2 hold240/A vssd1 vssd1 vccd1 vccd1 hold164/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10548_ _10391_/A _10686_/A _10548_/C vssd1 vssd1 vccd1 vccd1 _10686_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_106_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13267_ hold73/X hold287/X vssd1 vssd1 vccd1 vccd1 _13267_/X sky130_fd_sc_hd__and2b_1
X_10479_ curr_PC[6] _10480_/B vssd1 vssd1 vccd1 vccd1 _10479_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13172__A1 _13172_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12218_ _12218_/A _12218_/B vssd1 vssd1 vccd1 vccd1 _12218_/Y sky130_fd_sc_hd__nand2_1
X_13198_ _12496_/A _13598_/C hold47/X _13568_/A vssd1 vssd1 vccd1 vccd1 _13635_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12149_ _12311_/B1 _12227_/B hold174/A vssd1 vssd1 vccd1 vccd1 _12151_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12132__C1 _10866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11486__A1 _12760_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07690_ _08951_/A _07690_/B vssd1 vssd1 vccd1 vccd1 _07788_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09360_ _11732_/A fanout83/X fanout79/X _10814_/A1 vssd1 vssd1 vccd1 vccd1 _09361_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08311_ _08311_/A _08311_/B vssd1 vssd1 vccd1 vccd1 _08313_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_47_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09291_ _09414_/A _09291_/B vssd1 vssd1 vccd1 vccd1 _09293_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_74_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_13 instruction[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08242_ _08242_/A _08242_/B vssd1 vssd1 vccd1 vccd1 _08360_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_117_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_24 reg1_val[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 reg1_val[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_46 reg2_val[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_57 reg2_val[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_68 _09910_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08173_ _08173_/A _08173_/B vssd1 vssd1 vccd1 vccd1 _08174_/C sky130_fd_sc_hd__and2_1
XFILLER_0_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_79 reg1_val[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10749__B1 _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout124_A _07366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07020__B _07025_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07124_ instruction[11] _07129_/B vssd1 vssd1 vccd1 vccd1 dest_idx[0] sky130_fd_sc_hd__and2_4
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06968__A2 _06936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07055_ reg1_val[20] _07201_/A vssd1 vssd1 vccd1 vccd1 _07055_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10662__A _11719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07447__S _11913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07957_ _07958_/A _07958_/B vssd1 vssd1 vccd1 vccd1 _07957_/X sky130_fd_sc_hd__and2_1
X_06908_ reg1_val[16] _07297_/A vssd1 vssd1 vccd1 vccd1 _11772_/B sky130_fd_sc_hd__nand2_1
X_07888_ _10239_/A _07888_/B vssd1 vssd1 vccd1 vccd1 _07897_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07145__A2 _12578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09627_ _09627_/A _09627_/B vssd1 vssd1 vccd1 vccd1 _09630_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_69_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06839_ _06840_/A _06840_/B vssd1 vssd1 vccd1 vccd1 _06849_/C sky130_fd_sc_hd__and2_1
XFILLER_0_78_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09558_ _09559_/A _09559_/B _09559_/C vssd1 vssd1 vccd1 vccd1 _09811_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout37_A _07368_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08509_ _08507_/A _08507_/B _08575_/A vssd1 vssd1 vccd1 vccd1 _08518_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__10437__C1 _10631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09489_ reg1_val[4] reg1_val[27] _09493_/S vssd1 vssd1 vccd1 vccd1 _09489_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_92_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11520_ _11520_/A _11520_/B vssd1 vssd1 vccd1 vccd1 _11522_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_25_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08307__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout3_A fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07211__A _07230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11451_ _11221_/X _11339_/X _11341_/B vssd1 vssd1 vccd1 vccd1 _11451_/Y sky130_fd_sc_hd__a21oi_2
X_10402_ _07299_/Y fanout20/X fanout18/X _10814_/A1 vssd1 vssd1 vccd1 vccd1 _10403_/B
+ sky130_fd_sc_hd__o22a_2
X_11382_ curr_PC[12] curr_PC[13] _11382_/C vssd1 vssd1 vccd1 vccd1 _11597_/C sky130_fd_sc_hd__and3_1
XFILLER_0_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13121_ _13121_/A _13121_/B vssd1 vssd1 vccd1 vccd1 _13121_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10333_ reg1_val[5] curr_PC[5] vssd1 vssd1 vccd1 vccd1 _10334_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13154__A1 _10104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ _13057_/B _13052_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[13] sky130_fd_sc_hd__and2_4
X_10264_ _10271_/A vssd1 vssd1 vccd1 vccd1 _10264_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_103_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11704__A2 _09146_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12003_ _12417_/A _12003_/B vssd1 vssd1 vccd1 vccd1 _12004_/A sky130_fd_sc_hd__xnor2_1
X_10195_ _09860_/A _10180_/Y _10181_/X _09529_/B _10194_/X vssd1 vssd1 vccd1 vccd1
+ _10195_/Y sky130_fd_sc_hd__o221ai_2
XANTENNA__10912__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12665__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06928__C _13054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12905_ _12912_/A _12905_/B vssd1 vssd1 vccd1 vccd1 _12907_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_124_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12836_ _12837_/A _12837_/B _12837_/C vssd1 vssd1 vccd1 vccd1 _12844_/B sky130_fd_sc_hd__a21o_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10691__A2 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _12574_/B _12682_/D _12765_/Y _12766_/X vssd1 vssd1 vccd1 vccd1 _12768_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06944__B _06980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11718_ fanout54/X fanout34/X fanout32/X _12268_/A vssd1 vssd1 vccd1 vccd1 _11719_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_83_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12698_ reg1_val[28] reg1_val[29] _12698_/C vssd1 vssd1 vccd1 vccd1 _12782_/C sky130_fd_sc_hd__and3_1
XFILLER_0_84_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11649_ _11540_/A _11539_/B _11537_/X vssd1 vssd1 vccd1 vccd1 _11650_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_114_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13393__A1 _10239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13319_ _13459_/A _13319_/B vssd1 vssd1 vccd1 vccd1 _13641_/D sky130_fd_sc_hd__and2_1
XFILLER_0_122_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07267__S _07572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08860_ _08860_/A _08860_/B vssd1 vssd1 vccd1 vccd1 _08861_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09482__S _09839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07811_ _07811_/A _07811_/B vssd1 vssd1 vccd1 vccd1 _07813_/B sky130_fd_sc_hd__xnor2_1
X_08791_ _08791_/A _08791_/B vssd1 vssd1 vccd1 vccd1 _08793_/B sky130_fd_sc_hd__xnor2_1
X_07742_ _07819_/A _07819_/B vssd1 vssd1 vccd1 vccd1 _07830_/A sky130_fd_sc_hd__nor2_1
X_07673_ _07451_/X fanout24/X _08486_/B _09173_/B2 vssd1 vssd1 vccd1 vccd1 _07674_/B
+ sky130_fd_sc_hd__o22a_1
X_09412_ _09223_/A _09223_/B _09224_/X vssd1 vssd1 vccd1 vccd1 _09417_/A sky130_fd_sc_hd__o21bai_4
XANTENNA__07015__B _10456_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12408__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09343_ _09246_/A _09246_/B _09249_/A vssd1 vssd1 vccd1 vccd1 _09347_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_90_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06854__B _07230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09274_ _09275_/A _09275_/B vssd1 vssd1 vccd1 vccd1 _09274_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_90_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08225_ _08225_/A _08225_/B vssd1 vssd1 vccd1 vccd1 _08300_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08156_ _08156_/A _08156_/B vssd1 vssd1 vccd1 vccd1 _08158_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11395__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07107_ _07135_/S dest_pred_val _12406_/B1 vssd1 vssd1 vccd1 vccd1 take_branch sky130_fd_sc_hd__a21o_4
X_08087_ _08112_/A _08112_/B vssd1 vssd1 vccd1 vccd1 _08160_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_3_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07038_ _06976_/Y _07037_/X _10736_/A vssd1 vssd1 vccd1 vccd1 _10867_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08012__B1 _08246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12811__S _12825_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08797__A _09659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11698__B2 _10866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__B1 _10235_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ _08988_/A _08988_/B _08988_/C _09081_/A _09077_/A vssd1 vssd1 vccd1 vccd1
+ _08990_/B sky130_fd_sc_hd__a311o_1
XANTENNA__13439__A2 _13598_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08315__A1 _08866_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08315__B2 _09216_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07206__A _10239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10951_ _10952_/A _10952_/B vssd1 vssd1 vccd1 vccd1 _11029_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08866__A2 _08866_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10673__A2 _10787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13670_ _13735_/CLK hold199/X vssd1 vssd1 vccd1 vccd1 hold197/A sky130_fd_sc_hd__dfxtp_1
X_10882_ hold163/A hold180/A _10882_/C vssd1 vssd1 vccd1 vccd1 _11004_/B sky130_fd_sc_hd__or3_1
XFILLER_0_78_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12621_ _12621_/A _12677_/A _12621_/C vssd1 vssd1 vccd1 vccd1 _12677_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_66_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07826__B1 _08395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12552_ _12552_/A _12552_/B vssd1 vssd1 vccd1 vccd1 _12555_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_65_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11503_ _11503_/A _11503_/B vssd1 vssd1 vccd1 vccd1 _11525_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_80_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12782__A _13129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12483_ fanout12/X _12667_/A _09145_/Y fanout16/X vssd1 vssd1 vccd1 vccd1 _12484_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12178__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11434_ _11310_/A _11310_/B _11308_/A vssd1 vssd1 vccd1 vccd1 _11436_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_22_724 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11398__A _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11365_ _11362_/X _11364_/X _12225_/A vssd1 vssd1 vccd1 vccd1 _11365_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_104_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13104_ _13105_/A _13105_/B vssd1 vssd1 vccd1 vccd1 _13112_/A sky130_fd_sc_hd__nand2b_1
X_10316_ _09672_/X _09683_/X _10600_/S vssd1 vssd1 vccd1 vccd1 _10316_/X sky130_fd_sc_hd__mux2_1
X_11296_ _12557_/A fanout29/X fanout27/X _12557_/B vssd1 vssd1 vccd1 vccd1 _11297_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ reg1_val[11] _13036_/B vssd1 vssd1 vccd1 vccd1 _13037_/A sky130_fd_sc_hd__or2_1
X_10247_ fanout51/X fanout68/X fanout66/X fanout44/X vssd1 vssd1 vccd1 vccd1 _10248_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10178_ _10178_/A vssd1 vssd1 vccd1 vccd1 _10178_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_89_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08306__A1 _08806_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08306__B2 _08806_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07116__A _13141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12819_ _12995_/B _12820_/B vssd1 vssd1 vccd1 vccd1 _12830_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09267__C1 _13129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08490__B1 _08778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08010_ _07347_/X fanout28/X _08395_/B _09216_/B2 vssd1 vssd1 vccd1 vccd1 _08011_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09477__S _09493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12169__A2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09961_ _09961_/A _09961_/B vssd1 vssd1 vccd1 vccd1 _09963_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08912_ _08920_/A _08916_/B vssd1 vssd1 vccd1 vccd1 _08912_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09892_ _09893_/A _09893_/B vssd1 vssd1 vccd1 vccd1 _09892_/Y sky130_fd_sc_hd__nand2_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12341__A2 _07891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08843_ _08843_/A _08843_/B _08843_/C vssd1 vssd1 vccd1 vccd1 _08844_/B sky130_fd_sc_hd__or3_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10352__A1 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout191_A _12796_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10352__B2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08774_ _08774_/A _08774_/B vssd1 vssd1 vccd1 vccd1 _08804_/B sky130_fd_sc_hd__xor2_1
X_07725_ _09173_/B2 fanout83/X fanout79/X _07471_/Y vssd1 vssd1 vccd1 vccd1 _07726_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13462__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07656_ _07656_/A _07656_/B vssd1 vssd1 vccd1 vccd1 _07658_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06865__A _06886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07460__S _07572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09241__A _10944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07587_ _07588_/A _07588_/B vssd1 vssd1 vccd1 vccd1 _07948_/B sky130_fd_sc_hd__and2b_1
X_09326_ _09311_/A _09311_/B _09309_/X vssd1 vssd1 vccd1 vccd1 _09426_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_63_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11604__A1 _12557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11604__B2 _07597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09257_ _08271_/A _10536_/A2 fanout6/X _12982_/A vssd1 vssd1 vccd1 vccd1 _09258_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08481__B1 _09173_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08208_ _10236_/A _08208_/B vssd1 vssd1 vccd1 vccd1 _08214_/A sky130_fd_sc_hd__xnor2_2
X_09188_ _07873_/A _07872_/B _07872_/A vssd1 vssd1 vccd1 vccd1 _09193_/A sky130_fd_sc_hd__o21bai_4
XANTENNA__11368__B1 _12533_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08139_ _10078_/A _08139_/B vssd1 vssd1 vccd1 vccd1 _08176_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11150_ _11114_/A _11114_/B _10984_/X vssd1 vssd1 vccd1 vccd1 _11150_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_31_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10591__A1 _12515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10101_ _10102_/A _10102_/B vssd1 vssd1 vccd1 vccd1 _10103_/A sky130_fd_sc_hd__or2_1
X_11081_ _11082_/A _11082_/B vssd1 vssd1 vccd1 vccd1 _11083_/A sky130_fd_sc_hd__or2_1
XFILLER_0_101_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10032_ _12314_/A _10031_/X hold264/A vssd1 vssd1 vccd1 vccd1 _10032_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__08320__A _11286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09850__S _10007_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11983_ _10866_/B _11956_/X _11957_/Y _11982_/Y _11955_/X vssd1 vssd1 vccd1 vccd1
+ _11983_/X sky130_fd_sc_hd__o311a_1
XFILLER_0_98_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_4_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13719_/CLK sky130_fd_sc_hd__clkbuf_8
X_13722_ _13725_/CLK _13722_/D vssd1 vssd1 vccd1 vccd1 hold257/A sky130_fd_sc_hd__dfxtp_1
X_10934_ _10934_/A fanout6/X vssd1 vssd1 vccd1 vccd1 _10934_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12496__B _12666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13653_ _13659_/CLK _13653_/D vssd1 vssd1 vccd1 vccd1 hold214/A sky130_fd_sc_hd__dfxtp_1
X_10865_ _11562_/A _10864_/B _10864_/C vssd1 vssd1 vccd1 vccd1 _10866_/A sky130_fd_sc_hd__o21a_1
XANTENNA__10297__A _10577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12604_ _09529_/B _12591_/X _12597_/X _12603_/X vssd1 vssd1 vccd1 vccd1 _12604_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13584_ hold233/X _13584_/B vssd1 vssd1 vccd1 vccd1 _13584_/X sky130_fd_sc_hd__and2_1
XFILLER_0_54_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10796_ _10796_/A _10796_/B vssd1 vssd1 vccd1 vccd1 _10798_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12535_ reg1_val[26] _11688_/B _07252_/C _10889_/B vssd1 vssd1 vccd1 vccd1 _12535_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_121_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11071__A2 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12466_ hold278/A _12786_/B1 _12527_/B _12465_/Y _12748_/B1 vssd1 vssd1 vccd1 vccd1
+ _12475_/B sky130_fd_sc_hd__a311o_1
XFILLER_0_22_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11417_ _11417_/A _11417_/B vssd1 vssd1 vccd1 vccd1 _11418_/B sky130_fd_sc_hd__and2_1
XFILLER_0_111_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12397_ _06847_/A _09520_/X _12396_/X vssd1 vssd1 vccd1 vccd1 _12397_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_111_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07578__A2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11348_ _11864_/A _11348_/B _11600_/B vssd1 vssd1 vccd1 vccd1 _11348_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__12451__S _12515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11279_ _11279_/A _11279_/B vssd1 vssd1 vccd1 vccd1 _11290_/A sky130_fd_sc_hd__xor2_1
XANTENNA__08527__A1 _08821_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08527__B2 _08821_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13018_ _13017_/A _13014_/Y _13016_/B vssd1 vssd1 vccd1 vccd1 _13022_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_55_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07750__A2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07510_ _07517_/A _07517_/B vssd1 vssd1 vccd1 vccd1 _07510_/Y sky130_fd_sc_hd__nor2_1
X_08490_ _09216_/B2 _10538_/A _08778_/B _08868_/B1 vssd1 vssd1 vccd1 vccd1 _08491_/B
+ sky130_fd_sc_hd__o22a_1
X_07441_ _11884_/A _11884_/B _07637_/B vssd1 vssd1 vccd1 vccd1 _07445_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout19 _07493_/Y vssd1 vssd1 vccd1 vccd1 _08246_/B sky130_fd_sc_hd__buf_8
XFILLER_0_57_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07372_ reg1_val[24] reg1_val[25] vssd1 vssd1 vccd1 vccd1 _07377_/C sky130_fd_sc_hd__nor2_1
XANTENNA__11598__B1 _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09111_ _09111_/A _09111_/B vssd1 vssd1 vccd1 vccd1 _09113_/C sky130_fd_sc_hd__or2_1
XFILLER_0_127_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09042_ _08786_/A _08786_/B _08726_/A _08726_/B vssd1 vssd1 vccd1 vccd1 _09042_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11770__B1 _11866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13457__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09944_ _09944_/A _09944_/B vssd1 vssd1 vccd1 vccd1 _09945_/B sky130_fd_sc_hd__or2_1
XFILLER_0_0_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09236__A _10095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13511__B2 _13542_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09875_ _09866_/Y _09867_/X _09874_/X vssd1 vssd1 vccd1 vccd1 _09875_/Y sky130_fd_sc_hd__o21ai_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _08866_/B2 _09216_/B2 _08868_/B1 _08950_/B vssd1 vssd1 vccd1 vccd1 _08827_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09670__S _09703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08757_ _08762_/A _08755_/X _08743_/X vssd1 vssd1 vccd1 vccd1 _08784_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_68_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07708_ _07708_/A _07708_/B vssd1 vssd1 vccd1 vccd1 _07709_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_95_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08688_ _08728_/A _08728_/B vssd1 vssd1 vccd1 vccd1 _08729_/A sky130_fd_sc_hd__and2_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07639_ _12417_/A _07639_/B vssd1 vssd1 vccd1 vccd1 _12617_/A sky130_fd_sc_hd__nor2_1
XANTENNA__13205__B _13207_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10650_ _07306_/X fanout6/X _10649_/Y _10537_/A vssd1 vssd1 vccd1 vccd1 _10652_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11589__B1 _11588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09309_ _09310_/A _09310_/B vssd1 vssd1 vccd1 vccd1 _09309_/X sky130_fd_sc_hd__and2_1
XANTENNA__07257__A1 _07594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12250__A1 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10581_ _10300_/Y _10576_/Y _10580_/Y vssd1 vssd1 vccd1 vccd1 _10581_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12250__B2 _07699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12320_ _12710_/B2 _10744_/X _10758_/X _12537_/B2 _12319_/X vssd1 vssd1 vccd1 vccd1
+ _12320_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10541__A_N _09575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12002__A1 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12251_ _12417_/A _12251_/B vssd1 vssd1 vccd1 vccd1 _12253_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12002__B2 _12557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11202_ _11202_/A _11202_/B vssd1 vssd1 vccd1 vccd1 _11203_/B sky130_fd_sc_hd__or2_1
XANTENNA__12553__A2 _09145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12182_ _12182_/A _12182_/B vssd1 vssd1 vccd1 vccd1 _12197_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11133_ _13651_/Q _11248_/C vssd1 vssd1 vccd1 vccd1 _11133_/X sky130_fd_sc_hd__or2_1
X_11064_ _11064_/A _11064_/B vssd1 vssd1 vccd1 vccd1 _11065_/B sky130_fd_sc_hd__and2_1
X_10015_ _10016_/B _10016_/C _10016_/A vssd1 vssd1 vccd1 vccd1 _10017_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11966_ _11874_/A _11876_/B _11874_/B vssd1 vssd1 vccd1 vccd1 _11967_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_58_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06936__C _13048_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07496__A1 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10917_ _10917_/A _10917_/B vssd1 vssd1 vccd1 vccd1 _10929_/A sky130_fd_sc_hd__xnor2_1
X_13705_ _13705_/CLK _13705_/D vssd1 vssd1 vccd1 vccd1 hold245/A sky130_fd_sc_hd__dfxtp_2
XANTENNA__07496__B2 _09885_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11292__A2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11897_ _11843_/A _11843_/B _11844_/X vssd1 vssd1 vccd1 vccd1 _11942_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_128_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13636_ _13739_/CLK _13636_/D vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__dfxtp_1
X_10848_ _10849_/B _10849_/A vssd1 vssd1 vccd1 vccd1 _10976_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_128_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08445__B1 _08704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13567_ hold273/X _13584_/B _13566_/X _13599_/D vssd1 vssd1 vccd1 vccd1 hold274/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10779_ _10780_/A _10780_/B _10780_/C vssd1 vssd1 vccd1 vccd1 _10962_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__06952__B _06980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07799__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12518_ _12130_/A _09082_/X _09087_/X vssd1 vssd1 vccd1 vccd1 _12518_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__12792__A2 _07398_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13498_ _13259_/X _13498_/B vssd1 vssd1 vccd1 vccd1 _13499_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__12529__C1 _12748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12449_ _12480_/B _12447_/X _12448_/Y vssd1 vssd1 vccd1 vccd1 _12476_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08748__A1 _07238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08748__B2 _07239_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout209 _09381_/A vssd1 vssd1 vccd1 vccd1 _09671_/S sky130_fd_sc_hd__buf_4
X_07990_ _08071_/A _07988_/X _07985_/X vssd1 vssd1 vccd1 vccd1 _08092_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_66_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07971__A2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06941_ reg1_val[12] _07188_/B vssd1 vssd1 vccd1 vccd1 _06943_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11504__B1 fanout5/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09173__A1 _10049_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12701__C1 _09529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09173__B2 _09173_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09660_ _09660_/A _09660_/B vssd1 vssd1 vccd1 vccd1 _09660_/Y sky130_fd_sc_hd__xnor2_1
X_06872_ reg2_val[21] _06873_/B1 _06872_/B1 _06871_/Y vssd1 vssd1 vccd1 vccd1 _07201_/B
+ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__08895__A _10236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09490__S _09493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07723__A2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08611_ _08658_/A _08658_/B vssd1 vssd1 vccd1 vccd1 _08659_/A sky130_fd_sc_hd__nor2_1
X_09591_ _09591_/A _09591_/B vssd1 vssd1 vccd1 vccd1 _09599_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08542_ _08806_/B1 _07492_/Y _07556_/Y _08806_/A2 vssd1 vssd1 vccd1 vccd1 _08543_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10649__B fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07304__A _10095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08473_ _08473_/A _08473_/B vssd1 vssd1 vccd1 vccd1 _08475_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__13025__B _13025_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout154_A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07424_ _12421_/A _07424_/B vssd1 vssd1 vccd1 vccd1 _07652_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07355_ _07377_/A _07337_/B _07334_/D _07357_/A vssd1 vssd1 vccd1 vccd1 _12235_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11035__A2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12232__A1 _12314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07286_ _07521_/A _07213_/A _07201_/A vssd1 vssd1 vccd1 vccd1 _08197_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_31_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08135__A _08746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09025_ _09025_/A _09025_/B vssd1 vssd1 vccd1 vccd1 _10988_/A sky130_fd_sc_hd__or2_1
XFILLER_0_60_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07974__A _10095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09665__S _10004_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09936__B1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold230 hold230/A vssd1 vssd1 vccd1 vccd1 hold230/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 hold241/A vssd1 vssd1 vccd1 vccd1 hold241/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold252 hold252/A vssd1 vssd1 vccd1 vccd1 hold252/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 hold263/A vssd1 vssd1 vccd1 vccd1 hold263/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11496__A _11719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold274 hold274/A vssd1 vssd1 vccd1 vccd1 hold274/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 hold285/A vssd1 vssd1 vccd1 vccd1 hold285/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06907__A2_N _06906_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold296 hold296/A vssd1 vssd1 vccd1 vccd1 hold296/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09927_ _11076_/A _09927_/B vssd1 vssd1 vccd1 vccd1 _09932_/A sky130_fd_sc_hd__xnor2_1
X_09858_ _09858_/A _09858_/B vssd1 vssd1 vccd1 vccd1 _09858_/Y sky130_fd_sc_hd__xnor2_2
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08809_ _10236_/A _08809_/B vssd1 vssd1 vccd1 vccd1 _08845_/B sky130_fd_sc_hd__xnor2_1
X_09789_ _09789_/A _09789_/B vssd1 vssd1 vccd1 vccd1 _09806_/A sky130_fd_sc_hd__xor2_1
X_11820_ _11929_/B _11820_/B vssd1 vssd1 vccd1 vccd1 _11821_/B sky130_fd_sc_hd__or2_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _11751_/A _11751_/B vssd1 vssd1 vccd1 vccd1 _11753_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08675__B1 _08704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10077__A3 _10787_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09872__C1 _09871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10702_ _10702_/A _10702_/B vssd1 vssd1 vccd1 vccd1 _10703_/B sky130_fd_sc_hd__xnor2_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _11682_/A _11682_/B vssd1 vssd1 vccd1 vccd1 _11682_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13421_ _11913_/A _13445_/A2 hold114/X vssd1 vssd1 vccd1 vccd1 hold115/A sky130_fd_sc_hd__o21a_1
X_10633_ _10155_/C _10631_/X _10632_/X _10630_/Y vssd1 vssd1 vccd1 vccd1 _10724_/A
+ sky130_fd_sc_hd__o211a_4
XFILLER_0_63_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13352_ hold231/A _13506_/B2 _13506_/A2 hold200/X vssd1 vssd1 vccd1 vccd1 hold201/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10564_ _10564_/A _10564_/B vssd1 vssd1 vccd1 vccd1 _10565_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_91_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10785__A1 _10538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10785__B2 _08778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12303_ _12303_/A _12303_/B vssd1 vssd1 vccd1 vccd1 _12303_/Y sky130_fd_sc_hd__nand2_1
X_13283_ _13704_/Q hold13/X vssd1 vssd1 vccd1 vccd1 _13451_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_23_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10495_ _10495_/A _10495_/B vssd1 vssd1 vccd1 vccd1 _10496_/B sky130_fd_sc_hd__or2_1
XFILLER_0_51_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12234_ _12234_/A _12234_/B vssd1 vssd1 vccd1 vccd1 _12241_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07402__A1 _09381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07402__B2 _07699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12165_ _11601_/X _12373_/A vssd1 vssd1 vccd1 vccd1 _12165_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_102_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11116_ _11115_/A _11115_/B _11955_/A vssd1 vssd1 vccd1 vccd1 _11116_/Y sky130_fd_sc_hd__a21oi_1
X_12096_ _12096_/A _12096_/B vssd1 vssd1 vccd1 vccd1 _12097_/B sky130_fd_sc_hd__or2_1
XFILLER_0_127_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13683__CLK _13701_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11047_ _11047_/A _11825_/A vssd1 vssd1 vccd1 vccd1 _11048_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09604__A _09604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12998_ _12997_/A _12994_/Y _12996_/B vssd1 vssd1 vccd1 vccd1 _13002_/A sky130_fd_sc_hd__o21a_2
XANTENNA_wire122_A wire122/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11949_ _11760_/X _12125_/B _11947_/A vssd1 vssd1 vccd1 vccd1 _11949_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13619_ _13719_/CLK _13619_/D vssd1 vssd1 vccd1 vccd1 hold105/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07140_ _09524_/A _13748_/A vssd1 vssd1 vccd1 vccd1 _09520_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_42_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07071_ _12693_/A _07070_/X _07061_/Y vssd1 vssd1 vccd1 vccd1 _07071_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_2_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09485__S _09839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10528__B2 _10915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13190__A2 _13196_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07973_ _10235_/B2 _11732_/A fanout70/X _08873_/A2 vssd1 vssd1 vccd1 vccd1 _07974_/B
+ sky130_fd_sc_hd__o22a_1
X_09712_ _09484_/X _09536_/B _10004_/S vssd1 vssd1 vccd1 vccd1 _09712_/X sky130_fd_sc_hd__mux2_1
X_06924_ reg1_val[14] _07527_/A vssd1 vssd1 vccd1 vccd1 _06927_/A sky130_fd_sc_hd__or2_1
XANTENNA__07018__B _07110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12150__B1 _12533_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09643_ _09417_/A _09417_/B _09415_/X vssd1 vssd1 vccd1 vccd1 _09644_/B sky130_fd_sc_hd__a21oi_4
X_06855_ _07334_/B _07230_/A vssd1 vssd1 vccd1 vccd1 _06856_/B sky130_fd_sc_hd__and2_1
XANTENNA__06857__B _12981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09574_ fanout53/X fanout68/X fanout66/X fanout47/X vssd1 vssd1 vccd1 vccd1 _09575_/B
+ sky130_fd_sc_hd__o22a_1
X_06786_ instruction[41] _06781_/X _06784_/X vssd1 vssd1 vccd1 vccd1 _06989_/B sky130_fd_sc_hd__a21o_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08525_ _09591_/A _08525_/B vssd1 vssd1 vccd1 vccd1 _08607_/B sky130_fd_sc_hd__xnor2_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11256__A2 _12793_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12875__A _13036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13470__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08456_ _08456_/A _08456_/B vssd1 vssd1 vccd1 vccd1 _08458_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_65_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07407_ _09496_/S _07407_/B vssd1 vssd1 vccd1 vccd1 _09748_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_46_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08387_ _10225_/A _07541_/X _07545_/Y _07556_/Y vssd1 vssd1 vccd1 vccd1 _08388_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12756__A2 _11688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07338_ _07634_/B _13082_/B _07339_/D vssd1 vssd1 vccd1 vccd1 _07351_/A sky130_fd_sc_hd__or3_1
XFILLER_0_33_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07269_ reg1_val[4] reg1_val[5] _07265_/D reg1_val[6] vssd1 vssd1 vccd1 vccd1 _07270_/B
+ sky130_fd_sc_hd__o31ai_1
X_09008_ _09008_/A _09008_/B vssd1 vssd1 vccd1 vccd1 _09994_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__13166__C1 _13543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10280_ _10131_/A _10131_/B _10129_/X vssd1 vssd1 vccd1 vccd1 _10290_/A sky130_fd_sc_hd__a21o_1
XANTENNA__11954__A _12695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12921_ _12938_/A _12921_/B vssd1 vssd1 vccd1 vccd1 _12937_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_88_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11495__A2 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12852_ _12858_/B _12852_/B vssd1 vssd1 vccd1 vccd1 new_PC[7] sky130_fd_sc_hd__and2_4
XFILLER_0_87_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11803_ _11920_/A _11804_/B vssd1 vssd1 vccd1 vccd1 _11805_/A sky130_fd_sc_hd__and2_1
X_12783_ _12783_/A _12783_/B vssd1 vssd1 vccd1 vccd1 _12783_/X sky130_fd_sc_hd__xor2_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11734_ _11735_/A _11735_/B vssd1 vssd1 vccd1 vccd1 _11736_/A sky130_fd_sc_hd__nor2_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11665_ _11665_/A _11857_/A vssd1 vssd1 vccd1 vccd1 _11665_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10207__B1 _07471_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10616_ _10473_/A _10470_/Y _10472_/B vssd1 vssd1 vccd1 vccd1 _10620_/A sky130_fd_sc_hd__o21a_1
X_13404_ hold157/X _13416_/A2 _13420_/B1 hold120/X _13383_/A vssd1 vssd1 vccd1 vccd1
+ hold158/A sky130_fd_sc_hd__o221a_1
X_11596_ _07152_/X _11595_/X _07544_/A _10889_/B vssd1 vssd1 vccd1 vccd1 _11596_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_52_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10758__A1 _10603_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13335_ _13359_/A hold181/X vssd1 vssd1 vccd1 vccd1 _13649_/D sky130_fd_sc_hd__and2_1
XANTENNA__07623__A1 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10547_ _10546_/B _10546_/C _10546_/A vssd1 vssd1 vccd1 vccd1 _10548_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_24_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07623__B2 _13149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13266_ hold276/X hold68/X vssd1 vssd1 vccd1 vccd1 _13483_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_122_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10478_ _10442_/X _10443_/Y _10445_/Y _11866_/A _10477_/X vssd1 vssd1 vccd1 vccd1
+ _10478_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_32_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12217_ _12215_/X _12216_/X _12578_/A vssd1 vssd1 vccd1 vccd1 _12218_/B sky130_fd_sc_hd__mux2_1
XANTENNA__13172__A2 _13194_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13197_ hold46/X _13207_/B vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__or2_1
XFILLER_0_20_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12148_ hold212/A _13660_/Q _12148_/C vssd1 vssd1 vccd1 vccd1 _12227_/B sky130_fd_sc_hd__or3_1
X_12079_ _12557_/A fanout35/X _07699_/B _12557_/B vssd1 vssd1 vccd1 vccd1 _12080_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11885__A2_N _11688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11891__C1 _11890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12695__A _12695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08310_ _08311_/A _08311_/B vssd1 vssd1 vccd1 vccd1 _08310_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_87_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09290_ _09289_/A _09289_/C _09289_/B vssd1 vssd1 vccd1 vccd1 _09291_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_87_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08241_ _08242_/A _08242_/B vssd1 vssd1 vccd1 vccd1 _08241_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_14 instruction[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_25 reg1_val[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_36 reg1_val[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_47 reg2_val[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08172_ _08172_/A _08172_/B vssd1 vssd1 vccd1 vccd1 _08173_/B sky130_fd_sc_hd__or2_1
XANTENNA__07301__B _07535_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_58 reg2_val[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_69 _09706_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07123_ _07123_/A _07123_/B vssd1 vssd1 vccd1 vccd1 _07129_/B sky130_fd_sc_hd__or2_2
XFILLER_0_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout117_A _11508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06968__A3 _13025_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13148__C1 _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07054_ reg1_val[21] _07201_/B vssd1 vssd1 vccd1 vccd1 _07054_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_30_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07956_ _07956_/A _07956_/B vssd1 vssd1 vccd1 vccd1 _07958_/B sky130_fd_sc_hd__xnor2_4
X_06907_ _06905_/Y _06906_/B1 _06980_/B reg2_val[16] vssd1 vssd1 vccd1 vccd1 _06911_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_07887_ _08821_/A1 fanout49/X fanout45/X _08821_/B2 vssd1 vssd1 vccd1 vccd1 _07888_/B
+ sky130_fd_sc_hd__o22a_1
X_09626_ _09624_/X _09626_/B vssd1 vssd1 vccd1 vccd1 _09627_/B sky130_fd_sc_hd__nand2b_1
X_06838_ _07392_/A _07217_/A vssd1 vssd1 vccd1 vccd1 _06840_/B sky130_fd_sc_hd__nand2_1
X_09557_ _09557_/A _09557_/B vssd1 vssd1 vccd1 vccd1 _09559_/C sky130_fd_sc_hd__xor2_1
X_06769_ instruction[21] instruction[14] _07135_/S vssd1 vssd1 vccd1 vccd1 reg1_idx[3]
+ sky130_fd_sc_hd__mux2_8
X_08508_ _08574_/A _08574_/B vssd1 vssd1 vccd1 vccd1 _08575_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_77_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07699__A _09381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09488_ _09484_/X _09487_/X _10007_/S vssd1 vssd1 vccd1 vccd1 _09488_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_65_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08439_ _08438_/A _08505_/A _08451_/A vssd1 vssd1 vccd1 vccd1 _08439_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11450_ _11450_/A _11450_/B vssd1 vssd1 vccd1 vccd1 _11663_/A sky130_fd_sc_hd__or2_4
XFILLER_0_46_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10401_ _12253_/A _10401_/B vssd1 vssd1 vccd1 vccd1 _10410_/A sky130_fd_sc_hd__xnor2_4
X_11381_ _10730_/B _11348_/Y _11349_/X _11352_/Y _11380_/Y vssd1 vssd1 vccd1 vccd1
+ _11381_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_116_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13120_ _13120_/A _13120_/B vssd1 vssd1 vccd1 vccd1 _13123_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_61_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10332_ reg1_val[5] curr_PC[5] vssd1 vssd1 vccd1 vccd1 _10332_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13051_ _13051_/A _13051_/B _13051_/C vssd1 vssd1 vccd1 vccd1 _13052_/B sky130_fd_sc_hd__nand3_1
XANTENNA__13154__A2 _13194_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10263_ _10263_/A _10263_/B vssd1 vssd1 vccd1 vccd1 _10271_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07369__B1 _07366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12002_ fanout50/X fanout34/X fanout32/X _12557_/A vssd1 vssd1 vccd1 vccd1 _12003_/B
+ sky130_fd_sc_hd__o22a_1
X_10194_ _09839_/A _10193_/Y _10191_/X _10184_/X vssd1 vssd1 vccd1 vccd1 _10194_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10912__A1 _07477_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10912__B2 _07472_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12665__A1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12665__B2 _09145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12904_ _13059_/B _12904_/B vssd1 vssd1 vccd1 vccd1 _12905_/B sky130_fd_sc_hd__or2_1
XFILLER_0_69_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ _12844_/A _12835_/B vssd1 vssd1 vccd1 vccd1 _12837_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _12731_/A _12725_/Y _12765_/Y _12683_/X _12727_/B vssd1 vssd1 vccd1 vccd1
+ _12766_/X sky130_fd_sc_hd__a221o_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11717_ _11717_/A vssd1 vssd1 vccd1 vccd1 _11724_/A sky130_fd_sc_hd__inv_2
X_12697_ _09321_/A _12695_/X _12696_/Y vssd1 vssd1 vccd1 vccd1 _12714_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_71_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11648_ _11648_/A _11648_/B vssd1 vssd1 vccd1 vccd1 _11650_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_24_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11579_ hold300/A hold289/A _11579_/C vssd1 vssd1 vccd1 vccd1 _11881_/D sky130_fd_sc_hd__or3_2
XANTENNA__06960__B _06980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13318_ hold188/X _13450_/B fanout1/X _13463_/B2 vssd1 vssd1 vccd1 vccd1 _13319_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13249_ hold296/A hold126/X vssd1 vssd1 vccd1 vccd1 _13250_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_58_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07810_ _07798_/A _07798_/B _08022_/A vssd1 vssd1 vccd1 vccd1 _07838_/A sky130_fd_sc_hd__o21a_1
X_08790_ _08790_/A _08790_/B vssd1 vssd1 vccd1 vccd1 _08793_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_74_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07741_ _07741_/A _07741_/B vssd1 vssd1 vccd1 vccd1 _07819_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11459__A2 _11458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07672_ _07672_/A _07672_/B vssd1 vssd1 vccd1 vccd1 _07683_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09411_ _09297_/A _09297_/B _09296_/A vssd1 vssd1 vccd1 vccd1 _09421_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12408__A1 _07257_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12408__B2 _12496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09342_ _09342_/A _09342_/B vssd1 vssd1 vccd1 vccd1 _09410_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_59_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09511__B _13744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09273_ _11731_/A _09273_/B vssd1 vssd1 vccd1 vccd1 _09275_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_7_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08224_ _08224_/A _08224_/B vssd1 vssd1 vccd1 vccd1 _08226_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_28_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08155_ _08155_/A _08155_/B vssd1 vssd1 vccd1 vccd1 _08158_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11395__A1 _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07106_ instruction[1] _07123_/A vssd1 vssd1 vccd1 vccd1 _07106_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11395__B2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08086_ _10263_/A _08086_/B vssd1 vssd1 vccd1 vccd1 _08112_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07037_ _10588_/B _10588_/C _10592_/A vssd1 vssd1 vccd1 vccd1 _07037_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_30_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09673__S _09674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08012__A1 _13149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07982__A _09948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08012__B2 _08923_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__A1 _10235_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__B2 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08988_ _08988_/A _08988_/B _08988_/C vssd1 vssd1 vccd1 vccd1 _09074_/B sky130_fd_sc_hd__and3_1
X_07939_ _07940_/A _07940_/B _07940_/C vssd1 vssd1 vccd1 vccd1 _09190_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__08315__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10950_ _10950_/A _10950_/B vssd1 vssd1 vccd1 vccd1 _10952_/B sky130_fd_sc_hd__xnor2_1
X_09609_ _09609_/A _09609_/B vssd1 vssd1 vccd1 vccd1 _09610_/B sky130_fd_sc_hd__xnor2_1
X_10881_ _12648_/A _10879_/Y _10880_/Y _09529_/B vssd1 vssd1 vccd1 vccd1 _10897_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__10673__A3 _10787_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12620_ _12620_/A _12671_/A vssd1 vssd1 vccd1 vccd1 _12621_/C sky130_fd_sc_hd__and2_1
XANTENNA__08318__A _08746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07826__A1 _09216_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12551_ _12551_/A _12551_/B vssd1 vssd1 vccd1 vccd1 _12552_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_65_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07826__B2 _08868_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11502_ _11503_/A _11503_/B vssd1 vssd1 vccd1 vccd1 _11646_/B sky130_fd_sc_hd__and2b_1
X_12482_ _12414_/A _12414_/B _12412_/A vssd1 vssd1 vccd1 vccd1 _12494_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__12782__B _12782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11433_ _11302_/B _11302_/C _11302_/A vssd1 vssd1 vccd1 vccd1 _11436_/A sky130_fd_sc_hd__a21boi_2
XFILLER_0_124_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07876__B _11823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10583__A _10981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11364_ _09836_/X _11363_/X _11576_/A vssd1 vssd1 vccd1 vccd1 _11364_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_104_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13103_ _13084_/B _13102_/X _13129_/B _07634_/C vssd1 vssd1 vccd1 vccd1 _13105_/B
+ sky130_fd_sc_hd__a2bb2o_2
X_10315_ _09668_/X _09675_/X _10600_/S vssd1 vssd1 vccd1 vccd1 _10315_/X sky130_fd_sc_hd__mux2_1
X_11295_ _11603_/A _11295_/B vssd1 vssd1 vccd1 vccd1 _11299_/A sky130_fd_sc_hd__xnor2_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13034_ _13039_/B _13034_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[10] sky130_fd_sc_hd__and2_4
X_10246_ _11281_/A _10246_/B vssd1 vssd1 vccd1 vccd1 _10250_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_119_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_4_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10177_ _10600_/S _09473_/X _10176_/X vssd1 vssd1 vccd1 vccd1 _10178_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_100_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07762__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08306__A2 wire122/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09503__A1 _12648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07514__B1 _07535_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12818_ reg1_val[3] curr_PC[3] _12825_/S vssd1 vssd1 vccd1 vccd1 _12820_/B sky130_fd_sc_hd__mux2_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _12749_/A _12749_/B vssd1 vssd1 vccd1 vccd1 _12749_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_57_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08490__A1 _09216_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08490__B2 _08868_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13366__A2 _13542_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10493__A _11913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09960_ _09960_/A _09960_/B vssd1 vssd1 vccd1 vccd1 _09961_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09493__S _09493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08911_ _08911_/A _08911_/B vssd1 vssd1 vccd1 vccd1 _08916_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_0_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09891_ _12092_/A _09891_/B vssd1 vssd1 vccd1 vccd1 _09893_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _08814_/B _08814_/C _08814_/A vssd1 vssd1 vccd1 vccd1 _08842_/X sky130_fd_sc_hd__a21o_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12213__A _12695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10352__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ _10236_/A _08773_/B vssd1 vssd1 vccd1 vccd1 _08804_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13028__B _13029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout184_A _13450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07724_ _09575_/A _07724_/B vssd1 vssd1 vccd1 vccd1 _07731_/A sky130_fd_sc_hd__xnor2_1
X_07655_ _07655_/A _07655_/B vssd1 vssd1 vccd1 vccd1 _07658_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06865__B _13005_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07586_ _07696_/A _07585_/Y _07584_/A vssd1 vssd1 vccd1 vccd1 _07588_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_94_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09325_ _09325_/A _09325_/B vssd1 vssd1 vccd1 vccd1 _09427_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11604__A2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12883__A _13042_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07977__A _10078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09256_ _11958_/A _09254_/X _06790_/X vssd1 vssd1 vccd1 vccd1 fanout5/A sky130_fd_sc_hd__a21o_2
XANTENNA__08481__A1 _08873_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08481__B2 _08891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08207_ _08873_/A2 fanout82/X fanout76/X _08891_/B vssd1 vssd1 vccd1 vccd1 _08208_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_106_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09187_ _07930_/A _07930_/B _07944_/B _07945_/B _07945_/A vssd1 vssd1 vccd1 vccd1
+ _09197_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_90_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08138_ _08806_/A2 _07477_/X _13172_/A1 _08806_/B1 vssd1 vssd1 vccd1 vccd1 _08139_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08069_ _08156_/A _08156_/B _08058_/Y vssd1 vssd1 vccd1 vccd1 _08090_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_3_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12317__B1 _11688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10100_ _10100_/A _10100_/B vssd1 vssd1 vccd1 vccd1 _10102_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout97_A _11512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11080_ _10910_/A _10910_/B _10908_/Y vssd1 vssd1 vccd1 vccd1 _11082_/B sky130_fd_sc_hd__o21a_1
X_10031_ hold285/A hold262/A hold245/A vssd1 vssd1 vccd1 vccd1 _10031_/X sky130_fd_sc_hd__or3_1
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11982_ _07137_/Y _11968_/X _11981_/X _11962_/X vssd1 vssd1 vccd1 vccd1 _11982_/Y
+ sky130_fd_sc_hd__a211oi_2
X_13721_ _13725_/CLK _13721_/D vssd1 vssd1 vccd1 vccd1 hold292/A sky130_fd_sc_hd__dfxtp_1
X_10933_ _10778_/A _10778_/B _10777_/A vssd1 vssd1 vccd1 vccd1 _10939_/A sky130_fd_sc_hd__o21ai_2
X_10864_ _11562_/A _10864_/B _10864_/C vssd1 vssd1 vccd1 vccd1 _10864_/X sky130_fd_sc_hd__or3_1
X_13652_ _13659_/CLK hold211/X vssd1 vssd1 vccd1 vccd1 hold209/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10297__B _10631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12603_ _12593_/Y _12594_/X _12598_/X _12602_/X vssd1 vssd1 vccd1 vccd1 _12603_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11056__B1 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12399__A3 _12235_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10795_ _10666_/A _10666_/B _10665_/A vssd1 vssd1 vccd1 vccd1 _10796_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_109_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13583_ _13605_/A _13583_/B vssd1 vssd1 vccd1 vccd1 _13734_/D sky130_fd_sc_hd__and2_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12534_ _12534_/A _12534_/B _12754_/C vssd1 vssd1 vccd1 vccd1 _12534_/X sky130_fd_sc_hd__and3_1
XFILLER_0_109_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13348__A2 _13506_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12465_ _12786_/B1 _12527_/B hold278/A vssd1 vssd1 vccd1 vccd1 _12465_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12556__B1 _12557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11416_ _11417_/A _11417_/B vssd1 vssd1 vccd1 vccd1 _11538_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12396_ _07221_/A _12799_/A2 _12657_/B1 reg1_val[24] vssd1 vssd1 vccd1 vccd1 _12396_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_22_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11347_ _11554_/A _11347_/B vssd1 vssd1 vccd1 vccd1 _11600_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__07983__B1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09607__A _10522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11278_ _11279_/A _11279_/B vssd1 vssd1 vccd1 vccd1 _11388_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_39_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08527__A2 _09173_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13017_ _13017_/A _13017_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[7] sky130_fd_sc_hd__xor2_4
XANTENNA__13129__A _13129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10229_ _10229_/A _10229_/B vssd1 vssd1 vccd1 vccd1 _10233_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07735__B1 _11638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07440_ _07634_/B _07435_/B reg1_val[18] vssd1 vssd1 vccd1 vccd1 _11884_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07371_ reg1_val[27] _07865_/B vssd1 vssd1 vccd1 vccd1 _07641_/A sky130_fd_sc_hd__or2_2
XANTENNA__13587__A2 fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09110_ _09110_/A _09110_/B vssd1 vssd1 vccd1 vccd1 _09111_/B sky130_fd_sc_hd__and2_1
XANTENNA__09488__S _10007_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09041_ _09044_/A _09041_/B vssd1 vssd1 vccd1 vccd1 _09048_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_60_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12547__B1 _12971_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap153 _07399_/Y vssd1 vssd1 vccd1 vccd1 _09604_/A sky130_fd_sc_hd__buf_6
XFILLER_0_123_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09943_ _09944_/A _09944_/B vssd1 vssd1 vccd1 vccd1 _09945_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13511__A2 _13555_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ _12648_/A _09860_/B _09868_/Y _07016_/Y _09873_/X vssd1 vssd1 vccd1 vccd1
+ _09874_/X sky130_fd_sc_hd__o221a_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08825_ _08828_/A _08828_/B vssd1 vssd1 vccd1 vccd1 _08825_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_99_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08756_ _08756_/A _08756_/B vssd1 vssd1 vccd1 vccd1 _08762_/B sky130_fd_sc_hd__xnor2_1
X_07707_ _07707_/A _07707_/B _07718_/A vssd1 vssd1 vccd1 vccd1 _07708_/B sky130_fd_sc_hd__nand3_1
X_08687_ _08687_/A _08687_/B vssd1 vssd1 vccd1 vccd1 _08728_/B sky130_fd_sc_hd__xor2_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07638_ _07641_/C _07641_/D vssd1 vssd1 vccd1 vccd1 _07639_/B sky130_fd_sc_hd__and2_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07569_ _11508_/A _07569_/B vssd1 vssd1 vccd1 vccd1 _07583_/A sky130_fd_sc_hd__xnor2_1
X_09308_ _09308_/A _09308_/B vssd1 vssd1 vccd1 vccd1 _09310_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13502__A _13543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10580_ _10294_/X _10430_/X _10431_/X vssd1 vssd1 vccd1 vccd1 _10580_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_91_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout12_A fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12250__A2 _07597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09239_ _09239_/A _09239_/B vssd1 vssd1 vccd1 vccd1 _09264_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_23_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12250_ fanout35/X _07597_/X _07891_/X _07699_/B vssd1 vssd1 vccd1 vccd1 _12251_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12002__A2 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11201_ _11202_/A _11202_/B vssd1 vssd1 vccd1 vccd1 _11203_/A sky130_fd_sc_hd__nand2_1
X_12181_ _12258_/A _12181_/B vssd1 vssd1 vccd1 vccd1 _12182_/B sky130_fd_sc_hd__nor2_1
X_11132_ _11127_/X _11129_/Y _11131_/X _12648_/A vssd1 vssd1 vccd1 vccd1 _11132_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11063_ _11064_/A _11064_/B vssd1 vssd1 vccd1 vccd1 _11065_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11513__A1 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10014_ reg1_val[3] curr_PC[3] vssd1 vssd1 vccd1 vccd1 _10016_/C sky130_fd_sc_hd__nand2_1
XANTENNA__11513__B2 _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11965_ _11965_/A _11965_/B vssd1 vssd1 vccd1 vccd1 _11967_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_86_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13704_ _13705_/CLK hold125/X vssd1 vssd1 vccd1 vccd1 _13704_/Q sky130_fd_sc_hd__dfxtp_1
X_10916_ _10917_/A _10917_/B vssd1 vssd1 vccd1 vccd1 _10916_/X sky130_fd_sc_hd__and2_1
XANTENNA__07496__A2 _07491_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09890__B1 _07472_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11896_ _12372_/A _12372_/B _11896_/C _12163_/C vssd1 vssd1 vccd1 vccd1 _11988_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_0_67_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13635_ _13731_/CLK _13635_/D vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10847_ _10847_/A _10847_/B vssd1 vssd1 vccd1 vccd1 _10849_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08445__A1 _08866_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08445__B2 _09216_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13566_ hold278/A _13565_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13566_/X sky130_fd_sc_hd__mux2_1
X_10778_ _10778_/A _10778_/B vssd1 vssd1 vccd1 vccd1 _10780_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12517_ _12516_/A _12516_/B _12516_/Y _09507_/X vssd1 vssd1 vccd1 vccd1 _12517_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_124_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13497_ _13543_/A hold281/X vssd1 vssd1 vccd1 vccd1 _13715_/D sky130_fd_sc_hd__and2_1
XFILLER_0_54_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12448_ _12480_/B _12447_/X _10730_/B vssd1 vssd1 vccd1 vccd1 _12448_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__13558__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08748__A2 _07492_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07405__C1 _07398_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12379_ _12379_/A _12379_/B vssd1 vssd1 vccd1 vccd1 _12379_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_50_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11586__B _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06940_ _07535_/A _07476_/A vssd1 vssd1 vccd1 vccd1 _06943_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11504__A1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11504__B2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09173__A2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06871_ _06886_/A _13010_/B vssd1 vssd1 vccd1 vccd1 _06871_/Y sky130_fd_sc_hd__nor2_1
X_08610_ _08610_/A _08610_/B vssd1 vssd1 vccd1 vccd1 _08658_/B sky130_fd_sc_hd__xnor2_1
X_09590_ _10814_/A1 fanout83/X fanout79/X fanout42/X vssd1 vssd1 vccd1 vccd1 _09591_/B
+ sky130_fd_sc_hd__o22a_1
X_08541_ _08544_/A _08544_/B vssd1 vssd1 vccd1 vccd1 _08545_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08472_ _08472_/A _08472_/B vssd1 vssd1 vccd1 vccd1 _08475_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_106_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07423_ _09910_/A1 fanout14/X _09955_/A _07833_/B vssd1 vssd1 vccd1 vccd1 _07424_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10946__A _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07354_ _07360_/A _07360_/B vssd1 vssd1 vccd1 vccd1 _12093_/A sky130_fd_sc_hd__nand2_8
XFILLER_0_73_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07320__A _13015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13041__B _13042_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07285_ _10366_/A _07285_/B vssd1 vssd1 vccd1 vccd1 _07285_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_32_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09024_ _09023_/A _09023_/C _09023_/B vssd1 vssd1 vccd1 vccd1 _09025_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09936__A1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold220 hold220/A vssd1 vssd1 vccd1 vccd1 hold220/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09936__B2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold231 hold231/A vssd1 vssd1 vccd1 vccd1 hold231/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 hold242/A vssd1 vssd1 vccd1 vccd1 hold242/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 hold253/A vssd1 vssd1 vccd1 vccd1 hold253/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold264 hold264/A vssd1 vssd1 vccd1 vccd1 hold264/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 hold275/A vssd1 vssd1 vccd1 vccd1 hold275/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 hold286/A vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 hold297/A vssd1 vssd1 vccd1 vccd1 hold297/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09926_ fanout45/X fanout68/X fanout66/X fanout49/X vssd1 vssd1 vccd1 vccd1 _09927_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13496__B2 _13542_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09857_ _09855_/Y _09857_/B vssd1 vssd1 vccd1 vccd1 _09858_/B sky130_fd_sc_hd__nand2b_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07175__A1 _10239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08372__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08808_ _08873_/A2 _13149_/A _08923_/B1 _08891_/B vssd1 vssd1 vccd1 vccd1 _08809_/B
+ sky130_fd_sc_hd__o22a_1
X_09788_ _09788_/A _09788_/B vssd1 vssd1 vccd1 vccd1 _09789_/B sky130_fd_sc_hd__xnor2_1
X_08739_ _08739_/A _08739_/B vssd1 vssd1 vccd1 vccd1 _08766_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08124__B1 _09949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08675__A1 _09674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _11751_/A _11751_/B vssd1 vssd1 vccd1 vccd1 _11849_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__12471__A2 _12799_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08675__B2 _08873_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10482__A1 _12825_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10701_ _10702_/A _10798_/B _10701_/C vssd1 vssd1 vccd1 vccd1 _10701_/X sky130_fd_sc_hd__and3_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11681_ _11679_/Y _11681_/B vssd1 vssd1 vccd1 vccd1 _11682_/B sky130_fd_sc_hd__and2b_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13420_ hold151/A _13142_/A _13420_/B1 hold113/X _13430_/C1 vssd1 vssd1 vccd1 vccd1
+ hold114/A sky130_fd_sc_hd__o221a_1
X_10632_ _09325_/A _09325_/B _10150_/X _10631_/X vssd1 vssd1 vccd1 vccd1 _10632_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_102_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07230__A _07230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10563_ _10564_/A _10564_/B vssd1 vssd1 vccd1 vccd1 _10563_/Y sky130_fd_sc_hd__nor2_1
X_13351_ _13359_/A hold232/X vssd1 vssd1 vccd1 vccd1 _13657_/D sky130_fd_sc_hd__and2_1
XFILLER_0_36_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10785__A2 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12302_ _12515_/S _12301_/X _12300_/X vssd1 vssd1 vccd1 vccd1 _12303_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_23_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10494_ _10495_/A _10495_/B vssd1 vssd1 vccd1 vccd1 _10496_/A sky130_fd_sc_hd__nand2_1
X_13282_ hold245/X hold11/X vssd1 vssd1 vccd1 vccd1 _13451_/A sky130_fd_sc_hd__xor2_1
X_12233_ hold255/A _12314_/A _12313_/B _12796_/A1 vssd1 vssd1 vccd1 vccd1 _12234_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_121_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12164_ _12164_/A _12164_/B _12164_/C _12164_/D vssd1 vssd1 vccd1 vccd1 _12373_/A
+ sky130_fd_sc_hd__nor4_2
XANTENNA__07402__A2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11115_ _11115_/A _11115_/B vssd1 vssd1 vccd1 vccd1 _11115_/X sky130_fd_sc_hd__or2_1
X_12095_ _12096_/A _12096_/B vssd1 vssd1 vccd1 vccd1 _12187_/B sky130_fd_sc_hd__nand2_1
X_11046_ _11823_/A _11046_/B vssd1 vssd1 vccd1 vccd1 _11048_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07166__A1 _07535_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09604__B _10518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap112_A _07492_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12997_ _12997_/A _12997_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[3] sky130_fd_sc_hd__xnor2_4
XFILLER_0_98_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07124__B _07129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11948_ _11948_/A _12035_/A vssd1 vssd1 vccd1 vccd1 _12125_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11670__B1 _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11879_ _12311_/B1 _11972_/B hold203/A vssd1 vssd1 vccd1 vccd1 _11879_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__06963__B _10889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13142__A _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13618_ _13725_/CLK _13618_/D vssd1 vssd1 vccd1 vccd1 hold111/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13549_ hold266/A _13548_/Y hold234/X vssd1 vssd1 vccd1 vccd1 _13549_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07070_ _06848_/D _07069_/X _07062_/Y vssd1 vssd1 vccd1 vccd1 _07070_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_125_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07972_ _09575_/A _07972_/B vssd1 vssd1 vccd1 vccd1 _07978_/A sky130_fd_sc_hd__xnor2_2
X_09711_ _09507_/X _09702_/Y _09703_/X _09710_/X vssd1 vssd1 vccd1 vccd1 _09711_/X
+ sky130_fd_sc_hd__o31a_1
X_06923_ _06923_/A _07527_/A vssd1 vssd1 vccd1 vccd1 _06923_/X sky130_fd_sc_hd__or2_1
X_09642_ _09642_/A _09642_/B vssd1 vssd1 vccd1 vccd1 _09644_/A sky130_fd_sc_hd__xnor2_2
X_06854_ _07334_/B _07230_/A vssd1 vssd1 vccd1 vccd1 _06856_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_97_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13036__B _13036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09573_ _10095_/A _09573_/B vssd1 vssd1 vccd1 vccd1 _09577_/A sky130_fd_sc_hd__xnor2_1
X_06785_ instruction[1] instruction[2] instruction[25] pred_val vssd1 vssd1 vccd1
+ vccd1 _06785_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_0_26_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout264_A _13082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ _09674_/S fanout84/X _08580_/B _08873_/B2 vssd1 vssd1 vccd1 vccd1 _08525_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10464__A1 _12314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08455_ _08455_/A _08455_/B vssd1 vssd1 vccd1 vccd1 _08456_/B sky130_fd_sc_hd__or2_1
X_07406_ _10456_/S _07407_/B vssd1 vssd1 vccd1 vccd1 _07406_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_9_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08386_ _08389_/A _08389_/B vssd1 vssd1 vccd1 vccd1 _08391_/A sky130_fd_sc_hd__nor2_1
XANTENNA__09606__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07337_ _07377_/A _07337_/B vssd1 vssd1 vccd1 vccd1 _07337_/Y sky130_fd_sc_hd__nand2_1
X_07268_ _10095_/A vssd1 vssd1 vccd1 vccd1 _10542_/A sky130_fd_sc_hd__inv_6
XFILLER_0_60_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09007_ _08951_/A _08953_/Y _09005_/A vssd1 vssd1 vccd1 vccd1 _09008_/B sky130_fd_sc_hd__o21ba_1
X_07199_ _07200_/A _07200_/B vssd1 vssd1 vccd1 vccd1 _08933_/B sky130_fd_sc_hd__and2_4
XFILLER_0_13_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08593__B1 _08778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09909_ _09909_/A _09909_/B vssd1 vssd1 vccd1 vccd1 _09912_/A sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_4_9_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12920_ _12956_/A _12920_/B vssd1 vssd1 vccd1 vccd1 _12921_/B sky130_fd_sc_hd__or2_1
X_12851_ _12851_/A _12851_/B _12851_/C vssd1 vssd1 vccd1 vccd1 _12852_/B sky130_fd_sc_hd__nand3_1
X_11802_ wire101/X _11802_/B vssd1 vssd1 vccd1 vccd1 _11804_/B sky130_fd_sc_hd__nand2_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _13129_/A _12782_/B _12782_/C vssd1 vssd1 vccd1 vccd1 _12783_/B sky130_fd_sc_hd__and3_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _11733_/A _11733_/B vssd1 vssd1 vccd1 vccd1 _11735_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06783__B _12981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11664_ _11451_/Y _11857_/A _11662_/X vssd1 vssd1 vccd1 vccd1 _11664_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10207__A1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13403_ _07575_/B _13419_/A2 hold20/X vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__o21a_1
XANTENNA__10207__B2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10615_ _10605_/Y _10606_/X _10614_/X vssd1 vssd1 vccd1 vccd1 _10615_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11404__B1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11595_ _11955_/A _11560_/X _11561_/Y _11564_/X _11594_/X vssd1 vssd1 vccd1 vccd1
+ _11595_/X sky130_fd_sc_hd__o311a_1
XFILLER_0_107_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07895__A _09659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13334_ hold180/X _13506_/B2 _13506_/A2 hold163/X vssd1 vssd1 vccd1 vccd1 hold181/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07623__A2 _08873_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10546_ _10546_/A _10546_/B _10546_/C vssd1 vssd1 vccd1 vccd1 _10686_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_122_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13265_ hold68/X hold276/X vssd1 vssd1 vccd1 vccd1 _13265_/X sky130_fd_sc_hd__and2b_1
X_10477_ _12047_/C1 _10449_/X _10476_/X vssd1 vssd1 vccd1 vccd1 _10477_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_122_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12216_ _12136_/A _12134_/X _07054_/Y vssd1 vssd1 vccd1 vccd1 _12216_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_121_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13196_ _12413_/A _13196_/A2 hold40/X _13591_/A vssd1 vssd1 vccd1 vccd1 hold41/A
+ sky130_fd_sc_hd__o211a_1
X_12147_ hold266/A _12058_/A _12231_/B _12748_/B1 vssd1 vssd1 vccd1 vccd1 _12147_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12078_ _12666_/A _12078_/B vssd1 vssd1 vccd1 vccd1 _12082_/A sky130_fd_sc_hd__xnor2_1
X_11029_ _11029_/A _11029_/B _11029_/C vssd1 vssd1 vccd1 vccd1 _11030_/B sky130_fd_sc_hd__or3_1
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06898__B1 _06980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13571__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08240_ _08240_/A _08240_/B vssd1 vssd1 vccd1 vccd1 _08242_/B sky130_fd_sc_hd__xor2_2
XANTENNA__06906__A2_N _06980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_15 instruction[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 reg1_val[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_37 reg1_val[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08171_ _08130_/A _08129_/B _08129_/C vssd1 vssd1 vccd1 vccd1 _08174_/B sky130_fd_sc_hd__a21o_1
XANTENNA_48 reg2_val[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_59 reg2_val[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10749__A2 _12793_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09496__S _09496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07122_ instruction[13] _07122_/B vssd1 vssd1 vccd1 vccd1 dest_pred[2] sky130_fd_sc_hd__and2_4
XFILLER_0_6_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07053_ reg1_val[22] _07212_/B vssd1 vssd1 vccd1 vccd1 _07053_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_70_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09525__A _13744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07955_ _07956_/B _07956_/A vssd1 vssd1 vccd1 vccd1 _07955_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__06868__B _07201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13320__B1 _13450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06906_ reg2_val[16] _06980_/B _06906_/B1 _06905_/Y vssd1 vssd1 vccd1 vccd1 _07297_/A
+ sky130_fd_sc_hd__o2bb2a_2
X_07886_ _09951_/A _07886_/B vssd1 vssd1 vccd1 vccd1 _07900_/A sky130_fd_sc_hd__xnor2_2
X_09625_ _09625_/A _09625_/B vssd1 vssd1 vccd1 vccd1 _09626_/B sky130_fd_sc_hd__or2_1
X_06837_ _06840_/A vssd1 vssd1 vccd1 vccd1 _06837_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09556_ _09557_/B vssd1 vssd1 vccd1 vccd1 _09556_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06768_ instruction[20] instruction[13] _07135_/S vssd1 vssd1 vccd1 vccd1 reg1_idx[2]
+ sky130_fd_sc_hd__mux2_8
X_08507_ _08507_/A _08507_/B vssd1 vssd1 vccd1 vccd1 _08574_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07699__B _07699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07302__A1 _13015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09487_ _09485_/X _09486_/X _09688_/S vssd1 vssd1 vccd1 vccd1 _09487_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_92_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08438_ _08438_/A _08505_/A vssd1 vssd1 vccd1 vccd1 _08451_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_19_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08369_ _08370_/A _08370_/B vssd1 vssd1 vccd1 vccd1 _08369_/X sky130_fd_sc_hd__and2_1
XANTENNA__12825__S _12825_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10400_ fanout38/X _07543_/X fanout70/X fanout36/X vssd1 vssd1 vccd1 vccd1 _10401_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_61_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11380_ _11356_/Y _11357_/X _11379_/X vssd1 vssd1 vccd1 vccd1 _11380_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_0_21_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10331_ _10170_/A _10167_/Y _10169_/B vssd1 vssd1 vccd1 vccd1 _10335_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_14_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13050_ _13051_/A _13051_/B _13051_/C vssd1 vssd1 vccd1 vccd1 _13057_/B sky130_fd_sc_hd__a21o_1
X_10262_ _10814_/A1 fanout29/X _07453_/Y fanout42/X vssd1 vssd1 vccd1 vccd1 _10263_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07369__A1 _08866_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07369__B2 _08118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12001_ _12001_/A _12001_/B vssd1 vssd1 vccd1 vccd1 _12012_/A sky130_fd_sc_hd__nand2_1
X_10193_ _10458_/S _10192_/X _09537_/B vssd1 vssd1 vccd1 vccd1 _10193_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__10912__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06778__B _07110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12665__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12903_ _13059_/B _12904_/B vssd1 vssd1 vccd1 vccd1 _12912_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07541__A1 _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12834_ _13005_/B _12834_/B vssd1 vssd1 vccd1 vccd1 _12835_/B sky130_fd_sc_hd__or2_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11625__B1 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _12765_/A _12765_/B vssd1 vssd1 vccd1 vccd1 _12765_/Y sky130_fd_sc_hd__nor2_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _12092_/A _11716_/B vssd1 vssd1 vccd1 vccd1 _11717_/A sky130_fd_sc_hd__xnor2_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _09321_/A _12695_/X _11866_/A vssd1 vssd1 vccd1 vccd1 _12696_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13378__B1 _13584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11647_ _11647_/A _11647_/B vssd1 vssd1 vccd1 vccd1 _11648_/B sky130_fd_sc_hd__and2_1
XFILLER_0_64_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11578_ _11574_/Y _11577_/Y _12225_/A vssd1 vssd1 vccd1 vccd1 _11578_/X sky130_fd_sc_hd__mux2_1
X_13317_ _13589_/B _13316_/Y _13315_/X vssd1 vssd1 vccd1 vccd1 hold234/A sky130_fd_sc_hd__a21o_1
XFILLER_0_12_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10529_ _11823_/A _10529_/B vssd1 vssd1 vccd1 vccd1 _10531_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13248_ hold126/X hold296/A vssd1 vssd1 vccd1 vccd1 _13248_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_122_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13566__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10364__B1 _10536_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13179_ hold55/X _13191_/B vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__or2_1
X_07740_ _10542_/A _07740_/B vssd1 vssd1 vccd1 vccd1 _07819_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10116__B1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07671_ _07671_/A _07671_/B vssd1 vssd1 vccd1 vccd1 _07672_/B sky130_fd_sc_hd__or2_1
XANTENNA__07532__A1 _07572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09410_ _09410_/A _09410_/B vssd1 vssd1 vccd1 vccd1 _09423_/A sky130_fd_sc_hd__xor2_4
XANTENNA__12408__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09341_ _09342_/B _09342_/A vssd1 vssd1 vccd1 vccd1 _09341_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_87_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07296__B1 _07521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09272_ _09955_/A _07643_/B fanout13/X _09910_/A1 vssd1 vssd1 vccd1 vccd1 _09273_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08223_ _08223_/A _08223_/B vssd1 vssd1 vccd1 vccd1 _08226_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_7_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08154_ _08162_/A _08162_/B vssd1 vssd1 vccd1 vccd1 _08234_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12041__B1 _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11395__A2 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08796__B1 _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07105_ instruction[1] _07123_/A vssd1 vssd1 vccd1 vccd1 _07108_/D sky130_fd_sc_hd__and2_4
X_08085_ _13151_/A fanout28/X _08395_/B _08866_/A2 vssd1 vssd1 vccd1 vccd1 _08086_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07036_ _10447_/B _10447_/C _10449_/A vssd1 vssd1 vccd1 vccd1 _10588_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_2_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08012__A2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06879__A _06886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07220__B1 _07521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__A2 _10787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ _09068_/A _09077_/B _08572_/Y _09057_/B vssd1 vssd1 vccd1 vccd1 _08988_/C
+ sky130_fd_sc_hd__or4bb_1
X_07938_ _09119_/A _07938_/B vssd1 vssd1 vccd1 vccd1 _07940_/C sky130_fd_sc_hd__nand2_1
X_07869_ _07869_/A _11731_/A vssd1 vssd1 vccd1 vccd1 _07870_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09608_ _09609_/A _09609_/B vssd1 vssd1 vccd1 vccd1 _09608_/X sky130_fd_sc_hd__and2b_1
X_10880_ _12648_/A _10880_/B vssd1 vssd1 vccd1 vccd1 _10880_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_85_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout42_A _07282_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09539_ instruction[5] _07075_/Y _09509_/A _09503_/X _09538_/X vssd1 vssd1 vccd1
+ vccd1 _09539_/X sky130_fd_sc_hd__o311a_1
XFILLER_0_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12550_ _12551_/A _12551_/B vssd1 vssd1 vccd1 vccd1 _12552_/A sky130_fd_sc_hd__and2_1
XANTENNA__07826__A2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11501_ _11731_/A _11501_/B vssd1 vssd1 vccd1 vccd1 _11503_/B sky130_fd_sc_hd__xnor2_2
X_12481_ _12733_/A _12635_/A _12735_/A1 vssd1 vssd1 vccd1 vccd1 _12513_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_46_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11432_ _11319_/B _11319_/C _11319_/A vssd1 vssd1 vccd1 vccd1 _11443_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_61_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11363_ _10316_/X _10318_/X _11472_/S vssd1 vssd1 vccd1 vccd1 _11363_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13102_ _13102_/A _13102_/B _13102_/C _13102_/D vssd1 vssd1 vccd1 vccd1 _13102_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_0_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10314_ _11576_/A _10313_/A _09535_/Y vssd1 vssd1 vccd1 vccd1 _12525_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__11269__A2_N fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11294_ fanout54/X fanout38/X _07368_/Y _12268_/A vssd1 vssd1 vccd1 vccd1 _11295_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08539__B1 _09885_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13033_ _13033_/A _13033_/B _13033_/C vssd1 vssd1 vccd1 vccd1 _13034_/B sky130_fd_sc_hd__nand3_1
X_10245_ fanout53/X fanout83/X fanout79/X fanout47/X vssd1 vssd1 vccd1 vccd1 _10246_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06789__A _06936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10176_ _10176_/A _10176_/B vssd1 vssd1 vccd1 vccd1 _10176_/X sky130_fd_sc_hd__or2_1
XANTENNA__07762__A1 _08907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07762__B2 _08328_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10104__A _10104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout190 _09524_/Y vssd1 vssd1 vccd1 vccd1 _12795_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12817_ _12823_/B _12817_/B vssd1 vssd1 vccd1 vccd1 new_PC[2] sky130_fd_sc_hd__and2_4
XFILLER_0_84_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07278__B1 _07594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ hold233/A _12786_/B1 _12746_/X _12748_/B1 vssd1 vssd1 vccd1 vccd1 _12749_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08490__A2 _10538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10774__A _11913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12679_ _12677_/A _12677_/B _12677_/C vssd1 vssd1 vccd1 vccd1 _12680_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07450__B1 _07476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08910_ _08910_/A _08910_/B _08910_/C vssd1 vssd1 vccd1 vccd1 _08920_/A sky130_fd_sc_hd__or3_2
XFILLER_0_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ fanout14/X _07455_/Y _07472_/Y _07833_/B vssd1 vssd1 vccd1 vccd1 _09891_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07202__B1 _07521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08841_ _08814_/B _08814_/C _08814_/A vssd1 vssd1 vccd1 vccd1 _08976_/B sky130_fd_sc_hd__a21oi_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ _08891_/B _08866_/A2 _08923_/B1 _08873_/A2 vssd1 vssd1 vccd1 vccd1 _08773_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07723_ fanout76/X fanout68/X fanout66/X fanout74/X vssd1 vssd1 vccd1 vccd1 _07724_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08702__B1 _08778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout177_A _07476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13325__A _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07654_ _07654_/A _07654_/B vssd1 vssd1 vccd1 vccd1 _07655_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_95_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07585_ _07696_/B vssd1 vssd1 vccd1 vccd1 _07585_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_48_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09324_ _09825_/A _09204_/X _09986_/A _09828_/B _09828_/A vssd1 vssd1 vccd1 vccd1
+ _09325_/B sky130_fd_sc_hd__o32a_1
XFILLER_0_75_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09255_ _11958_/A _09254_/X _06790_/X vssd1 vssd1 vccd1 vccd1 fanout7/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_63_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08481__A2 _10049_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06881__B _07281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08206_ _08205_/B _08205_/C _08205_/A vssd1 vssd1 vccd1 vccd1 _08217_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_62_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07469__S _11709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09186_ _09186_/A _09186_/B vssd1 vssd1 vccd1 vccd1 _09198_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_31_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08769__B1 _08868_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08137_ _10236_/A _08137_/B vssd1 vssd1 vccd1 vccd1 _08140_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09430__A1 _12695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08068_ _08068_/A _08068_/B vssd1 vssd1 vccd1 vccd1 _08156_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_31_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12317__A1 _07230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07019_ instruction[41] _06781_/X _06784_/X _06895_/Y _07110_/A vssd1 vssd1 vccd1
+ vccd1 _07025_/C sky130_fd_sc_hd__a2111o_4
XFILLER_0_101_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10328__B1 _12657_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10030_ _07010_/B _12793_/A2 _11586_/B vssd1 vssd1 vccd1 vccd1 _10030_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__08941__B1 _07420_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11981_ _09521_/Y _11970_/Y _11971_/X _11980_/X vssd1 vssd1 vccd1 vccd1 _11981_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13720_ _13725_/CLK _13720_/D vssd1 vssd1 vccd1 vccd1 hold296/A sky130_fd_sc_hd__dfxtp_2
X_10932_ _10932_/A _10932_/B vssd1 vssd1 vccd1 vccd1 _10941_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08329__A _09950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13651_ _13659_/CLK hold242/X vssd1 vssd1 vccd1 vccd1 _13651_/Q sky130_fd_sc_hd__dfxtp_1
X_10863_ _10863_/A _10863_/B vssd1 vssd1 vccd1 vccd1 _10863_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_39_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12602_ _09839_/A _10180_/Y _10193_/Y _09860_/A _12601_/X vssd1 vssd1 vccd1 vccd1
+ _12602_/X sky130_fd_sc_hd__o221a_1
XANTENNA__11056__A1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11056__B2 _12557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13582_ hold268/X _13584_/B _13581_/X _13599_/D vssd1 vssd1 vccd1 vccd1 _13583_/B
+ sky130_fd_sc_hd__a22o_1
X_10794_ _10794_/A _10794_/B vssd1 vssd1 vccd1 vccd1 _10796_/A sky130_fd_sc_hd__xnor2_2
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12533_ hold166/A _12374_/A _12592_/B _12533_/B1 vssd1 vssd1 vccd1 vccd1 _12533_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_81_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12005__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12464_ hold269/A _12464_/B vssd1 vssd1 vccd1 vccd1 _12527_/B sky130_fd_sc_hd__or2_1
XANTENNA__12556__A1 _12557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11415_ _11415_/A _11415_/B vssd1 vssd1 vccd1 vccd1 _11417_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12395_ hold216/A _12374_/A _12467_/B _12795_/A1 vssd1 vssd1 vccd1 vccd1 _12395_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11346_ _10860_/B _11343_/Y _11345_/X vssd1 vssd1 vccd1 vccd1 _11347_/B sky130_fd_sc_hd__o21bai_4
XFILLER_0_22_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07983__A1 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07983__B2 _08328_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11277_ _12417_/A _11277_/B vssd1 vssd1 vccd1 vccd1 _11279_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12314__A _12314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13016_ _13014_/Y _13016_/B vssd1 vssd1 vccd1 vccd1 _13017_/B sky130_fd_sc_hd__nand2b_2
X_10228_ _10229_/A _10229_/B vssd1 vssd1 vccd1 vccd1 _10392_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__13129__B _13129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07735__A1 _07300_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07196__C1 _07201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07735__B2 _08806_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07127__B _07129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10159_ _11562_/A _10160_/B _10160_/C vssd1 vssd1 vccd1 vccd1 _10159_/Y sky130_fd_sc_hd__o21ai_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09623__A _10263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13145__A _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07370_ _10119_/A _07370_/B vssd1 vssd1 vccd1 vccd1 _07425_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06982__A _07556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12795__A1 _12795_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09040_ _09039_/A _09039_/B _11460_/B vssd1 vssd1 vccd1 vccd1 _11562_/B sky130_fd_sc_hd__o21ba_2
XFILLER_0_44_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmax_cap121 _07455_/Y vssd1 vssd1 vccd1 vccd1 _13166_/A1 sky130_fd_sc_hd__buf_4
XFILLER_0_111_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07423__B1 _09955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmax_cap176 _07185_/C vssd1 vssd1 vccd1 vccd1 _07187_/B sky130_fd_sc_hd__buf_1
X_09942_ _11072_/A _09942_/B vssd1 vssd1 vccd1 vccd1 _09944_/B sky130_fd_sc_hd__xnor2_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ _09496_/S _11793_/B _11587_/A2 _07015_/Y _09872_/X vssd1 vssd1 vccd1 vccd1
+ _09873_/X sky130_fd_sc_hd__o221a_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout294_A _12578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08923__B1 _08923_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08824_ _09659_/B _08824_/B vssd1 vssd1 vccd1 vccd1 _08828_/B sky130_fd_sc_hd__xnor2_2
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09533__A _10457_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08755_ _08755_/A _08755_/B _08756_/B vssd1 vssd1 vccd1 vccd1 _08755_/X sky130_fd_sc_hd__and3_1
X_07706_ _07707_/B _07718_/A _07707_/A vssd1 vssd1 vccd1 vccd1 _07708_/A sky130_fd_sc_hd__a21o_1
X_08686_ _08686_/A _08686_/B vssd1 vssd1 vccd1 vccd1 _08728_/A sky130_fd_sc_hd__xor2_1
XANTENNA__12483__B1 _09145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07637_ _12647_/A _07637_/B vssd1 vssd1 vccd1 vccd1 _07641_/D sky130_fd_sc_hd__nand2_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07568_ fanout85/X fanout83/X fanout82/X fanout79/X vssd1 vssd1 vccd1 vccd1 _07569_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13432__C1 _13568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09307_ _09308_/B _09308_/A vssd1 vssd1 vccd1 vccd1 _09307_/Y sky130_fd_sc_hd__nand2b_1
X_07499_ _07499_/A _07499_/B vssd1 vssd1 vccd1 vccd1 _07500_/B sky130_fd_sc_hd__or2_1
XFILLER_0_90_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09238_ _09238_/A _09238_/B vssd1 vssd1 vccd1 vccd1 _09239_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07662__B1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12538__A1 _12710_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09169_ _09169_/A _09169_/B vssd1 vssd1 vccd1 vccd1 _09184_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11200_ _11326_/D _11200_/B vssd1 vssd1 vccd1 vccd1 _11202_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_114_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12180_ _12180_/A _12180_/B vssd1 vssd1 vccd1 vccd1 _12181_/B sky130_fd_sc_hd__and2_1
X_11131_ _10192_/X _11130_/X _11576_/A vssd1 vssd1 vccd1 vccd1 _11131_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09706__A2 _12314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11062_ _11062_/A _11062_/B vssd1 vssd1 vccd1 vccd1 _11064_/B sky130_fd_sc_hd__or2_1
XFILLER_0_101_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10013_ reg1_val[3] curr_PC[3] vssd1 vssd1 vccd1 vccd1 _10016_/B sky130_fd_sc_hd__or2_1
XANTENNA__12710__B2 _12710_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11964_ reg1_val[19] curr_PC[19] vssd1 vssd1 vccd1 vccd1 _11965_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13703_ _13742_/CLK hold34/X vssd1 vssd1 vccd1 vccd1 hold123/A sky130_fd_sc_hd__dfxtp_1
X_10915_ _10915_/A _11825_/A vssd1 vssd1 vccd1 vccd1 _10917_/B sky130_fd_sc_hd__nor2_1
X_11895_ _10342_/A _11891_/X _11894_/X vssd1 vssd1 vccd1 vccd1 dest_val[18] sky130_fd_sc_hd__o21ai_4
XANTENNA__09890__A1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09890__B2 _07833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13634_ _13731_/CLK hold41/X vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__dfxtp_1
X_10846_ _10847_/A _10847_/B vssd1 vssd1 vccd1 vccd1 _10976_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12777__A1 _10734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13565_ _13565_/A _13565_/B vssd1 vssd1 vccd1 vccd1 _13565_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__08445__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10777_ _10777_/A _10777_/B vssd1 vssd1 vccd1 vccd1 _10778_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10788__B1 _07546_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12516_ _12516_/A _12516_/B vssd1 vssd1 vccd1 vccd1 _12516_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07410__B _07535_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13496_ hold280/X _13555_/A2 _13495_/X _13542_/B2 vssd1 vssd1 vccd1 vccd1 hold281/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12447_ _12373_/A _12480_/A _12373_/B _12056_/B vssd1 vssd1 vccd1 vccd1 _12447_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_112_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12378_ _12130_/A _09082_/B _09082_/C _10866_/B vssd1 vssd1 vccd1 vccd1 _12379_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_50_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11329_ _11329_/A _11329_/B vssd1 vssd1 vccd1 vccd1 _11331_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12701__A1 _12648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11504__A2 _09146_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06870_ instruction[0] instruction[1] instruction[2] instruction[31] pred_val vssd1
+ vssd1 vccd1 vccd1 _13010_/B sky130_fd_sc_hd__o311a_4
XANTENNA__06977__A _13015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07572__S _07572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09353__A _10095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08540_ _10236_/A _08540_/B vssd1 vssd1 vccd1 vccd1 _08544_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08471_ _08471_/A _08471_/B vssd1 vssd1 vccd1 vccd1 _09077_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07422_ _07422_/A _07422_/B vssd1 vssd1 vccd1 vccd1 _07422_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_9_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_358 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07353_ _07360_/A _07360_/B vssd1 vssd1 vccd1 vccd1 _11512_/A sky130_fd_sc_hd__and2_4
XFILLER_0_33_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07284_ _10366_/A _07285_/B vssd1 vssd1 vccd1 vccd1 _09929_/A sky130_fd_sc_hd__and2_1
XFILLER_0_127_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06998__A2 _06936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09023_ _09023_/A _09023_/B _09023_/C vssd1 vssd1 vccd1 vccd1 _09025_/A sky130_fd_sc_hd__and3_1
XFILLER_0_32_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold210 hold210/A vssd1 vssd1 vccd1 vccd1 hold210/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09936__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold221 hold221/A vssd1 vssd1 vccd1 vccd1 hold221/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08432__A _09373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold232 hold232/A vssd1 vssd1 vccd1 vccd1 hold232/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold243 hold243/A vssd1 vssd1 vccd1 vccd1 hold243/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 hold254/A vssd1 vssd1 vccd1 vccd1 hold254/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 hold265/A vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold276 hold301/X vssd1 vssd1 vccd1 vccd1 hold276/X sky130_fd_sc_hd__buf_1
Xhold287 hold287/A vssd1 vssd1 vccd1 vccd1 hold287/X sky130_fd_sc_hd__dlygate4sd3_1
X_09925_ _10537_/A _09925_/B vssd1 vssd1 vccd1 vccd1 _09935_/A sky130_fd_sc_hd__xnor2_2
Xhold298 hold298/A vssd1 vssd1 vccd1 vccd1 hold298/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12889__A _13048_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13496__A2 _13555_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11793__A _11793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09856_ reg1_val[2] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _09857_/B sky130_fd_sc_hd__nand2_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08372__A1 _08866_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08807_ _08857_/A _08807_/B vssd1 vssd1 vccd1 vccd1 _08845_/A sky130_fd_sc_hd__xor2_1
XANTENNA__08372__B2 _08950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09787_ _09788_/A _09788_/B vssd1 vssd1 vccd1 vccd1 _09787_/Y sky130_fd_sc_hd__nand2_1
X_06999_ _06928_/A _06936_/B _13005_/B _06997_/X vssd1 vssd1 vccd1 vccd1 _07363_/B
+ sky130_fd_sc_hd__a31oi_4
XANTENNA__11259__A1 _10603_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08738_ _10542_/A _08738_/B vssd1 vssd1 vccd1 vccd1 _08766_/A sky130_fd_sc_hd__xnor2_2
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _08951_/A _08669_/B vssd1 vssd1 vccd1 vccd1 _08715_/A sky130_fd_sc_hd__xnor2_2
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08675__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09872__B2 _12796_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _10798_/B _10701_/C vssd1 vssd1 vccd1 vccd1 _10702_/B sky130_fd_sc_hd__nand2_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ reg1_val[16] curr_PC[16] vssd1 vssd1 vccd1 vccd1 _11681_/B sky130_fd_sc_hd__nand2_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07511__A _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12759__A1 _12759_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10631_ _10631_/A _10857_/A _10981_/A _10981_/B vssd1 vssd1 vccd1 vccd1 _10631_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_76_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13420__A2 _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13350_ hold195/X _13463_/B2 _13450_/B hold231/X vssd1 vssd1 vccd1 vccd1 hold232/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10562_ _10391_/A _10391_/B _10393_/B _10394_/X vssd1 vssd1 vccd1 vccd1 _10564_/B
+ sky130_fd_sc_hd__a31oi_2
XFILLER_0_24_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12301_ _12218_/A _12215_/X _06863_/A vssd1 vssd1 vccd1 vccd1 _12301_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_63_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13281_ hold11/X hold245/X vssd1 vssd1 vccd1 vccd1 _13281_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_16_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10493_ _11913_/A _10493_/B vssd1 vssd1 vccd1 vccd1 _10495_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13184__A1 _11922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12232_ _12314_/A _12313_/B hold255/A vssd1 vssd1 vccd1 vccd1 _12234_/A sky130_fd_sc_hd__a21oi_1
X_12163_ _12163_/A _12163_/B _12163_/C vssd1 vssd1 vccd1 vccd1 _12164_/D sky130_fd_sc_hd__or3_1
X_11114_ _11114_/A _11114_/B vssd1 vssd1 vccd1 vccd1 _11115_/B sky130_fd_sc_hd__or2_2
X_12094_ _12094_/A _12094_/B vssd1 vssd1 vccd1 vccd1 _12096_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12144__C1 _09529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11045_ _11527_/A fanout16/X _07877_/X _11423_/A vssd1 vssd1 vccd1 vccd1 _11046_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07108__D _07108_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12447__B1 _12056_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12996_ _12994_/Y _12996_/B vssd1 vssd1 vccd1 vccd1 _12997_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09901__A _10266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11947_ _11947_/A vssd1 vssd1 vccd1 vccd1 _11947_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11670__A1 _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11878_ hold200/A hold231/A _11878_/C vssd1 vssd1 vccd1 vccd1 _11972_/B sky130_fd_sc_hd__or3_1
XFILLER_0_39_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13617_ _13719_/CLK _13617_/D vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__dfxtp_1
X_10829_ _10828_/B _10828_/C _10828_/A vssd1 vssd1 vccd1 vccd1 _10829_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07140__B _13748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13548_ _13548_/A _13548_/B vssd1 vssd1 vccd1 vccd1 _13548_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12981__B _12982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13479_ _13479_/A _13479_/B vssd1 vssd1 vccd1 vccd1 _13479_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11186__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08051__B1 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07971_ fanout85/X fanout68/X fanout66/X fanout82/X vssd1 vssd1 vccd1 vccd1 _07972_/B
+ sky130_fd_sc_hd__o22a_1
X_09710_ _07024_/Y _11587_/A2 _09704_/X _07026_/B _09709_/X vssd1 vssd1 vccd1 vccd1
+ _09710_/X sky130_fd_sc_hd__o221a_1
X_06922_ _07527_/A vssd1 vssd1 vccd1 vccd1 _07526_/A sky130_fd_sc_hd__inv_2
XFILLER_0_93_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09641_ _09641_/A _09641_/B vssd1 vssd1 vccd1 vccd1 _09642_/B sky130_fd_sc_hd__xor2_2
X_06853_ reg2_val[23] _07110_/A _06872_/B1 _06852_/Y vssd1 vssd1 vccd1 vccd1 _07230_/A
+ sky130_fd_sc_hd__o2bb2a_4
X_09572_ fanout51/X _10235_/A1 _10235_/B2 fanout44/X vssd1 vssd1 vccd1 vccd1 _09573_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_93_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06784_ instruction[1] instruction[2] instruction[25] pred_val vssd1 vssd1 vccd1
+ vccd1 _06784_/X sky130_fd_sc_hd__o211a_2
XFILLER_0_26_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08523_ _11286_/A _08523_/B vssd1 vssd1 vccd1 vccd1 _08607_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11110__B1 _11109_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08454_ _08454_/A _08454_/B vssd1 vssd1 vccd1 vccd1 _08455_/B sky130_fd_sc_hd__and2_1
XFILLER_0_9_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07405_ _10004_/S _09703_/B _11463_/A _07398_/B vssd1 vssd1 vccd1 vccd1 _07407_/B
+ sky130_fd_sc_hd__o211a_4
XFILLER_0_92_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08385_ _08746_/A _08385_/B vssd1 vssd1 vccd1 vccd1 _08389_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09606__A1 _09955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09606__B2 _09910_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07336_ _07377_/A _07377_/B vssd1 vssd1 vccd1 vccd1 _07336_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_61_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07267_ _13015_/A _07266_/X _07572_/S vssd1 vssd1 vccd1 vccd1 _07267_/X sky130_fd_sc_hd__mux2_2
XANTENNA__10692__A _11709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09006_ _09005_/Y _09006_/B vssd1 vssd1 vccd1 vccd1 _09994_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__13166__A1 _13166_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09258__A _09949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07198_ _07198_/A _07198_/B vssd1 vssd1 vccd1 vccd1 _07198_/Y sky130_fd_sc_hd__nand2_8
XANTENNA__11177__B1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08593__A1 _08923_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08593__B2 _08866_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09908_ _09908_/A _09908_/B vssd1 vssd1 vccd1 vccd1 _09909_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11954__C _12164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09705__B _12578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout72_A _07546_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09839_ _09839_/A _09839_/B vssd1 vssd1 vccd1 vccd1 _09839_/Y sky130_fd_sc_hd__nor2_1
X_12850_ _12851_/A _12851_/B _12851_/C vssd1 vssd1 vccd1 vccd1 _12858_/B sky130_fd_sc_hd__a21o_1
X_11801_ _07446_/Y fanout7/X _11800_/X _11913_/A vssd1 vssd1 vccd1 vccd1 _11920_/A
+ sky130_fd_sc_hd__a22o_2
X_12781_ _12781_/A _12781_/B vssd1 vssd1 vccd1 vccd1 _12781_/Y sky130_fd_sc_hd__nand2_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10867__A _12515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11732_ _11732_/A _11825_/A vssd1 vssd1 vccd1 vccd1 _11733_/B sky130_fd_sc_hd__nor2_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _11663_/A _11761_/A vssd1 vssd1 vccd1 vccd1 _11857_/A sky130_fd_sc_hd__nor2_1
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13402_ hold19/X _13416_/A2 _13420_/B1 hold157/A _13383_/A vssd1 vssd1 vccd1 vccd1
+ hold20/A sky130_fd_sc_hd__o221a_1
XANTENNA__10207__A2 _10915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10614_ _06979_/B _11587_/A2 _10607_/Y _06977_/Y _10613_/X vssd1 vssd1 vccd1 vccd1
+ _10614_/X sky130_fd_sc_hd__o221a_1
XANTENNA__11404__A1 _07282_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11404__B2 _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11594_ _09529_/B _11578_/X _11593_/X _11569_/X vssd1 vssd1 vccd1 vccd1 _11594_/X
+ sky130_fd_sc_hd__o211a_1
X_13333_ _13359_/A _13333_/B vssd1 vssd1 vccd1 vccd1 _13648_/D sky130_fd_sc_hd__and2_1
X_10545_ _10544_/B _10544_/C _10544_/A vssd1 vssd1 vccd1 vccd1 _10546_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_122_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13264_ hold295/A hold111/X vssd1 vssd1 vccd1 vccd1 _13488_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10476_ _12759_/A1 _12462_/B _10458_/X _10321_/X _10475_/Y vssd1 vssd1 vccd1 vccd1
+ _10476_/X sky130_fd_sc_hd__a221o_1
XANTENNA__11168__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12215_ _12136_/A _12133_/X _06876_/A vssd1 vssd1 vccd1 vccd1 _12215_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_122_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10107__A _10522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13195_ hold39/X _13207_/B vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__or2_1
XFILLER_0_121_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09781__B1 _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09526__A1_N _09501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12146_ _12058_/A _12231_/B hold266/A vssd1 vssd1 vccd1 vccd1 _12146_/Y sky130_fd_sc_hd__a21oi_1
X_12077_ _07230_/Y fanout8/X fanout3/X _12189_/A vssd1 vssd1 vccd1 vccd1 _12078_/B
+ sky130_fd_sc_hd__a22o_1
X_11028_ _11029_/A _11029_/B _11029_/C vssd1 vssd1 vccd1 vccd1 _11209_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12979_ _12979_/A _12979_/B vssd1 vssd1 vccd1 vccd1 _12980_/B sky130_fd_sc_hd__xor2_2
XANTENNA__06974__B _06980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08247__A _10266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12992__A _12992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_16 instruction[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_27 reg1_val[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_38 reg1_val[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08170_ _08232_/A _08232_/B vssd1 vssd1 vccd1 vccd1 _08236_/A sky130_fd_sc_hd__or2_1
XANTENNA_49 reg2_val[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07121_ instruction[12] _07122_/B vssd1 vssd1 vccd1 vccd1 dest_pred[1] sky130_fd_sc_hd__and2_4
XFILLER_0_27_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07150__A_N _13744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07052_ reg1_val[23] _07230_/A vssd1 vssd1 vccd1 vccd1 _07052_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_2_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10017__A _12648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10906__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08710__A _09950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07954_ _07954_/A _07954_/B vssd1 vssd1 vccd1 vccd1 _07956_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06905_ _06928_/B _12806_/A vssd1 vssd1 vccd1 vccd1 _06905_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13047__B _13048_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07885_ fanout51/X _08866_/B2 _08950_/B fanout44/X vssd1 vssd1 vccd1 vccd1 _07886_/B
+ sky130_fd_sc_hd__o22a_1
X_09624_ _09625_/A _09625_/B vssd1 vssd1 vccd1 vccd1 _09624_/X sky130_fd_sc_hd__and2_1
X_06836_ reg1_val[26] _07252_/C vssd1 vssd1 vccd1 vccd1 _06840_/A sky130_fd_sc_hd__nand2_2
X_09555_ _09555_/A _09555_/B vssd1 vssd1 vccd1 vccd1 _09557_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06767_ instruction[23] instruction[16] _07135_/S vssd1 vssd1 vccd1 vccd1 reg1_idx[5]
+ sky130_fd_sc_hd__mux2_8
XANTENNA__09827__A1 _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08506_ _08506_/A _08506_/B vssd1 vssd1 vccd1 vccd1 _08574_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11634__A1 _10944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09486_ reg1_val[3] reg1_val[28] _09493_/S vssd1 vssd1 vccd1 vccd1 _09486_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08437_ _08504_/A _08504_/B vssd1 vssd1 vccd1 vccd1 _08505_/A sky130_fd_sc_hd__and2_1
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08368_ _08368_/A _08368_/B vssd1 vssd1 vccd1 vccd1 _08370_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11014__C _11014_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07319_ _13015_/A reg1_val[10] _07320_/C _07320_/D vssd1 vssd1 vccd1 vccd1 _07571_/A
+ sky130_fd_sc_hd__nor4_4
XANTENNA__08263__B1 _13168_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08299_ _08299_/A _08299_/B vssd1 vssd1 vccd1 vccd1 _08365_/B sky130_fd_sc_hd__or2_1
XFILLER_0_61_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10330_ _06994_/A _11587_/A2 _10324_/Y _06996_/B _10329_/X vssd1 vssd1 vccd1 vccd1
+ _10330_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_0_21_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10261_ _10275_/A vssd1 vssd1 vccd1 vccd1 _10261_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_103_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07369__A2 fanout39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12000_ _12000_/A _12000_/B vssd1 vssd1 vccd1 vccd1 _12001_/B sky130_fd_sc_hd__nand2_1
X_10192_ _11472_/S _10008_/X _09534_/C vssd1 vssd1 vccd1 vccd1 _10192_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07236__A _08951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12902_ reg1_val[15] curr_PC[15] _12978_/S vssd1 vssd1 vccd1 vccd1 _12904_/B sky130_fd_sc_hd__mux2_1
X_12833_ _13005_/B _12834_/B vssd1 vssd1 vccd1 vccd1 _12844_/A sky130_fd_sc_hd__nand2_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13075__B1 _13129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11625__A1 _07230_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ fanout5/X _12764_/B vssd1 vssd1 vccd1 vccd1 _12768_/A sky130_fd_sc_hd__nand2_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11625__B2 _12331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11715_ _12331_/A fanout15/X fanout31/X _12413_/A vssd1 vssd1 vccd1 vccd1 _11716_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ _12695_/A _12695_/B vssd1 vssd1 vccd1 vccd1 _12695_/X sky130_fd_sc_hd__and2_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11646_ _11646_/A _11646_/B _11646_/C _11646_/D vssd1 vssd1 vccd1 vccd1 _11647_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_52_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09451__C1 _10457_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11577_ _10458_/S _11575_/X _11576_/X vssd1 vssd1 vccd1 vccd1 _11577_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_3_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13316_ hold233/X hold172/X vssd1 vssd1 vccd1 vccd1 _13316_/Y sky130_fd_sc_hd__nand2b_1
X_10528_ _07472_/Y fanout16/X _07877_/X _10915_/A vssd1 vssd1 vccd1 vccd1 _10529_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13247_ _13247_/A _13247_/B vssd1 vssd1 vccd1 vccd1 _13527_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10459_ hold182/A hold238/A _10459_/C vssd1 vssd1 vccd1 vccd1 _10604_/B sky130_fd_sc_hd__or3_1
XFILLER_0_20_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13178_ _11638_/A _13194_/A2 hold127/X _13539_/A vssd1 vssd1 vccd1 vccd1 _13625_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08530__A _09950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10364__A1 _10536_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10364__B2 _10536_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12129_ _12129_/A _12164_/C vssd1 vssd1 vccd1 vccd1 _12129_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07146__A _12971_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10116__A1 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10116__B2 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07670_ _07749_/A _07669_/Y _07668_/A vssd1 vssd1 vccd1 vccd1 _07686_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09361__A _09591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09340_ _09340_/A _09340_/B vssd1 vssd1 vccd1 vccd1 _09342_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09271_ _09151_/A _09151_/B _09149_/Y vssd1 vssd1 vccd1 vccd1 _09275_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__11115__B _11115_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08222_ _08222_/A _08222_/B vssd1 vssd1 vccd1 vccd1 _08229_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_90_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08153_ _08222_/A _08222_/B _08132_/X vssd1 vssd1 vccd1 vccd1 _08162_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12041__A1 _12695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08796__A1 _09501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10052__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07104_ instruction[5] _07104_/B vssd1 vssd1 vccd1 vccd1 dest_pred_val sky130_fd_sc_hd__xnor2_4
XANTENNA__08796__B2 _08271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09993__B1 _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08084_ _10266_/A _08084_/B vssd1 vssd1 vccd1 vccd1 _08112_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07035_ _07000_/Y _07034_/X _10311_/A vssd1 vssd1 vccd1 vccd1 _10447_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06879__B _13000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07220__A1 _07213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10181__S _12648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ _09068_/A _09077_/B _08568_/Y vssd1 vssd1 vccd1 vccd1 _08988_/B sky130_fd_sc_hd__or3b_1
XANTENNA__09760__A3 _10787_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07937_ _07937_/A _07937_/B vssd1 vssd1 vccd1 vccd1 _07938_/B sky130_fd_sc_hd__or2_1
XANTENNA__12897__A _13054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11304__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07868_ _07637_/B _07866_/X _07865_/X vssd1 vssd1 vccd1 vccd1 _07868_/Y sky130_fd_sc_hd__o21ai_2
X_09607_ _10522_/B _09607_/B vssd1 vssd1 vccd1 vccd1 _09609_/B sky130_fd_sc_hd__xnor2_1
X_06819_ _06817_/Y _06872_/B1 _06873_/B1 reg2_val[28] vssd1 vssd1 vccd1 vccd1 _09254_/C
+ sky130_fd_sc_hd__a2bb2o_2
X_07799_ _08821_/B2 fanout42/X fanout40/X _08821_/A1 vssd1 vssd1 vccd1 vccd1 _07800_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12804__A0 _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09538_ _09499_/Y _09860_/A _12783_/A _09839_/A _09528_/X vssd1 vssd1 vccd1 vccd1
+ _09538_/X sky130_fd_sc_hd__o221a_1
XANTENNA__10210__A _12253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09469_ _09467_/X _09468_/X _09688_/S vssd1 vssd1 vccd1 vccd1 _09469_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_66_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11500_ _11922_/A _07643_/B fanout12/X wire101/X vssd1 vssd1 vccd1 vccd1 _11501_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12480_ _12480_/A _12480_/B vssd1 vssd1 vccd1 vccd1 _12635_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_81_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11431_ _11431_/A _11431_/B vssd1 vssd1 vccd1 vccd1 _11445_/A sky130_fd_sc_hd__and2_1
XFILLER_0_123_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10043__B1 _12825_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11362_ _11362_/A _11362_/B vssd1 vssd1 vccd1 vccd1 _11362_/X sky130_fd_sc_hd__xor2_1
X_13101_ _13101_/A _13106_/A vssd1 vssd1 vccd1 vccd1 _13105_/A sky130_fd_sc_hd__nand2_2
XANTENNA__11791__B1 _11774_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10313_ _10313_/A vssd1 vssd1 vccd1 vccd1 _10313_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10880__A _12648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11293_ _12093_/A _11293_/B vssd1 vssd1 vccd1 vccd1 _11301_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08539__A1 _08891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13032_ _13033_/A _13033_/C _13033_/B vssd1 vssd1 vccd1 vccd1 _13039_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08539__B2 _08873_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ _10244_/A vssd1 vssd1 vccd1 vccd1 _10252_/A sky130_fd_sc_hd__inv_2
X_10175_ _11575_/S _10171_/X _10174_/Y _11576_/A vssd1 vssd1 vccd1 vccd1 _10175_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07762__A2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout180 _07163_/X vssd1 vssd1 vccd1 vccd1 _09373_/A sky130_fd_sc_hd__buf_8
XANTENNA__10104__B _10518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout191 _12796_/A1 vssd1 vssd1 vccd1 vccd1 _12748_/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12816_ _12816_/A _12816_/B _12816_/C vssd1 vssd1 vccd1 vccd1 _12817_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_84_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _12786_/B1 _12746_/X hold233/A vssd1 vssd1 vccd1 vccd1 _12749_/A sky130_fd_sc_hd__a21oi_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12678_ _12677_/A _12677_/B _12677_/C vssd1 vssd1 vccd1 vccd1 _12731_/A sky130_fd_sc_hd__o21a_1
XANTENNA__08525__A _09591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11629_ _11743_/A _11629_/B vssd1 vssd1 vccd1 vccd1 _11631_/B sky130_fd_sc_hd__or2_1
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10034__B1 _12657_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11782__B1 _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10790__A _11286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09727__B1 _09885_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10337__A1 _10320_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10337__B2 _09523_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _08843_/B _08843_/C _08843_/A vssd1 vssd1 vccd1 vccd1 _08844_/A sky130_fd_sc_hd__o21ai_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07202__A1 _07213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _08774_/A _08774_/B vssd1 vssd1 vccd1 vccd1 _08771_/X sky130_fd_sc_hd__and2_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07722_ _07656_/A _07722_/B vssd1 vssd1 vccd1 vccd1 _07744_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__08702__A1 _08873_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08702__B2 _13149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07653_ _07653_/A _07653_/B vssd1 vssd1 vccd1 vccd1 _07659_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_95_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11126__A _11126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07584_ _07584_/A _07584_/B vssd1 vssd1 vccd1 vccd1 _07696_/B sky130_fd_sc_hd__or2_1
XFILLER_0_87_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09323_ _09313_/A _09313_/B _09201_/X vssd1 vssd1 vccd1 vccd1 _09828_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_47_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09254_ _09254_/A _09254_/B _09254_/C _09254_/D vssd1 vssd1 vccd1 vccd1 _09254_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_16_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08435__A _10236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08205_ _08205_/A _08205_/B _08205_/C vssd1 vssd1 vccd1 vccd1 _08257_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09185_ _09185_/A _09185_/B vssd1 vssd1 vccd1 vccd1 _09186_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_7_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08769__A1 _08821_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08769__B2 _08821_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08136_ _08873_/A2 fanout76/X fanout74/X _08891_/B vssd1 vssd1 vccd1 vccd1 _08137_/B
+ sky130_fd_sc_hd__o22a_1
X_08067_ _08133_/A _08133_/B _08063_/Y vssd1 vssd1 vccd1 vccd1 _08156_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_113_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12317__A2 _12799_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07018_ reg2_val[1] _07110_/A vssd1 vssd1 vccd1 vccd1 _07025_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_113_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08941__A1 _08271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08941__B2 _09501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ _08970_/A _08970_/B _09019_/A vssd1 vssd1 vccd1 vccd1 _08971_/B sky130_fd_sc_hd__a21o_1
X_11980_ _11980_/A _11980_/B _11980_/C vssd1 vssd1 vccd1 vccd1 _11980_/X sky130_fd_sc_hd__or3_1
XANTENNA__12420__A _12420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10931_ _10931_/A _10931_/B vssd1 vssd1 vccd1 vccd1 _10932_/B sky130_fd_sc_hd__and2_1
XFILLER_0_98_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11036__A _11719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10862_ _12742_/A _10900_/A _10900_/B vssd1 vssd1 vccd1 vccd1 _10863_/B sky130_fd_sc_hd__or3_1
X_13650_ _13659_/CLK hold165/X vssd1 vssd1 vccd1 vccd1 hold240/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _06801_/Y _09516_/X _12599_/Y _06802_/A _12600_/X vssd1 vssd1 vccd1 vccd1
+ _12601_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_94_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11056__A2 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13581_ hold247/X _13580_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13581_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10793_ _10791_/X _10793_/B vssd1 vssd1 vccd1 vccd1 _10794_/B sky130_fd_sc_hd__and2b_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12532_ _12374_/A _12592_/B hold166/A vssd1 vssd1 vccd1 vccd1 _12532_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08209__B1 _08778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12463_ _12782_/B _12461_/Y _12462_/Y _09529_/B vssd1 vssd1 vccd1 vccd1 _12475_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__12005__A1 _12331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12005__B2 _07230_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09957__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11414_ _11415_/A _11415_/B vssd1 vssd1 vccd1 vccd1 _11538_/A sky130_fd_sc_hd__nor2_1
X_12394_ _12374_/A _12467_/B hold216/A vssd1 vssd1 vccd1 vccd1 _12394_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11345_ _11109_/Y _11556_/A _11344_/Y vssd1 vssd1 vccd1 vccd1 _11345_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07983__A2 _08907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11276_ _07310_/Y fanout34/X fanout32/X _07282_/X vssd1 vssd1 vccd1 vccd1 _11277_/B
+ sky130_fd_sc_hd__o22a_1
X_13015_ _13015_/A _13015_/B vssd1 vssd1 vccd1 vccd1 _13016_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_120_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10227_ _11823_/A _10227_/B vssd1 vssd1 vccd1 vccd1 _10229_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13686__CLK _13701_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07735__A2 _10536_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10158_ _10045_/X _10200_/B _10157_/Y vssd1 vssd1 vccd1 vccd1 _10158_/Y sky130_fd_sc_hd__a21oi_1
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__buf_1
X_10089_ _11281_/A _10089_/B vssd1 vssd1 vccd1 vccd1 _10091_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07424__A _12421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13145__B _13193_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07423__A1 _09910_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07423__B2 _07833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09941_ fanout53/X fanout75/X _08704_/B fanout47/X vssd1 vssd1 vccd1 vccd1 _09942_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07318__B _07535_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ reg1_val[2] _11688_/B _09870_/Y _12796_/A1 _09871_/Y vssd1 vssd1 vccd1 vccd1
+ _09872_/X sky130_fd_sc_hd__o221a_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08923__A1 _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _08271_/A _07492_/Y _10637_/A _09501_/A vssd1 vssd1 vccd1 vccd1 _08824_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08923__B2 _08907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08754_ _08790_/A _08790_/B _08747_/Y vssd1 vssd1 vccd1 vccd1 _08762_/A sky130_fd_sc_hd__o21a_1
X_07705_ _07717_/A _07717_/B vssd1 vssd1 vccd1 vccd1 _07718_/A sky130_fd_sc_hd__nand2_1
X_08685_ _08685_/A _08685_/B vssd1 vssd1 vccd1 vccd1 _08687_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12483__A1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12483__B2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07636_ _12656_/A _12656_/B _07637_/B vssd1 vssd1 vccd1 vccd1 _07641_/C sky130_fd_sc_hd__a21o_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07567_ _07948_/A _07567_/B vssd1 vssd1 vccd1 vccd1 _07588_/A sky130_fd_sc_hd__or2_1
XANTENNA__13432__B1 _13444_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09306_ _09306_/A _09306_/B vssd1 vssd1 vccd1 vccd1 _09308_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_76_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07498_ _07499_/A _07499_/B vssd1 vssd1 vccd1 vccd1 _07500_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_36_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09237_ _09238_/A _09238_/B vssd1 vssd1 vccd1 vccd1 _09237_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07662__A1 _11047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07662__B2 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09939__B1 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12538__A2 _10320_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09168_ _09168_/A _09168_/B vssd1 vssd1 vccd1 vccd1 _09169_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_50_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08119_ _08933_/B _07300_/Y _11638_/A _07175_/X vssd1 vssd1 vccd1 vccd1 _08120_/B
+ sky130_fd_sc_hd__a22o_1
X_09099_ _07959_/A _07959_/B _07957_/X vssd1 vssd1 vccd1 vccd1 _09203_/A sky130_fd_sc_hd__a21oi_4
X_11130_ _10002_/X _10006_/X _11575_/S vssd1 vssd1 vccd1 vccd1 _11130_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_101_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11061_ _11061_/A _11061_/B vssd1 vssd1 vccd1 vccd1 _11062_/B sky130_fd_sc_hd__and2_1
X_10012_ reg1_val[3] curr_PC[3] vssd1 vssd1 vccd1 vccd1 _10012_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07244__A _08951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11963_ reg1_val[19] curr_PC[19] vssd1 vssd1 vccd1 vccd1 _11965_/A sky130_fd_sc_hd__or2_1
XFILLER_0_58_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13702_ _13705_/CLK _13702_/D vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__dfxtp_1
X_10914_ _10914_/A _10914_/B vssd1 vssd1 vccd1 vccd1 _10917_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_98_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11894_ _12327_/A _11894_/B _12070_/C vssd1 vssd1 vccd1 vccd1 _11894_/X sky130_fd_sc_hd__or3_1
XANTENNA__09890__A2 _07455_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10845_ _10845_/A _10845_/B vssd1 vssd1 vccd1 vccd1 _10847_/B sky130_fd_sc_hd__xnor2_1
X_13633_ _13731_/CLK _13633_/D vssd1 vssd1 vccd1 vccd1 hold118/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10237__B1 _12667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08075__A _11286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10776_ _10776_/A _10776_/B vssd1 vssd1 vccd1 vccd1 _10777_/B sky130_fd_sc_hd__or2_1
X_13564_ _13591_/A hold279/X vssd1 vssd1 vccd1 vccd1 _13730_/D sky130_fd_sc_hd__and2_1
XANTENNA__11985__B1 _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12515_ _07079_/Y _12514_/Y _12515_/S vssd1 vssd1 vccd1 vccd1 _12516_/B sky130_fd_sc_hd__mux2_1
X_13495_ hold253/X _13494_/Y hold234/X vssd1 vssd1 vccd1 vccd1 _13495_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_109_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12446_ _12570_/A _12446_/B vssd1 vssd1 vccd1 vccd1 _12480_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_35_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07405__A1 _10004_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12377_ _12130_/A _09082_/B _09082_/C vssd1 vssd1 vccd1 vccd1 _12379_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11328_ _11329_/A _11329_/B vssd1 vssd1 vccd1 vccd1 _11440_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09158__A1 _13129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11259_ _10603_/S _10009_/X _09537_/B vssd1 vssd1 vccd1 vccd1 _11259_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_120_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06977__B _07492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07154__A _12578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08470_ _08470_/A _08470_/B vssd1 vssd1 vccd1 vccd1 _09068_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_77_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07421_ _07422_/A _07422_/B vssd1 vssd1 vccd1 vccd1 _07421_/X sky130_fd_sc_hd__and2_2
XANTENNA__13701__CLK _13701_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07352_ _07351_/A _07351_/B _07637_/B vssd1 vssd1 vccd1 vccd1 _07360_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_17_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07283_ _07283_/A _07283_/B vssd1 vssd1 vccd1 vccd1 _11922_/A sky130_fd_sc_hd__nand2_8
XFILLER_0_5_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09022_ _09019_/A _09019_/B _08882_/X _08900_/X vssd1 vssd1 vccd1 vccd1 _09023_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_115_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06998__A3 _13005_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11728__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold200 hold200/A vssd1 vssd1 vccd1 vccd1 hold200/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold211 hold211/A vssd1 vssd1 vccd1 vccd1 hold211/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_4_3_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13708_/CLK sky130_fd_sc_hd__clkbuf_8
Xhold222 hold237/X vssd1 vssd1 vccd1 vccd1 hold222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 hold233/A vssd1 vssd1 vccd1 vccd1 hold233/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10400__B1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold244 hold244/A vssd1 vssd1 vccd1 vccd1 hold244/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 hold255/A vssd1 vssd1 vccd1 vccd1 hold255/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 hold266/A vssd1 vssd1 vccd1 vccd1 hold266/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold277 hold277/A vssd1 vssd1 vccd1 vccd1 hold277/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 hold288/A vssd1 vssd1 vccd1 vccd1 hold288/X sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ _12496_/A _10536_/A1 _10536_/B2 _07257_/X vssd1 vssd1 vccd1 vccd1 _09925_/B
+ sky130_fd_sc_hd__a22o_1
Xhold299 hold299/A vssd1 vssd1 vccd1 vccd1 hold299/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11793__B _11793_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09855_ reg1_val[2] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _09855_/Y sky130_fd_sc_hd__nor2_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06907__B1 _06980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11900__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08372__A2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08806_ _09703_/B _08806_/A2 _08806_/B1 _07399_/Y vssd1 vssd1 vccd1 vccd1 _08807_/B
+ sky130_fd_sc_hd__a22o_1
X_09786_ _09786_/A _09786_/B vssd1 vssd1 vccd1 vccd1 _09788_/B sky130_fd_sc_hd__xnor2_2
X_06998_ _06928_/A _06936_/B _13005_/B _06997_/X vssd1 vssd1 vccd1 vccd1 _06998_/X
+ sky130_fd_sc_hd__a31o_1
X_08737_ _08873_/A2 _08866_/A2 _09216_/B2 _08891_/B vssd1 vssd1 vccd1 vccd1 _08738_/B
+ sky130_fd_sc_hd__o22a_1
X_08668_ _08866_/B2 _10049_/A2 _09173_/B2 _08950_/B vssd1 vssd1 vccd1 vccd1 _08669_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09872__A2 _11688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07619_ _07672_/A _07619_/B vssd1 vssd1 vccd1 vccd1 _07620_/B sky130_fd_sc_hd__xnor2_2
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08599_ _08857_/A _08599_/B vssd1 vssd1 vccd1 vccd1 _08647_/A sky130_fd_sc_hd__xnor2_2
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10630_ _10438_/A _10629_/Y _10628_/Y vssd1 vssd1 vccd1 vccd1 _10630_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12129__B _12164_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10561_ _10383_/A _10383_/B _10381_/Y vssd1 vssd1 vccd1 vccd1 _10564_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_8_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12300_ _12218_/A _12216_/X _07053_/Y _12578_/A vssd1 vssd1 vccd1 vccd1 _12300_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13280_ hold262/X hold9/X vssd1 vssd1 vccd1 vccd1 _13455_/B sky130_fd_sc_hd__nand2b_1
X_10492_ _12087_/A fanout29/X fanout27/X _12103_/A vssd1 vssd1 vccd1 vccd1 _10493_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12231_ hold266/A _12231_/B vssd1 vssd1 vccd1 vccd1 _12313_/B sky130_fd_sc_hd__or2_1
XFILLER_0_121_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13184__A2 _13194_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12392__B1 _12748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12162_ _12406_/B1 _12159_/X _12325_/C _12161_/Y vssd1 vssd1 vccd1 vccd1 dest_val[21]
+ sky130_fd_sc_hd__o22ai_4
XFILLER_0_102_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11113_ _11342_/A _11113_/B _11113_/C vssd1 vssd1 vccd1 vccd1 _11114_/B sky130_fd_sc_hd__and3_1
X_12093_ _12093_/A _12094_/B vssd1 vssd1 vccd1 vccd1 _12187_/A sky130_fd_sc_hd__nand2_1
X_11044_ _11802_/B _11044_/B vssd1 vssd1 vccd1 vccd1 _11050_/A sky130_fd_sc_hd__xnor2_1
X_12995_ reg1_val[3] _12995_/B vssd1 vssd1 vccd1 vccd1 _12996_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_59_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11946_ _11757_/Y _11852_/Y _11854_/B vssd1 vssd1 vccd1 vccd1 _11947_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_86_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11877_ _11377_/Y _11876_/X _12525_/A vssd1 vssd1 vccd1 vccd1 _11877_/X sky130_fd_sc_hd__mux2_1
X_13616_ _13731_/CLK hold75/X vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__dfxtp_1
X_10828_ _10828_/A _10828_/B _10828_/C vssd1 vssd1 vccd1 vccd1 _10964_/B sky130_fd_sc_hd__or3_1
XFILLER_0_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08823__B1 _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13547_ _13547_/A hold267/X vssd1 vssd1 vccd1 vccd1 _13726_/D sky130_fd_sc_hd__and2_1
X_10759_ _12537_/B2 _10744_/X _10758_/X _12710_/B2 _10757_/X vssd1 vssd1 vccd1 vccd1
+ _10759_/X sky130_fd_sc_hd__a221o_1
XANTENNA__12981__C _12981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10630__B1 _10628_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13478_ _13267_/X _13478_/B vssd1 vssd1 vccd1 vccd1 _13479_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_23_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12429_ _12429_/A _12429_/B vssd1 vssd1 vccd1 vccd1 _12431_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11186__A1 _11638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11186__B2 _11527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07149__A _13744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11894__A _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07970_ _07970_/A _07970_/B vssd1 vssd1 vccd1 vccd1 _07991_/A sky130_fd_sc_hd__xor2_1
X_06921_ _06936_/A _06936_/B _13059_/B _06920_/X vssd1 vssd1 vccd1 vccd1 _07527_/A
+ sky130_fd_sc_hd__a31o_4
X_09640_ _09641_/A _09641_/B vssd1 vssd1 vccd1 vccd1 _09640_/Y sky130_fd_sc_hd__nor2_1
X_06852_ _06928_/B _13020_/B vssd1 vssd1 vccd1 vccd1 _06852_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10303__A _10857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09571_ _09579_/A vssd1 vssd1 vccd1 vccd1 _09571_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06783_ instruction[25] _12981_/C vssd1 vssd1 vccd1 vccd1 _12982_/B sky130_fd_sc_hd__and2_2
X_08522_ _09910_/A1 _07541_/X _07545_/Y _07420_/Y vssd1 vssd1 vccd1 vccd1 _08523_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11110__A1 _10854_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08708__A _09371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07612__A _09575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08453_ _08453_/A _08453_/B vssd1 vssd1 vccd1 vccd1 _08456_/A sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout152_A _13147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07404_ _07425_/A _07425_/B vssd1 vssd1 vccd1 vccd1 _07504_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_92_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08384_ _10522_/A _10538_/A _08778_/B _09885_/B1 vssd1 vssd1 vccd1 vccd1 _08385_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09606__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07335_ reg1_val[22] reg1_val[23] _13082_/B _07339_/D vssd1 vssd1 vccd1 vccd1 _07634_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_0_33_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07266_ _13015_/A _07320_/C vssd1 vssd1 vccd1 vccd1 _07266_/X sky130_fd_sc_hd__xor2_2
XANTENNA__08443__A _09591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09005_ _09005_/A _09005_/B vssd1 vssd1 vccd1 vccd1 _09005_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13166__A2 _13194_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07197_ _07198_/A _07198_/B vssd1 vssd1 vccd1 vccd1 _07197_/X sky130_fd_sc_hd__and2_1
XANTENNA__11177__A1 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11177__B2 _12557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08593__A2 _10538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09274__A _09275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09907_ _09907_/A _09907_/B vssd1 vssd1 vccd1 vccd1 _09908_/B sky130_fd_sc_hd__or2_1
XANTENNA__10688__B1 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11309__A _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09838_ _09839_/B vssd1 vssd1 vccd1 vccd1 _09838_/Y sky130_fd_sc_hd__inv_2
X_09769_ _11732_/A fanout24/X _08486_/B _10814_/A1 vssd1 vssd1 vccd1 vccd1 _09770_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12839__S _12867_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11800_ _11800_/A fanout5/X vssd1 vssd1 vccd1 vccd1 _11800_/X sky130_fd_sc_hd__or2_1
X_12780_ _12780_/A _12780_/B vssd1 vssd1 vccd1 vccd1 _12781_/B sky130_fd_sc_hd__xnor2_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _11731_/A _11731_/B vssd1 vssd1 vccd1 vccd1 _11733_/A sky130_fd_sc_hd__xnor2_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11044__A _11802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11662_ _11450_/A _11550_/Y _11552_/B vssd1 vssd1 vccd1 vccd1 _11662_/X sky130_fd_sc_hd__o21a_1
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13401_ _10537_/A _13419_/A2 hold65/X vssd1 vssd1 vccd1 vccd1 _13682_/D sky130_fd_sc_hd__o21a_1
X_10613_ _10611_/Y _10612_/X _10609_/X vssd1 vssd1 vccd1 vccd1 _10613_/X sky130_fd_sc_hd__o21ba_1
X_11593_ _09860_/A _11577_/Y _11592_/Y _09493_/S _11590_/X vssd1 vssd1 vccd1 vccd1
+ _11593_/X sky130_fd_sc_hd__o221a_1
XANTENNA__11404__A2 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10544_ _10544_/A _10544_/B _10544_/C vssd1 vssd1 vccd1 vccd1 _10546_/B sky130_fd_sc_hd__nand3_2
X_13332_ hold222/X _13506_/B2 _13506_/A2 hold180/X vssd1 vssd1 vccd1 vccd1 _13333_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10612__B1 _12748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08281__A1 _10266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10475_ _10460_/Y _10461_/X _10474_/X vssd1 vssd1 vccd1 vccd1 _10475_/Y sky130_fd_sc_hd__o21ai_1
X_13263_ hold111/X hold295/A vssd1 vssd1 vccd1 vccd1 _13263_/X sky130_fd_sc_hd__and2b_1
XANTENNA__11168__A1 _12103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11168__B2 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12214_ _12214_/A _12214_/B vssd1 vssd1 vccd1 vccd1 _12214_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13194_ _12331_/A _13194_/A2 hold119/X _13591_/A vssd1 vssd1 vccd1 vccd1 _13633_/D
+ sky130_fd_sc_hd__o211a_1
X_12145_ hold275/A _12145_/B vssd1 vssd1 vccd1 vccd1 _12231_/B sky130_fd_sc_hd__or2_1
XFILLER_0_20_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12076_ _12668_/A _12076_/B vssd1 vssd1 vccd1 vccd1 _12085_/A sky130_fd_sc_hd__xnor2_1
X_11027_ _11027_/A _11027_/B vssd1 vssd1 vccd1 vccd1 _11029_/C sky130_fd_sc_hd__xor2_1
XANTENNA__08528__A _09373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12978_ reg1_val[27] curr_PC[27] _12978_/S vssd1 vssd1 vccd1 vccd1 _12979_/B sky130_fd_sc_hd__mux2_2
XANTENNA__13153__B _13193_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11929_ _11929_/A _11929_/B vssd1 vssd1 vccd1 vccd1 _11931_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_74_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07151__B _13748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_17 instruction[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 reg1_val[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13396__A2 _13141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_39 reg1_val[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07120_ instruction[11] _07122_/B vssd1 vssd1 vccd1 vccd1 dest_pred[0] sky130_fd_sc_hd__and2_4
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07051_ _07050_/A _07050_/B _07099_/B vssd1 vssd1 vccd1 vccd1 _07059_/A sky130_fd_sc_hd__o21bai_1
XANTENNA__13148__A2 _13193_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_646 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10906__A1 _07526_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10906__B2 _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07607__A _10078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07953_ _07783_/A _07783_/B _07781_/X vssd1 vssd1 vccd1 vccd1 _07954_/B sky130_fd_sc_hd__a21oi_4
X_06904_ instruction[26] _12981_/C vssd1 vssd1 vccd1 vccd1 _12985_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11129__A _12648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13320__A2 _13463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07884_ _07884_/A _07884_/B vssd1 vssd1 vccd1 vccd1 _07929_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09623_ _10263_/A _09623_/B vssd1 vssd1 vccd1 vccd1 _09625_/B sky130_fd_sc_hd__xnor2_1
X_06835_ _06833_/Y _06872_/B1 _06873_/B1 reg2_val[26] vssd1 vssd1 vccd1 vccd1 _07252_/C
+ sky130_fd_sc_hd__a2bb2o_4
X_09554_ _09555_/A _09555_/B vssd1 vssd1 vccd1 vccd1 _09554_/Y sky130_fd_sc_hd__nand2_1
X_06766_ instruction[0] pred_val instruction[2] _06775_/B vssd1 vssd1 vccd1 vccd1
+ _07135_/S sky130_fd_sc_hd__and4_4
XANTENNA__09827__A2 _09650_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08505_ _08505_/A _08505_/B vssd1 vssd1 vccd1 vccd1 _08507_/B sky130_fd_sc_hd__or2_1
XANTENNA__13063__B _13129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10179__S _10457_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09485_ reg1_val[2] reg1_val[29] _09839_/A vssd1 vssd1 vccd1 vccd1 _09485_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_13_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08436_ _08436_/A _08436_/B vssd1 vssd1 vccd1 vccd1 _08504_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_108_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08367_ _08367_/A _08367_/B vssd1 vssd1 vccd1 vccd1 _08370_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_19_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07488__S _12093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07318_ _07334_/B _07535_/B vssd1 vssd1 vccd1 vccd1 _07414_/A sky130_fd_sc_hd__nand2_2
XANTENNA__08263__A1 _08806_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08263__B2 _08806_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08298_ _08299_/A _08299_/B vssd1 vssd1 vccd1 vccd1 _08298_/X sky130_fd_sc_hd__and2_1
XFILLER_0_103_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07249_ _08821_/B2 fanout53/X fanout47/X _08821_/A1 vssd1 vssd1 vccd1 vccd1 _07250_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10208__A _11719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10260_ _10058_/A _10058_/B _10056_/Y vssd1 vssd1 vccd1 vccd1 _10275_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__09212__B1 _10349_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ _07003_/B _11587_/A2 _10185_/Y _07001_/Y _10190_/X vssd1 vssd1 vccd1 vccd1
+ _10191_/X sky130_fd_sc_hd__o221a_1
XANTENNA__09732__A _12092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12901_ _12907_/B _12901_/B vssd1 vssd1 vccd1 vccd1 new_PC[14] sky130_fd_sc_hd__and2_4
XANTENNA__06962__A_N _10889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ reg1_val[5] curr_PC[5] _12867_/S vssd1 vssd1 vccd1 vccd1 _12834_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_69_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13075__B2 _07435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _12732_/Y _12733_/X _12374_/A vssd1 vssd1 vccd1 vccd1 _12763_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11625__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _11714_/A _11714_/B vssd1 vssd1 vccd1 vccd1 _11727_/A sky130_fd_sc_hd__xnor2_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _12693_/A _12693_/B _12693_/Y _09506_/X vssd1 vssd1 vccd1 vccd1 _12714_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11645_ _11646_/A _11646_/B _11646_/C _11646_/D vssd1 vssd1 vccd1 vccd1 _11647_/A
+ sky130_fd_sc_hd__o22ai_1
XFILLER_0_25_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11576_ _11576_/A _11576_/B vssd1 vssd1 vccd1 vccd1 _11576_/X sky130_fd_sc_hd__or2_1
X_13315_ hold172/X hold233/X vssd1 vssd1 vccd1 vccd1 _13315_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_122_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10527_ _12421_/A _10527_/B vssd1 vssd1 vccd1 vccd1 _10531_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10458_ _10455_/X _10457_/X _10458_/S vssd1 vssd1 vccd1 vccd1 _10458_/X sky130_fd_sc_hd__mux2_1
X_13246_ hold292/A hold55/X vssd1 vssd1 vccd1 vccd1 _13247_/B sky130_fd_sc_hd__and2b_1
X_10389_ _10390_/A _10390_/B vssd1 vssd1 vccd1 vccd1 _10391_/A sky130_fd_sc_hd__nand2_1
X_13177_ hold126/X _13191_/B vssd1 vssd1 vccd1 vccd1 hold127/A sky130_fd_sc_hd__or2_1
XANTENNA__10364__A2 _12667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12128_ _12129_/A _12164_/C vssd1 vssd1 vccd1 vccd1 _12128_/X sky130_fd_sc_hd__and2_1
X_12059_ hold275/A _12058_/X _09521_/Y vssd1 vssd1 vccd1 vccd1 _12059_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10116__A2 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08190__B1 _08580_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06985__B _07556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09270_ _10522_/B _09270_/B vssd1 vssd1 vccd1 vccd1 _09276_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_59_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08221_ _08243_/A _08243_/B _08189_/X vssd1 vssd1 vccd1 vccd1 _08229_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_118_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08152_ _08152_/A _08152_/B vssd1 vssd1 vccd1 vccd1 _08222_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_7_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10052__A1 _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07103_ _09524_/A _07087_/Y _07099_/X _09509_/A _07101_/X vssd1 vssd1 vccd1 vccd1
+ _07104_/B sky130_fd_sc_hd__o221a_2
XFILLER_0_15_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08796__A2 wire122/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08083_ _08873_/B2 fanout21/X _08246_/B _07406_/Y vssd1 vssd1 vccd1 vccd1 _08084_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10052__B2 _10374_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout115_A _07471_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07034_ _07007_/Y _07033_/X _10165_/A vssd1 vssd1 vccd1 vccd1 _07034_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_113_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08985_ _08572_/Y _09057_/B _08568_/Y vssd1 vssd1 vccd1 vccd1 _09065_/B sky130_fd_sc_hd__a21o_1
X_07936_ _07937_/A _07937_/B vssd1 vssd1 vccd1 vccd1 _09119_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11304__A1 _11527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11304__B2 _07526_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07867_ _07637_/B _07866_/X _07865_/X vssd1 vssd1 vccd1 vccd1 _11823_/A sky130_fd_sc_hd__o21a_4
XANTENNA__12389__S _12782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09606_ _09955_/A fanout9/X fanout4/X _09910_/A1 vssd1 vssd1 vccd1 vccd1 _09607_/B
+ sky130_fd_sc_hd__a22o_1
X_06818_ reg2_val[28] _06873_/B1 _06872_/B1 _06817_/Y vssd1 vssd1 vccd1 vccd1 _07062_/B
+ sky130_fd_sc_hd__o2bb2a_2
X_07798_ _07798_/A _07798_/B vssd1 vssd1 vccd1 vccd1 _08021_/A sky130_fd_sc_hd__xor2_1
X_09537_ _11576_/B _09537_/B vssd1 vssd1 vccd1 vccd1 _12783_/A sky130_fd_sc_hd__nand2_2
X_06749_ _09694_/A vssd1 vssd1 vccd1 vccd1 _12985_/A sky130_fd_sc_hd__inv_2
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09468_ reg1_val[9] reg1_val[22] _09493_/S vssd1 vssd1 vccd1 vccd1 _09468_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_109_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout28_A _07447_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07800__A _10239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08419_ _09671_/S fanout24/X _08486_/B _08873_/B2 vssd1 vssd1 vccd1 vccd1 _08420_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09399_ _10119_/A _09399_/B vssd1 vssd1 vccd1 vccd1 _09401_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11430_ _11430_/A _11430_/B vssd1 vssd1 vccd1 vccd1 _11431_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10043__B2 _10040_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11361_ reg1_val[12] curr_PC[12] _11244_/X vssd1 vssd1 vccd1 vccd1 _11362_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13100_ reg1_val[24] _13136_/A vssd1 vssd1 vccd1 vccd1 _13106_/A sky130_fd_sc_hd__nand2_1
X_10312_ _11472_/S _09851_/X _09534_/C vssd1 vssd1 vccd1 vccd1 _10313_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__11791__B2 _12047_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11292_ fanout46/X fanout20/X fanout18/X fanout50/X vssd1 vssd1 vccd1 vccd1 _11293_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08631__A _09948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08539__A2 _10049_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13031_ _13027_/A _13031_/B vssd1 vssd1 vccd1 vccd1 _13033_/C sky130_fd_sc_hd__nand2b_1
X_10243_ _10507_/A _10243_/B vssd1 vssd1 vccd1 vccd1 _10244_/A sky130_fd_sc_hd__xnor2_1
X_10174_ _11575_/S _10174_/B vssd1 vssd1 vccd1 vccd1 _10174_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_28_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout170 _12759_/A1 vssd1 vssd1 vccd1 vccd1 _09463_/S sky130_fd_sc_hd__clkbuf_8
Xfanout181 _10240_/A vssd1 vssd1 vccd1 vccd1 _09948_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_89_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout192 _09522_/Y vssd1 vssd1 vccd1 vccd1 _12796_/A1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10401__A _12253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08078__A _09591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09511__A_N _13748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12815_ _12816_/A _12816_/B _12816_/C vssd1 vssd1 vccd1 vccd1 _12823_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_97_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ hold299/A _12746_/B vssd1 vssd1 vccd1 vccd1 _12746_/X sky130_fd_sc_hd__or2_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12677_ _12677_/A _12677_/B _12677_/C vssd1 vssd1 vccd1 vccd1 _12680_/A sky130_fd_sc_hd__or3_1
XFILLER_0_37_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11628_ _11628_/A _11628_/B vssd1 vssd1 vccd1 vccd1 _11629_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_114_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11559_ _11761_/A _11559_/B vssd1 vssd1 vccd1 vccd1 _11561_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_123_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07986__B1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10585__A2 _10727_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09727__A1 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09727__B2 _07699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13229_ hold103/X hold255/X vssd1 vssd1 vccd1 vccd1 _13229_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_20_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07157__A _12982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08770_ _09373_/A _08770_/B vssd1 vssd1 vccd1 vccd1 _08774_/B sky130_fd_sc_hd__xnor2_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06961__A1 _06936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07721_ _07721_/A _07721_/B vssd1 vssd1 vccd1 vccd1 _07722_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_79_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08702__A2 _10538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07652_ _07652_/A _07652_/B vssd1 vssd1 vccd1 vccd1 _07653_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07583_ _07583_/A _07583_/B vssd1 vssd1 vccd1 vccd1 _07584_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_48_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09322_ _09094_/B _09094_/C _09825_/A _09205_/X _09986_/A vssd1 vssd1 vccd1 vccd1
+ _09325_/A sky130_fd_sc_hd__a2111o_1
XFILLER_0_63_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09253_ _10239_/A _09253_/B vssd1 vssd1 vccd1 vccd1 _09260_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__10457__S _10457_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08204_ _08201_/B _08201_/C _08201_/A vssd1 vssd1 vccd1 vccd1 _08205_/C sky130_fd_sc_hd__a21o_1
X_09184_ _09184_/A _09184_/B vssd1 vssd1 vccd1 vccd1 _09185_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10025__A1 _10734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08769__A2 _09216_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08135_ _08746_/A _08135_/B vssd1 vssd1 vccd1 vccd1 _08140_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10981__A _10981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11773__A1 _12515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08066_ _08951_/A _08066_/B vssd1 vssd1 vccd1 vccd1 _08133_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07017_ reg1_val[2] _09496_/S vssd1 vssd1 vccd1 vccd1 _07097_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09718__A1 _12537_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08941__A2 _09910_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08968_ _09016_/A _09016_/C _09016_/B vssd1 vssd1 vccd1 vccd1 _09019_/A sky130_fd_sc_hd__a21boi_2
XANTENNA__09282__A _10266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07919_ _10119_/A _07919_/B vssd1 vssd1 vccd1 vccd1 _07921_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08899_ _08970_/A _08970_/B vssd1 vssd1 vccd1 vccd1 _08971_/A sky130_fd_sc_hd__or2_1
X_10930_ _10931_/A _10931_/B vssd1 vssd1 vccd1 vccd1 _10932_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_98_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10861_ _11562_/A _10900_/A _10900_/B vssd1 vssd1 vccd1 vccd1 _10863_/A sky130_fd_sc_hd__o21ai_1
X_12600_ _07251_/A _12799_/A2 _12657_/B1 reg1_val[27] _12971_/S vssd1 vssd1 vccd1
+ vccd1 _12600_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_94_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _13580_/A _13580_/B vssd1 vssd1 vccd1 vccd1 _13580_/Y sky130_fd_sc_hd__nor2_1
X_10792_ _10791_/B _10791_/C _10537_/A vssd1 vssd1 vccd1 vccd1 _10793_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_109_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07530__A _11126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12531_ _12531_/A vssd1 vssd1 vccd1 vccd1 _12592_/B sky130_fd_sc_hd__inv_2
XFILLER_0_47_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08209__A1 _10049_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08209__B2 _09173_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12462_ _12782_/B _12462_/B vssd1 vssd1 vccd1 vccd1 _12462_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13202__A1 _12614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12005__A2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09957__A1 _10225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11413_ _11413_/A _11413_/B vssd1 vssd1 vccd1 vccd1 _11415_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09957__B2 _10104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12393_ hold229/A _13663_/Q _12393_/C vssd1 vssd1 vccd1 vccd1 _12467_/B sky130_fd_sc_hd__or3_1
XFILLER_0_105_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11344_ _11103_/X _11221_/X _11222_/X vssd1 vssd1 vccd1 vccd1 _11344_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09709__A1 _10007_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11275_ _11388_/A _11275_/B vssd1 vssd1 vccd1 vccd1 _11279_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13014_ reg1_val[7] _13015_/B vssd1 vssd1 vccd1 vccd1 _13014_/Y sky130_fd_sc_hd__nor2_1
X_10226_ wire122/X fanout16/X _07877_/X _07495_/X vssd1 vssd1 vccd1 vccd1 _10227_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07196__A1 _07594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08393__B1 _08486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10157_ _10045_/X _10200_/B _10730_/B vssd1 vssd1 vccd1 vccd1 _10157_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
X_10088_ fanout56/X fanout83/X fanout79/X fanout53/X vssd1 vssd1 vccd1 vccd1 _10089_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13441__A1 _11823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13161__B _13193_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12729_ _12628_/Y _12730_/C _12680_/A _12626_/A vssd1 vssd1 vccd1 vccd1 _12731_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap112 _07492_/Y vssd1 vssd1 vccd1 vccd1 _10374_/B2 sky130_fd_sc_hd__buf_6
XFILLER_0_20_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08271__A _08271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07423__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09940_ _09940_/A _09940_/B vssd1 vssd1 vccd1 vccd1 _09944_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12704__B1 _12748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09871_ _09871_/A _09871_/B _12235_/C vssd1 vssd1 vccd1 vccd1 _09871_/Y sky130_fd_sc_hd__nand3_2
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08384__B1 _08778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ _09373_/A _08822_/B vssd1 vssd1 vccd1 vccd1 _08828_/A sky130_fd_sc_hd__xnor2_2
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08753_ _08753_/A _08753_/B vssd1 vssd1 vccd1 vccd1 _08790_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08136__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout182_A _13444_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07704_ _07704_/A _07704_/B vssd1 vssd1 vccd1 vccd1 _07717_/B sky130_fd_sc_hd__xnor2_1
X_08684_ _08712_/A _08712_/B vssd1 vssd1 vccd1 vccd1 _08687_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12483__A2 _12667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07635_ _07462_/B _07377_/B _07376_/C _12647_/A vssd1 vssd1 vccd1 vccd1 _12656_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07566_ _07566_/A _07566_/B _07655_/A vssd1 vssd1 vccd1 vccd1 _07567_/B sky130_fd_sc_hd__and3_1
XFILLER_0_76_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08446__A _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09305_ _09193_/A _09193_/B _09191_/Y vssd1 vssd1 vccd1 vccd1 _09306_/B sky130_fd_sc_hd__a21boi_4
XFILLER_0_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07497_ _10266_/A _07497_/B vssd1 vssd1 vccd1 vccd1 _07499_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09236_ _10095_/A _09236_/B vssd1 vssd1 vccd1 vccd1 _09238_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_106_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07662__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09939__A1 _10814_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09167_ _09168_/A _09168_/B vssd1 vssd1 vccd1 vccd1 _09167_/X sky130_fd_sc_hd__and2_1
XANTENNA__09939__B2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11600__A _11600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08118_ _09381_/A _08118_/B vssd1 vssd1 vccd1 vccd1 _08224_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08181__A _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09098_ _09321_/A _12695_/B vssd1 vssd1 vccd1 vccd1 _12742_/B sky130_fd_sc_hd__nor2_1
X_08049_ _09575_/A _08049_/B vssd1 vssd1 vccd1 vccd1 _08054_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11060_ _11061_/A _11061_/B vssd1 vssd1 vccd1 vccd1 _11062_/A sky130_fd_sc_hd__nor2_1
X_10011_ _09858_/A _09855_/Y _09857_/B vssd1 vssd1 vccd1 vccd1 _10016_/A sky130_fd_sc_hd__o21a_1
XANTENNA__08127__B1 wire101/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11047__A _11047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11962_ _11961_/A _11961_/B _11961_/Y _12047_/C1 vssd1 vssd1 vccd1 vccd1 _11962_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12474__A2 _12754_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13701_ _13701_/CLK hold27/X vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__dfxtp_1
X_10913_ _11825_/A _10913_/B vssd1 vssd1 vccd1 vccd1 _10914_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11893_ curr_PC[18] _11893_/B vssd1 vssd1 vccd1 vccd1 _12070_/C sky130_fd_sc_hd__and2_1
XFILLER_0_79_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13632_ _13731_/CLK _13632_/D vssd1 vssd1 vccd1 vccd1 hold103/A sky130_fd_sc_hd__dfxtp_1
X_10844_ _10845_/B _10845_/A vssd1 vssd1 vccd1 vccd1 _10844_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10237__A1 _10536_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10237__B2 _10536_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13563_ hold278/X _13584_/B _13562_/X _13563_/B2 vssd1 vssd1 vccd1 vccd1 hold279/A
+ sky130_fd_sc_hd__a22o_1
X_10775_ _10776_/A _10776_/B vssd1 vssd1 vccd1 vccd1 _10777_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12514_ _12452_/A _12450_/X _06831_/B vssd1 vssd1 vccd1 vccd1 _12514_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13494_ _13494_/A _13494_/B vssd1 vssd1 vccd1 vccd1 _13494_/Y sky130_fd_sc_hd__xnor2_1
X_12445_ _11766_/B _12125_/X _12682_/B _12444_/X vssd1 vssd1 vccd1 vccd1 _12446_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07405__A2 _09703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12376_ _12480_/A _12376_/B vssd1 vssd1 vccd1 vccd1 _12376_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11327_ _11440_/A _11327_/B vssd1 vssd1 vccd1 vccd1 _11329_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_120_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11258_ _09521_/Y _11252_/Y _11253_/X _11257_/X vssd1 vssd1 vccd1 vccd1 _11258_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10209_ fanout39/X _11423_/A fanout74/X fanout36/X vssd1 vssd1 vccd1 vccd1 _10210_/B
+ sky130_fd_sc_hd__o22a_1
X_11189_ _11825_/A _11189_/B vssd1 vssd1 vccd1 vccd1 _11191_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12995__B _12995_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09650__A _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10476__A1 _12759_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07420_ _10457_/S _07420_/B vssd1 vssd1 vccd1 vccd1 _07420_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__09618__B1 _08246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08266__A _10236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07170__A _08203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07351_ _07351_/A _07351_/B vssd1 vssd1 vccd1 vccd1 _07351_/X sky130_fd_sc_hd__and2_1
XFILLER_0_128_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07282_ _07283_/A _07283_/B vssd1 vssd1 vccd1 vccd1 _07282_/X sky130_fd_sc_hd__and2_4
XFILLER_0_128_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09021_ _09021_/A _09021_/B vssd1 vssd1 vccd1 vccd1 _10864_/C sky130_fd_sc_hd__xor2_2
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11728__A1 _11922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11420__A _11802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11728__B2 wire101/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold201 hold201/A vssd1 vssd1 vccd1 vccd1 hold201/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 hold212/A vssd1 vssd1 vccd1 vccd1 hold212/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold223 hold223/A vssd1 vssd1 vccd1 vccd1 hold223/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10400__A1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold234 hold234/A vssd1 vssd1 vccd1 vccd1 hold234/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10400__B2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold245 hold245/A vssd1 vssd1 vccd1 vccd1 hold245/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold256 hold256/A vssd1 vssd1 vccd1 vccd1 hold256/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 hold267/A vssd1 vssd1 vccd1 vccd1 hold267/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 hold278/A vssd1 vssd1 vccd1 vccd1 hold278/X sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ _09923_/A _09923_/B vssd1 vssd1 vccd1 vccd1 _09964_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_0_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold289 hold289/A vssd1 vssd1 vccd1 vccd1 hold289/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13350__B1 _13450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09854_ _09696_/A _09696_/B _09695_/A vssd1 vssd1 vccd1 vccd1 _09858_/A sky130_fd_sc_hd__o21a_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12251__A _12417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11900__A1 _07230_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08805_ _08811_/B _08811_/A vssd1 vssd1 vccd1 vccd1 _08805_/Y sky130_fd_sc_hd__nand2b_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11900__B2 _12189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ _09785_/A _09785_/B vssd1 vssd1 vccd1 vccd1 _09786_/B sky130_fd_sc_hd__xor2_4
X_06997_ reg2_val[4] _07110_/A vssd1 vssd1 vccd1 vccd1 _06997_/X sky130_fd_sc_hd__and2_1
X_08736_ _08739_/A _08739_/B vssd1 vssd1 vccd1 vccd1 _08755_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10467__B2 _10465_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08667_ _08670_/A _08670_/B vssd1 vssd1 vccd1 vccd1 _08667_/Y sky130_fd_sc_hd__nand2_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13082__A _13082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07618_ _07672_/A _07619_/B vssd1 vssd1 vccd1 vccd1 _07618_/X sky130_fd_sc_hd__or2_1
XFILLER_0_95_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13405__A1 _11076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ _08806_/A2 _10225_/A _07556_/Y _08806_/B1 vssd1 vssd1 vccd1 vccd1 _08599_/B
+ sky130_fd_sc_hd__a22o_1
X_07549_ _07541_/X _07544_/Y _07545_/Y _11638_/A vssd1 vssd1 vccd1 vccd1 _07550_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10560_ _10412_/A _10412_/B _10413_/X vssd1 vssd1 vccd1 vccd1 _10565_/A sky130_fd_sc_hd__o21bai_1
XFILLER_0_63_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout10_A _09146_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09219_ _09219_/A _09219_/B vssd1 vssd1 vccd1 vccd1 _09220_/B sky130_fd_sc_hd__or2_1
XFILLER_0_51_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10491_ _11603_/A _10491_/B vssd1 vssd1 vccd1 vccd1 _10495_/A sky130_fd_sc_hd__xnor2_1
X_12230_ _12230_/A _12230_/B vssd1 vssd1 vccd1 vccd1 _12241_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_102_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12161_ curr_PC[21] _12160_/B _10342_/A vssd1 vssd1 vccd1 vccd1 _12161_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__12860__S _12867_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11112_ _11113_/B _11113_/C _11342_/A vssd1 vssd1 vccd1 vccd1 _11114_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12092_ _12092_/A _12092_/B vssd1 vssd1 vccd1 vccd1 _12094_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12144__A1 _12782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11043_ _11309_/A fanout9/X fanout4/X _07477_/X vssd1 vssd1 vccd1 vccd1 _11044_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12994_ reg1_val[3] _12995_/B vssd1 vssd1 vccd1 vccd1 _12994_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_98_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11945_ _11943_/Y _11945_/B vssd1 vssd1 vccd1 vccd1 _12035_/B sky130_fd_sc_hd__nand2b_4
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11505__A _11709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08086__A _10263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11876_ _11876_/A _11876_/B vssd1 vssd1 vccd1 vccd1 _11876_/X sky130_fd_sc_hd__xor2_1
XANTENNA__11670__A3 _12163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13615_ _13736_/CLK _13615_/D vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__dfxtp_1
X_10827_ _10827_/A _10827_/B vssd1 vssd1 vccd1 vccd1 _10828_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_67_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13546_ hold266/X _13555_/A2 _13545_/X _13563_/B2 vssd1 vssd1 vccd1 vccd1 hold267/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08823__A1 _08271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10758_ _10603_/S _10602_/X _09537_/B vssd1 vssd1 vccd1 vccd1 _10758_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_27_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08823__B2 _09501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13477_ _13591_/A hold288/X vssd1 vssd1 vccd1 vccd1 _13711_/D sky130_fd_sc_hd__and2_1
XFILLER_0_42_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10689_ _11913_/A _10689_/B vssd1 vssd1 vccd1 vccd1 _10690_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12428_ _12429_/B _12429_/A vssd1 vssd1 vccd1 vccd1 _12502_/B sky130_fd_sc_hd__and2b_1
XANTENNA__11186__A2 _07643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08051__A2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12359_ _12437_/B _12359_/B vssd1 vssd1 vccd1 vccd1 _12362_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_77_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13332__B1 _13506_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06920_ reg2_val[14] _06920_/B vssd1 vssd1 vccd1 vccd1 _06920_/X sky130_fd_sc_hd__and2_1
XANTENNA__12071__A _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06851_ instruction[33] _12981_/C vssd1 vssd1 vccd1 vccd1 _13020_/B sky130_fd_sc_hd__and2_4
X_09570_ _10078_/A _09570_/B vssd1 vssd1 vccd1 vccd1 _09579_/A sky130_fd_sc_hd__xnor2_1
X_06782_ instruction[1] instruction[2] instruction[0] pred_val vssd1 vssd1 vccd1 vccd1
+ _07110_/B sky130_fd_sc_hd__or4bb_1
X_08521_ _08521_/A _08521_/B vssd1 vssd1 vccd1 vccd1 _08560_/A sky130_fd_sc_hd__xnor2_1
X_08452_ _08501_/A _08501_/B _08439_/X vssd1 vssd1 vccd1 vccd1 _08460_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07403_ _10050_/A _07403_/B vssd1 vssd1 vccd1 vccd1 _07425_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08383_ _10944_/A _08383_/B vssd1 vssd1 vccd1 vccd1 _08389_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07331__C _07435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout145_A _09575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07334_ _07357_/A _07334_/B _07337_/B _07334_/D vssd1 vssd1 vccd1 vccd1 _07377_/B
+ sky130_fd_sc_hd__and4_2
XFILLER_0_45_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10621__A1 _12525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07265_ reg1_val[4] reg1_val[5] reg1_val[6] _07265_/D vssd1 vssd1 vccd1 vccd1 _07320_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_0_5_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09004_ _09004_/A _09004_/B vssd1 vssd1 vccd1 vccd1 _09005_/B sky130_fd_sc_hd__and2_1
XFILLER_0_116_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07196_ _07594_/B _07287_/A _07287_/B _07201_/B vssd1 vssd1 vccd1 vccd1 _07198_/B
+ sky130_fd_sc_hd__a211o_2
XANTENNA__08578__B1 _07545_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11177__A2 _10787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10385__B1 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09906_ _09907_/A _09907_/B vssd1 vssd1 vccd1 vccd1 _09908_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_67_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10688__A1 _12103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09837_ _10458_/S _09836_/X _09537_/B vssd1 vssd1 vccd1 vccd1 _09839_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__10688__B2 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11309__B _11802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08750__B1 _09173_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09768_ _11508_/A _09768_/B vssd1 vssd1 vccd1 vccd1 _09776_/A sky130_fd_sc_hd__xnor2_4
XANTENNA_fanout58_A _10522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08719_ _08719_/A _08719_/B vssd1 vssd1 vccd1 vccd1 _08727_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_68_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09699_ hold188/A _10606_/A2 _13642_/Q vssd1 vssd1 vccd1 vccd1 _09699_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _07198_/Y _07643_/B fanout12/X _11997_/A vssd1 vssd1 vccd1 vccd1 _11731_/B
+ sky130_fd_sc_hd__a22o_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12719__A1_N fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _11659_/Y _11661_/B vssd1 vssd1 vccd1 vccd1 _11856_/A sky130_fd_sc_hd__nand2b_2
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13400_ hold64/X _13416_/A2 _13420_/B1 hold19/X _13383_/A vssd1 vssd1 vccd1 vccd1
+ hold65/A sky130_fd_sc_hd__o221a_1
XFILLER_0_126_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10612_ hold301/A _12786_/B1 _10752_/B _12748_/B1 vssd1 vssd1 vccd1 vccd1 _10612_/X
+ sky130_fd_sc_hd__a31o_1
X_11592_ _11683_/B vssd1 vssd1 vccd1 vccd1 _11592_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_106_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13331_ _13359_/A hold223/X vssd1 vssd1 vccd1 vccd1 _13647_/D sky130_fd_sc_hd__and2_1
X_10543_ _10542_/B _10542_/C _10542_/A vssd1 vssd1 vccd1 vccd1 _10544_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_36_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13262_ hold253/X hold105/X vssd1 vssd1 vccd1 vccd1 _13493_/B sky130_fd_sc_hd__nand2b_1
X_10474_ _12648_/A _09529_/B _10473_/Y _10468_/X vssd1 vssd1 vccd1 vccd1 _10474_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_20_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11168__A2 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12213_ _12695_/A _12213_/B vssd1 vssd1 vccd1 vccd1 _12214_/B sky130_fd_sc_hd__nand2_1
X_13193_ hold118/X _13193_/B vssd1 vssd1 vccd1 vccd1 hold119/A sky130_fd_sc_hd__or2_1
XFILLER_0_32_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10376__B1 _07478_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12144_ _12782_/B _12142_/Y _12143_/Y _09529_/B vssd1 vssd1 vccd1 vccd1 _12144_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__09781__A2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12075_ _12413_/A fanout16/X fanout12/X _12331_/A vssd1 vssd1 vccd1 vccd1 _12076_/B
+ sky130_fd_sc_hd__a22o_1
X_11026_ _11027_/A _11027_/B vssd1 vssd1 vccd1 vccd1 _11209_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08809__A _10236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12977_ _12974_/B _12976_/B _12974_/A vssd1 vssd1 vccd1 vccd1 _12980_/A sky130_fd_sc_hd__o21ba_2
XFILLER_0_86_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11928_ _11807_/A _11807_/B _11805_/B vssd1 vssd1 vccd1 vccd1 _11931_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_47_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11859_ _11662_/X _12037_/A _11858_/A _11453_/X _11855_/X vssd1 vssd1 vccd1 vccd1
+ _11859_/Y sky130_fd_sc_hd__a221oi_1
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_18 instruction[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_29 reg1_val[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13529_ hold257/X _13555_/A2 _13528_/X _13542_/B2 vssd1 vssd1 vccd1 vccd1 hold258/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07050_ _07050_/A _07050_/B vssd1 vssd1 vccd1 vccd1 _07050_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_70_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10906__A2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07952_ _07952_/A _07952_/B vssd1 vssd1 vccd1 vccd1 _07954_/A sky130_fd_sc_hd__xnor2_4
X_06903_ instruction[26] _12981_/C vssd1 vssd1 vccd1 vccd1 _12806_/A sky130_fd_sc_hd__and2_2
X_07883_ _07874_/A _07874_/B _07884_/B vssd1 vssd1 vccd1 vccd1 _09113_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__08732__B1 _07420_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09622_ fanout28/X fanout76/X fanout74/X _08395_/B vssd1 vssd1 vccd1 vccd1 _09623_/B
+ sky130_fd_sc_hd__o22a_1
X_06834_ reg2_val[26] _06873_/B1 _06872_/B1 _06833_/Y vssd1 vssd1 vccd1 vccd1 _07217_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_78_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09553_ _12092_/A _09553_/B vssd1 vssd1 vccd1 vccd1 _09555_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06765_ pred_val instruction[1] vssd1 vssd1 vccd1 vccd1 _06775_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08504_ _08504_/A _08504_/B vssd1 vssd1 vccd1 vccd1 _08505_/B sky130_fd_sc_hd__nor2_1
X_09484_ _09482_/X _09483_/X _13145_/A vssd1 vssd1 vccd1 vccd1 _09484_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08435_ _10236_/A _08435_/B vssd1 vssd1 vccd1 vccd1 _08504_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10984__A _11225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08366_ _08293_/A _08292_/B _08292_/C vssd1 vssd1 vccd1 vccd1 _08367_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_46_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07317_ _07316_/A _07644_/B _07263_/Y _07656_/A _07656_/B vssd1 vssd1 vccd1 vccd1
+ _07506_/A sky130_fd_sc_hd__a32o_2
XFILLER_0_46_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_441 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08263__A2 _13166_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08297_ _08297_/A _08297_/B vssd1 vssd1 vccd1 vccd1 _08299_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07248_ _08951_/A _07248_/B vssd1 vssd1 vccd1 vccd1 _07264_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09212__A1 _07833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07179_ _10457_/S _09496_/S _10007_/S _13145_/A vssd1 vssd1 vccd1 vccd1 _07186_/B
+ sky130_fd_sc_hd__and4_4
XANTENNA__09212__B2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10190_ _07363_/B _11793_/B _10187_/Y _10188_/X _10189_/X vssd1 vssd1 vccd1 vccd1
+ _10190_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_112_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12900_ _12900_/A _12900_/B _12900_/C vssd1 vssd1 vccd1 vccd1 _12901_/B sky130_fd_sc_hd__nand3_1
XANTENNA__08629__A _10944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12831_ _12837_/B _12831_/B vssd1 vssd1 vccd1 vccd1 new_PC[4] sky130_fd_sc_hd__and2_4
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11055__A _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _09254_/A _12799_/A2 _12736_/Y _12761_/X _12971_/S vssd1 vssd1 vccd1 vccd1
+ dest_val[30] sky130_fd_sc_hd__o221a_4
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _11714_/A _11714_/B vssd1 vssd1 vccd1 vccd1 _11838_/B sky130_fd_sc_hd__nand2b_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _12693_/A _12693_/B vssd1 vssd1 vccd1 vccd1 _12693_/Y sky130_fd_sc_hd__nand2_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11644_ _11528_/A _11528_/B _11531_/A vssd1 vssd1 vccd1 vccd1 _11648_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11575_ _10598_/X _10600_/X _11575_/S vssd1 vssd1 vccd1 vccd1 _11575_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_24_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13314_ _13585_/A _13585_/B _13211_/A vssd1 vssd1 vccd1 vccd1 _13589_/B sky130_fd_sc_hd__o21ai_1
X_10526_ _07416_/X _11423_/A _07543_/X _07422_/Y vssd1 vssd1 vccd1 vccd1 _10527_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13245_ hold55/X hold292/A vssd1 vssd1 vccd1 vccd1 _13247_/A sky130_fd_sc_hd__and2b_1
X_10457_ _09713_/X _10456_/X _10457_/S vssd1 vssd1 vccd1 vccd1 _10457_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12614__A _12614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13176_ _11527_/A _13194_/A2 hold91/X _13543_/A vssd1 vssd1 vccd1 vccd1 _13624_/D
+ sky130_fd_sc_hd__o211a_1
X_10388_ _11913_/A _10388_/B vssd1 vssd1 vccd1 vccd1 _10390_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12127_ _12440_/A _12127_/B vssd1 vssd1 vccd1 vccd1 _12164_/C sky130_fd_sc_hd__xnor2_4
X_12058_ _12058_/A _12145_/B vssd1 vssd1 vccd1 vccd1 _12058_/X sky130_fd_sc_hd__and2_1
X_11009_ hold280/A _11252_/B _11251_/C _11008_/Y _12748_/B1 vssd1 vssd1 vccd1 vccd1
+ _11014_/B sky130_fd_sc_hd__a311o_1
XFILLER_0_79_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08190__A1 _09216_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08190__B2 _08868_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13066__A2 _13059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08220_ _08220_/A _08220_/B vssd1 vssd1 vccd1 vccd1 _08243_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_7_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08151_ _08225_/A _08225_/B _08143_/X vssd1 vssd1 vccd1 vccd1 _08222_/A sky130_fd_sc_hd__a21o_1
XANTENNA__11412__B _11413_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12041__A3 _12164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07102_ instruction[3] _13748_/A vssd1 vssd1 vccd1 vccd1 _09509_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10052__A2 _07643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08082_ _08088_/B _08088_/A vssd1 vssd1 vccd1 vccd1 _08082_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_30_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07033_ _07014_/Y _07032_/X _10026_/A vssd1 vssd1 vccd1 vccd1 _07033_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_113_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout108_A _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07205__B1 _08821_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08984_ _09049_/A _08980_/X _09049_/B _08657_/X _08981_/A vssd1 vssd1 vccd1 vccd1
+ _09057_/B sky130_fd_sc_hd__a32o_2
X_07935_ _09591_/A _07935_/B vssd1 vssd1 vccd1 vccd1 _07937_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08705__A0 _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10979__A _10981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07508__A1 _11126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11304__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07866_ reg1_val[29] _12656_/A vssd1 vssd1 vccd1 vccd1 _07866_/X sky130_fd_sc_hd__xor2_2
X_09605_ _09377_/A _09377_/B _09375_/Y vssd1 vssd1 vccd1 vccd1 _09609_/A sky130_fd_sc_hd__o21a_1
X_06817_ _06886_/A _13048_/B vssd1 vssd1 vccd1 vccd1 _06817_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_3_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07797_ _07993_/A _07993_/B _07793_/X vssd1 vssd1 vccd1 vccd1 _07798_/B sky130_fd_sc_hd__a21oi_2
X_09536_ _11576_/A _09536_/B vssd1 vssd1 vccd1 vccd1 _09537_/B sky130_fd_sc_hd__or2_4
X_06748_ _12982_/A vssd1 vssd1 vccd1 vccd1 _06748_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09467_ reg1_val[8] reg1_val[23] _09493_/S vssd1 vssd1 vccd1 vccd1 _09467_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_65_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08418_ _08418_/A _08418_/B vssd1 vssd1 vccd1 vccd1 _08427_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11603__A _11603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09398_ fanout39/X _07451_/X _10915_/A _08118_/B vssd1 vssd1 vccd1 vccd1 _09399_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08349_ _08349_/A _08349_/B _08349_/C vssd1 vssd1 vccd1 vccd1 _08353_/A sky130_fd_sc_hd__and3_1
XFILLER_0_34_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11360_ _11360_/A _11360_/B vssd1 vssd1 vccd1 vccd1 _11362_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10311_ _10311_/A _10311_/B vssd1 vssd1 vccd1 vccd1 _10311_/X sky130_fd_sc_hd__xor2_1
X_11291_ _11290_/B _11290_/C _11290_/A vssd1 vssd1 vccd1 vccd1 _11302_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13030_ _13030_/A _13039_/A vssd1 vssd1 vccd1 vccd1 _13033_/B sky130_fd_sc_hd__nand2_1
X_10242_ fanout45/X fanout75/X _08704_/B fanout49/X vssd1 vssd1 vccd1 vccd1 _10243_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10173_ _10600_/S _09458_/X _10172_/X vssd1 vssd1 vccd1 vccd1 _10174_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10751__B1 _12657_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10889__A _10889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout160 _13445_/A2 vssd1 vssd1 vccd1 vccd1 _13419_/A2 sky130_fd_sc_hd__buf_4
Xfanout171 _12759_/A1 vssd1 vssd1 vccd1 vccd1 _12710_/B2 sky130_fd_sc_hd__buf_4
Xfanout182 _13444_/B1 vssd1 vssd1 vccd1 vccd1 _13420_/B1 sky130_fd_sc_hd__buf_4
Xfanout193 _09519_/Y vssd1 vssd1 vccd1 vccd1 _11586_/B sky130_fd_sc_hd__buf_4
X_12814_ _12823_/A _12814_/B vssd1 vssd1 vccd1 vccd1 _12816_/C sky130_fd_sc_hd__nand2_1
XANTENNA__13453__C1 _13463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _09716_/Y _12744_/X _12782_/B vssd1 vssd1 vccd1 vccd1 _12745_/X sky130_fd_sc_hd__mux2_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _12724_/B _12676_/B vssd1 vssd1 vccd1 vccd1 _12677_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_127_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11627_ _11628_/A _11628_/B vssd1 vssd1 vccd1 vccd1 _11743_/A sky130_fd_sc_hd__and2_1
XFILLER_0_52_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11558_ _11113_/C _11556_/Y _11557_/X _11555_/Y vssd1 vssd1 vccd1 vccd1 _11559_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__08822__A _09373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07986__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11782__A2 _12793_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07986__B2 _08866_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10509_ _10510_/A _10510_/B vssd1 vssd1 vccd1 vccd1 _10511_/A sky130_fd_sc_hd__or2_1
XFILLER_0_100_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11489_ curr_PC[14] _11597_/C vssd1 vssd1 vccd1 vccd1 _11490_/B sky130_fd_sc_hd__and2_1
XFILLER_0_110_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09727__A2 _10522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13228_ _13226_/X _13228_/B vssd1 vssd1 vccd1 vccd1 _13557_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__13159__B _13193_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07157__B _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13159_ hold73/X _13193_/B vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__or2_1
XFILLER_0_0_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06961__A2 _06936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07720_ _07842_/A _07842_/B _07716_/X vssd1 vssd1 vccd1 vccd1 _07776_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__12495__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08269__A _09948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09360__B1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07173__A _10239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07651_ _07651_/A _07651_/B vssd1 vssd1 vccd1 vccd1 _07851_/A sky130_fd_sc_hd__xor2_4
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12247__B1 _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07582_ _11286_/A _07582_/B vssd1 vssd1 vccd1 vccd1 _07696_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13444__C1 _13444_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09321_ _09321_/A _12780_/A _12695_/B _12743_/A vssd1 vssd1 vccd1 vccd1 _09881_/A
+ sky130_fd_sc_hd__or4b_4
XANTENNA__12798__A1 _09507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11423__A _11423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09252_ _09582_/A fanout51/X fanout44/X _07200_/Y vssd1 vssd1 vccd1 vccd1 _09253_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_8_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08203_ _08203_/A _08203_/B vssd1 vssd1 vccd1 vccd1 _08205_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09183_ _09184_/A _09184_/B vssd1 vssd1 vccd1 vccd1 _09185_/A sky130_fd_sc_hd__and2_1
XFILLER_0_90_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout225_A _06906_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08134_ _09173_/B2 _10538_/A _08778_/B _11047_/A vssd1 vssd1 vccd1 vccd1 _08135_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10981__B _10981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08065_ _08866_/B2 fanout42/X fanout40/X _07240_/X vssd1 vssd1 vccd1 vccd1 _08066_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07016_ reg1_val[2] _10456_/S vssd1 vssd1 vccd1 vccd1 _07016_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_3_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08967_ _08929_/X _08967_/B vssd1 vssd1 vccd1 vccd1 _09013_/B sky130_fd_sc_hd__and2b_1
X_07918_ _08118_/B _07491_/X _07557_/Y fanout39/X vssd1 vssd1 vccd1 vccd1 _07919_/B
+ sky130_fd_sc_hd__o22a_1
X_08898_ _08898_/A _08898_/B vssd1 vssd1 vccd1 vccd1 _08970_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10502__A _11281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07849_ _07966_/B _07966_/A vssd1 vssd1 vccd1 vccd1 _07849_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_98_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07901__A1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07901__B2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10860_ _11106_/A _10860_/B vssd1 vssd1 vccd1 vccd1 _10900_/B sky130_fd_sc_hd__xnor2_4
XANTENNA_fanout40_A _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08907__A _08907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09519_ _09520_/A _09520_/B vssd1 vssd1 vccd1 vccd1 _09519_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_94_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10791_ _10537_/A _10791_/B _10791_/C vssd1 vssd1 vccd1 vccd1 _10791_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_94_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ hold207/A _12530_/B vssd1 vssd1 vccd1 vccd1 _12531_/A sky130_fd_sc_hd__nor2_1
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07665__B1 _08704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07530__B _07572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12461_ _12461_/A _12461_/B vssd1 vssd1 vccd1 vccd1 _12461_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__08209__A2 _10538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13202__A2 _13598_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11412_ _11413_/A _11413_/B vssd1 vssd1 vccd1 vccd1 _11530_/A sky130_fd_sc_hd__nor2_1
XANTENNA__09957__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12392_ hold269/A _12786_/B1 _12464_/B _12748_/B1 vssd1 vssd1 vccd1 vccd1 _12392_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11343_ _11343_/A _11556_/A vssd1 vssd1 vccd1 vccd1 _11343_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_105_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12164__A _12164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09709__A2 _11793_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11274_ _11274_/A _11274_/B vssd1 vssd1 vccd1 vccd1 _11275_/B sky130_fd_sc_hd__or2_1
XFILLER_0_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13013_ _13012_/A _13009_/Y _13011_/B vssd1 vssd1 vccd1 vccd1 _13017_/A sky130_fd_sc_hd__o21a_2
X_10225_ _10225_/A _10518_/A vssd1 vssd1 vccd1 vccd1 _10229_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08393__A1 _08873_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08393__B2 _13149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09590__B1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10156_ _10156_/A _10156_/B vssd1 vssd1 vccd1 vccd1 _10200_/B sky130_fd_sc_hd__nor2_1
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11508__A _11508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10087_ _11913_/A _10087_/B vssd1 vssd1 vccd1 vccd1 _10091_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__12229__B1 _12533_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10989_ _06963_/Y _10868_/X _06966_/B vssd1 vssd1 vccd1 vccd1 _10990_/B sky130_fd_sc_hd__o21a_1
XANTENNA__13441__A2 _13598_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12728_ _12728_/A _12765_/A vssd1 vssd1 vccd1 vccd1 _12730_/C sky130_fd_sc_hd__or2_1
XFILLER_0_84_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12659_ _06848_/D _12709_/A2 _10022_/Y _09504_/Y _12658_/Y vssd1 vssd1 vccd1 vccd1
+ _12659_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_127_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06771__S _07135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap102 _07300_/Y vssd1 vssd1 vccd1 vccd1 _13180_/A1 sky130_fd_sc_hd__buf_6
XFILLER_0_111_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08271__B wire101/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ hold285/A _09870_/B vssd1 vssd1 vccd1 vccd1 _09870_/Y sky130_fd_sc_hd__xnor2_2
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12802__A _12982_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08384__A1 _10522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _08821_/A1 _08866_/A2 _08923_/B1 _08821_/B2 vssd1 vssd1 vccd1 vccd1 _08822_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08384__B2 _09885_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ _08777_/A _08777_/B vssd1 vssd1 vccd1 vccd1 _08790_/A sky130_fd_sc_hd__nand2b_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08136__A1 _08873_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07703_ _12092_/A _07703_/B vssd1 vssd1 vccd1 vccd1 _07717_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08136__B2 _08891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08683_ _10236_/A _08683_/B vssd1 vssd1 vccd1 vccd1 _08712_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11140__B1 _11587_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07634_ reg1_val[28] _07634_/B _07634_/C _07634_/D vssd1 vssd1 vccd1 vccd1 _12656_/A
+ sky130_fd_sc_hd__or4_4
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07565_ _07566_/B _07655_/A _07566_/A vssd1 vssd1 vccd1 vccd1 _07948_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__12249__A _12420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13432__A2 _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09304_ _09304_/A _09304_/B vssd1 vssd1 vccd1 vccd1 _09306_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_91_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07496_ fanout21/X _07491_/X _08246_/B _09885_/B1 vssd1 vssd1 vccd1 vccd1 _07497_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_75_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09235_ fanout45/X _10235_/A1 _10235_/B2 fanout49/X vssd1 vssd1 vccd1 vccd1 _09236_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13196__A1 _12413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09166_ _09289_/A _09166_/B vssd1 vssd1 vccd1 vccd1 _09168_/B sky130_fd_sc_hd__or2_1
XANTENNA__09939__A2 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08117_ _08223_/A _08223_/B _08114_/Y vssd1 vssd1 vccd1 vccd1 _08152_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_9_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08072__B1 _08486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11600__B _11600_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09097_ _09097_/A _12583_/B _12584_/A _09096_/X vssd1 vssd1 vccd1 vccd1 _12695_/B
+ sky130_fd_sc_hd__or4bb_1
XFILLER_0_4_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08048_ _11047_/A fanout68/X fanout66/X fanout85/X vssd1 vssd1 vccd1 vccd1 _08049_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09572__B1 _10235_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout88_A _11507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10010_ _10003_/X _10009_/X _10458_/S vssd1 vssd1 vccd1 vccd1 _10010_/X sky130_fd_sc_hd__mux2_2
X_09999_ _09997_/X _09998_/X _10600_/S vssd1 vssd1 vccd1 vccd1 _09999_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08127__A1 _07239_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08127__B2 _07238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11961_ _11961_/A _11961_/B vssd1 vssd1 vccd1 vccd1 _11961_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11047__B _11825_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10912_ _07477_/X fanout9/X fanout4/X _07472_/Y vssd1 vssd1 vccd1 vccd1 _10913_/B
+ sky130_fd_sc_hd__a22o_1
X_13700_ _13700_/CLK _13700_/D vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13543__A _13543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11892_ curr_PC[18] _11893_/B vssd1 vssd1 vccd1 vccd1 _11894_/B sky130_fd_sc_hd__nor2_1
X_13631_ _13731_/CLK hold50/X vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10890__C1 _12327_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10843_ _10843_/A _10843_/B vssd1 vssd1 vccd1 vccd1 _10845_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13423__A2 _13445_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10237__A2 _12614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13562_ hold269/X _13561_/X fanout2/X vssd1 vssd1 vccd1 vccd1 _13562_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10774_ _11913_/A _10774_/B vssd1 vssd1 vccd1 vccd1 _10776_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12513_ _12513_/A _12635_/B vssd1 vssd1 vccd1 vccd1 _12513_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13493_ _13261_/X _13493_/B vssd1 vssd1 vccd1 vccd1 _13494_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_109_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12444_ _12124_/Y _12682_/B _12443_/Y vssd1 vssd1 vccd1 vccd1 _12444_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12375_ _12480_/A _12376_/B vssd1 vssd1 vccd1 vccd1 _12375_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_105_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10945__B1 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11326_ _11326_/A _11326_/B _11326_/C _11326_/D vssd1 vssd1 vccd1 vccd1 _11327_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_22_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11257_ _07321_/X _07533_/X _12235_/C _11256_/X vssd1 vssd1 vccd1 vccd1 _11257_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_0_66_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10208_ _11719_/A _10208_/B vssd1 vssd1 vccd1 vccd1 _10212_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11188_ _07526_/Y fanout9/X fanout4/X _11309_/A vssd1 vssd1 vccd1 vccd1 _11189_/B
+ sky130_fd_sc_hd__a22o_1
X_10139_ _09975_/A _09975_/B _09973_/X vssd1 vssd1 vccd1 vccd1 _10140_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__07435__B _07435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09931__A _10542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09650__B _09650_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07451__A _10889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10881__C1 _09529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09618__A1 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09618__B2 _07522_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07350_ _07483_/A _07377_/A _07337_/B _07348_/A vssd1 vssd1 vccd1 vccd1 _07351_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_57_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07281_ _07281_/A _07310_/B _07281_/C vssd1 vssd1 vccd1 vccd1 _07283_/B sky130_fd_sc_hd__or3_4
XFILLER_0_31_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09020_ _10731_/B _10731_/C vssd1 vssd1 vccd1 vccd1 _10864_/B sky130_fd_sc_hd__and2_1
XANTENNA__13178__A1 _11638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11728__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold202 hold202/A vssd1 vssd1 vccd1 vccd1 hold202/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10936__B1 _11027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold213 hold213/A vssd1 vssd1 vccd1 vccd1 hold213/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12235__C _12235_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold224 hold224/A vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07801__B1 _11638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10400__A2 _07543_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold235 hold297/A vssd1 vssd1 vccd1 vccd1 hold235/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold246 hold246/A vssd1 vssd1 vccd1 vccd1 hold246/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold257 hold257/A vssd1 vssd1 vccd1 vccd1 hold257/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 hold299/X vssd1 vssd1 vccd1 vccd1 hold268/X sky130_fd_sc_hd__buf_1
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09922_ _09922_/A _09922_/B vssd1 vssd1 vccd1 vccd1 _09923_/B sky130_fd_sc_hd__nor2_1
Xhold279 hold279/A vssd1 vssd1 vccd1 vccd1 hold279/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12689__B1 _10730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07626__A _10119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09853_ _09846_/X _09852_/X _10458_/S vssd1 vssd1 vccd1 vccd1 _09853_/X sky130_fd_sc_hd__mux2_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08804_ _08804_/A _08804_/B vssd1 vssd1 vccd1 vccd1 _08811_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07345__B _07594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09784_ _09785_/A _09785_/B vssd1 vssd1 vccd1 vccd1 _09784_/Y sky130_fd_sc_hd__nor2_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06996_ _06996_/A _06996_/B vssd1 vssd1 vccd1 vccd1 _10311_/A sky130_fd_sc_hd__nor2_1
X_08735_ _09373_/A _08735_/B vssd1 vssd1 vccd1 vccd1 _08739_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__13363__A _13543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ _09659_/B _08666_/B vssd1 vssd1 vccd1 vccd1 _08670_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10467__A2 _11793_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07361__A _12253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07617_ _07617_/A _07617_/B vssd1 vssd1 vccd1 vccd1 _07619_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__13082__B _13082_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08597_ _08600_/A _08600_/B vssd1 vssd1 vccd1 vccd1 _08597_/Y sky130_fd_sc_hd__nand2_1
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13405__A2 _13445_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07548_ _06911_/B _07296_/Y _07297_/Y _07189_/Y vssd1 vssd1 vccd1 vccd1 _07548_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_119_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07479_ fanout24/X _11047_/A _08486_/B fanout85/X vssd1 vssd1 vccd1 vccd1 _07480_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_64_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09218_ _09219_/A _09219_/B vssd1 vssd1 vccd1 vccd1 _09220_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_106_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10490_ _07299_/Y fanout36/X fanout70/X fanout38/X vssd1 vssd1 vccd1 vccd1 _10491_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_32_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09149_ _09150_/A _09150_/B vssd1 vssd1 vccd1 vccd1 _09149_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10227__A _11823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09793__B1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12160_ curr_PC[21] _12160_/B vssd1 vssd1 vccd1 vccd1 _12325_/C sky130_fd_sc_hd__and2_2
X_11111_ _11111_/A vssd1 vssd1 vccd1 vccd1 _11113_/C sky130_fd_sc_hd__inv_2
X_12091_ fanout15/X _12614_/A _12667_/A fanout31/X vssd1 vssd1 vccd1 vccd1 _12092_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11042_ _11161_/B _11042_/B vssd1 vssd1 vccd1 vccd1 _11066_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_99_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12993_ _12992_/A _12989_/Y _12991_/B vssd1 vssd1 vccd1 vccd1 _12997_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_99_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07859__B1 _07522_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11944_ _11944_/A _11944_/B _11944_/C vssd1 vssd1 vccd1 vccd1 _11945_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_86_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11875_ _11779_/A _11776_/Y _11778_/B vssd1 vssd1 vccd1 vccd1 _11876_/B sky130_fd_sc_hd__o21ai_1
X_10826_ _10828_/B vssd1 vssd1 vccd1 vccd1 _10964_/A sky130_fd_sc_hd__inv_2
X_13614_ _13719_/CLK hold80/X vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__dfxtp_1
X_10757_ _09523_/Y _10747_/Y _10748_/X _10756_/Y vssd1 vssd1 vccd1 vccd1 _10757_/X
+ sky130_fd_sc_hd__a31o_1
X_13545_ hold275/A _13544_/X fanout1/X vssd1 vssd1 vccd1 vccd1 _13545_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08823__A2 _07492_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13476_ hold287/X _13550_/A2 _13475_/X _13563_/B2 vssd1 vssd1 vccd1 vccd1 hold288/A
+ sky130_fd_sc_hd__a22o_1
X_10688_ _12103_/A fanout29/X fanout27/X fanout54/X vssd1 vssd1 vccd1 vccd1 _10689_/B
+ sky130_fd_sc_hd__o22a_1
X_12427_ _12502_/A _12427_/B vssd1 vssd1 vccd1 vccd1 _12429_/B sky130_fd_sc_hd__or2_1
XFILLER_0_22_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10918__B1 _08246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12358_ _12358_/A _12358_/B _12358_/C vssd1 vssd1 vccd1 vccd1 _12359_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_77_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11309_ _11309_/A _11802_/B vssd1 vssd1 vccd1 vccd1 _11310_/B sky130_fd_sc_hd__nand2_1
X_12289_ _12440_/A _12440_/B vssd1 vssd1 vccd1 vccd1 _12290_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07446__A _11913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13167__B _13191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07165__B _07572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06850_ _06850_/A _06850_/B vssd1 vssd1 vccd1 vccd1 _07099_/A sky130_fd_sc_hd__or2_1
X_06781_ instruction[1] instruction[2] instruction[0] pred_val vssd1 vssd1 vccd1 vccd1
+ _06781_/X sky130_fd_sc_hd__and4bb_2
XFILLER_0_26_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08520_ _08520_/A _08520_/B vssd1 vssd1 vccd1 vccd1 _08573_/A sky130_fd_sc_hd__xnor2_2
X_08451_ _08451_/A _08451_/B vssd1 vssd1 vccd1 vccd1 _08501_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07402_ _09381_/A fanout35/X _08873_/B2 _07699_/B vssd1 vssd1 vccd1 vccd1 _07403_/B
+ sky130_fd_sc_hd__o22a_1
X_08382_ _08923_/B1 fanout84/X _08580_/B _08866_/A2 vssd1 vssd1 vccd1 vccd1 _08383_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07333_ reg1_val[20] reg1_val[21] vssd1 vssd1 vccd1 vccd1 _07339_/D sky130_fd_sc_hd__or2_1
XANTENNA__08275__B1 _11638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout138_A _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07264_ _07264_/A _07264_/B vssd1 vssd1 vccd1 vccd1 _07316_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10621__A2 _12760_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09003_ _09003_/A _09003_/B vssd1 vssd1 vccd1 vccd1 _09082_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07195_ _07201_/A _07213_/A _07521_/A _06875_/B vssd1 vssd1 vccd1 vccd1 _07198_/A
+ sky130_fd_sc_hd__a211o_2
XANTENNA__08578__A1 _07399_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08578__B2 _09910_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11177__A3 _10787_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10385__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10385__B2 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09527__B1 _09523_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09905_ _10119_/A _09905_/B vssd1 vssd1 vccd1 vccd1 _09907_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09836_ _11575_/S _09835_/X _09534_/C vssd1 vssd1 vccd1 vccd1 _09836_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10688__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11885__B2 _10889_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08750__A1 _08907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08750__B2 _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ fanout42/X fanout83/X fanout79/X fanout40/X vssd1 vssd1 vccd1 vccd1 _09768_/B
+ sky130_fd_sc_hd__o22a_2
X_06979_ _06977_/Y _06979_/B vssd1 vssd1 vccd1 vccd1 _10592_/A sky130_fd_sc_hd__and2b_1
X_08718_ _08730_/A _08730_/B vssd1 vssd1 vccd1 vccd1 _08719_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09698_ _12525_/A _09692_/X _09697_/Y _12760_/A1 vssd1 vssd1 vccd1 vccd1 _09698_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08649_ _08646_/A _08646_/B _08698_/A vssd1 vssd1 vccd1 vccd1 _08660_/A sky130_fd_sc_hd__a21bo_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ _11660_/A _11660_/B _11660_/C vssd1 vssd1 vccd1 vccd1 _11661_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_49_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ _12786_/B1 _10752_/B hold301/A vssd1 vssd1 vccd1 vccd1 _10611_/Y sky130_fd_sc_hd__a21oi_1
X_11591_ _10458_/S _09497_/X _09537_/B vssd1 vssd1 vccd1 vccd1 _11683_/B sky130_fd_sc_hd__o21a_1
X_13330_ hold182/X _13506_/B2 _13506_/A2 hold222/X vssd1 vssd1 vccd1 vccd1 hold223/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10542_ _10542_/A _10542_/B _10542_/C vssd1 vssd1 vccd1 vccd1 _10544_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_51_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13261_ hold105/X hold253/X vssd1 vssd1 vccd1 vccd1 _13261_/X sky130_fd_sc_hd__and2b_1
X_10473_ _10473_/A _10473_/B vssd1 vssd1 vccd1 vccd1 _10473_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12212_ _12695_/A _12165_/Y _12372_/C _11955_/A vssd1 vssd1 vccd1 vccd1 _12212_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_121_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13192_ _07230_/Y _13194_/A2 hold104/X _13591_/A vssd1 vssd1 vccd1 vccd1 _13632_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_121_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10376__A1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10376__B2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12143_ _12782_/B _12143_/B vssd1 vssd1 vccd1 vccd1 _12143_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09518__B1 _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07266__A _13015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12074_ _12025_/A _12025_/B _12023_/Y vssd1 vssd1 vccd1 vccd1 _12117_/A sky130_fd_sc_hd__a21o_1
X_11025_ _10927_/A _10926_/B _10924_/X vssd1 vssd1 vccd1 vccd1 _11027_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12976_ _12976_/A _12976_/B vssd1 vssd1 vccd1 vccd1 new_PC[26] sky130_fd_sc_hd__xnor2_4
XFILLER_0_87_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11927_ _11830_/A _11830_/B _11828_/Y vssd1 vssd1 vccd1 vccd1 _11933_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11858_ _11858_/A vssd1 vssd1 vccd1 vccd1 _11858_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13450__B _13450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10809_ _10809_/A _10809_/B vssd1 vssd1 vccd1 vccd1 _10828_/A sky130_fd_sc_hd__nand2_1
XANTENNA_19 instruction[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11789_ _09521_/Y _11786_/X _11788_/Y _09523_/Y vssd1 vssd1 vccd1 vccd1 _11789_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13528_ hold292/A _13527_/X fanout1/X vssd1 vssd1 vccd1 vccd1 _13528_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_27_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13459_ _13459_/A hold286/X vssd1 vssd1 vccd1 vccd1 _13707_/D sky130_fd_sc_hd__and2_1
XFILLER_0_112_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10367__B2 _10236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07951_ _07951_/A _07951_/B vssd1 vssd1 vccd1 vccd1 _07952_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__06991__B1 _12782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06902_ _06902_/A _06902_/B vssd1 vssd1 vccd1 vccd1 _11774_/A sky130_fd_sc_hd__and2_2
XFILLER_0_128_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07882_ _07882_/A _07882_/B vssd1 vssd1 vccd1 vccd1 _07884_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08732__A1 _08806_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07904__A _09575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08732__B2 _08806_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09621_ _10119_/A _09621_/B vssd1 vssd1 vccd1 vccd1 _09625_/A sky130_fd_sc_hd__xnor2_1
X_06833_ _06928_/B _13036_/B vssd1 vssd1 vccd1 vccd1 _06833_/Y sky130_fd_sc_hd__nor2_1
X_09552_ _07833_/B wire122/X _10637_/A fanout14/X vssd1 vssd1 vccd1 vccd1 _09553_/B
+ sky130_fd_sc_hd__a22o_1
X_06764_ rst vssd1 vssd1 vccd1 vccd1 _06764_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08503_ _08503_/A _08503_/B vssd1 vssd1 vccd1 vccd1 _08507_/A sky130_fd_sc_hd__xnor2_1
X_09483_ _09694_/A _13129_/A _09839_/A vssd1 vssd1 vccd1 vccd1 _09483_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08434_ _08873_/A2 _09173_/B2 _11047_/A _08891_/B vssd1 vssd1 vccd1 vccd1 _08435_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_53_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08735__A _09373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10984__B _10984_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08365_ _08298_/X _08365_/B vssd1 vssd1 vccd1 vccd1 _09081_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_92_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07316_ _07316_/A _07316_/B vssd1 vssd1 vccd1 vccd1 _07656_/B sky130_fd_sc_hd__xnor2_1
X_08296_ _08360_/A _08360_/B _08241_/Y vssd1 vssd1 vccd1 vccd1 _08299_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07247_ fanout49/X _08950_/B fanout45/X _08866_/B2 vssd1 vssd1 vccd1 vccd1 _07248_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07178_ _07544_/A _07527_/A vssd1 vssd1 vccd1 vccd1 _07188_/C sky130_fd_sc_hd__or2_1
XANTENNA__09212__A2 _10374_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11555__B1 _11553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10505__A _11709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout70_A _07548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09819_ _09819_/A _09819_/B vssd1 vssd1 vccd1 vccd1 _09821_/B sky130_fd_sc_hd__xnor2_4
X_12830_ _12830_/A _12830_/B _12830_/C vssd1 vssd1 vccd1 vccd1 _12831_/B sky130_fd_sc_hd__nand3_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08487__A0 _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _12781_/A _12743_/Y _12760_/X _12741_/X vssd1 vssd1 vccd1 vccd1 _12761_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _11712_/A _11712_/B vssd1 vssd1 vccd1 vccd1 _11714_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_68_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _07083_/Y _12691_/Y _12738_/S vssd1 vssd1 vccd1 vccd1 _12693_/B sky130_fd_sc_hd__mux2_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _11525_/A _11525_/B _11532_/Y vssd1 vssd1 vccd1 vccd1 _11652_/A sky130_fd_sc_hd__a21bo_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09987__B1 _09824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11574_ _11574_/A _11574_/B vssd1 vssd1 vccd1 vccd1 _11574_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10525_ _12551_/A _10525_/B vssd1 vssd1 vccd1 vccd1 _10533_/A sky130_fd_sc_hd__xnor2_1
X_13313_ _13313_/A _13580_/A vssd1 vssd1 vccd1 vccd1 _13585_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13244_ _13244_/A _13244_/B vssd1 vssd1 vccd1 vccd1 _13531_/A sky130_fd_sc_hd__nor2_1
X_10456_ _09847_/X _09850_/X _10456_/S vssd1 vssd1 vccd1 vccd1 _10456_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10349__A1 _10349_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12614__B _12764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13175_ hold90/X _13191_/B vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__or2_1
X_10387_ _07282_/X fanout29/X fanout27/X fanout40/X vssd1 vssd1 vccd1 vccd1 _10388_/B
+ sky130_fd_sc_hd__o22a_1
X_12126_ _11766_/B _12125_/X _12124_/Y vssd1 vssd1 vccd1 vccd1 _12127_/B sky130_fd_sc_hd__a21oi_2
X_12057_ hold298/A _12057_/B vssd1 vssd1 vccd1 vccd1 _12145_/B sky130_fd_sc_hd__or2_1
XANTENNA__07724__A _09575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11008_ _11252_/B _11251_/C hold280/A vssd1 vssd1 vccd1 vccd1 _11008_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__08190__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11246__A _12525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08478__B1 _13168_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12274__A1 _12189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12959_ reg1_val[24] curr_PC[24] _12978_/S vssd1 vssd1 vccd1 vccd1 _12960_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_90_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11482__C1 _11481_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08150_ _08150_/A _08150_/B vssd1 vssd1 vccd1 vccd1 _08225_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07101_ instruction[3] _13748_/A _07101_/C vssd1 vssd1 vccd1 vccd1 _07101_/X sky130_fd_sc_hd__or3_1
X_08081_ _08079_/Y _08115_/B _08076_/X vssd1 vssd1 vccd1 vccd1 _08088_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_3_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09993__A3 _10726_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12805__A _12806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09386__A _09386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07032_ _07022_/Y _09703_/C _07097_/B vssd1 vssd1 vccd1 vccd1 _07032_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_30_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07205__A1 _08821_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07205__B2 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08983_ _08983_/A _09052_/A vssd1 vssd1 vccd1 vccd1 _09049_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10044__B _10726_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10760__A1 _12760_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07934_ fanout83/X fanout76/X fanout74/X fanout79/X vssd1 vssd1 vccd1 vccd1 _07935_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10979__B _11106_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09902__B1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07865_ reg1_val[29] _07865_/B vssd1 vssd1 vccd1 vccd1 _07865_/X sky130_fd_sc_hd__or2_1
XFILLER_0_98_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09604_ _09604_/A _10518_/A vssd1 vssd1 vccd1 vccd1 _09610_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11156__A _11281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06816_ instruction[38] _12981_/C vssd1 vssd1 vccd1 vccd1 _13048_/B sky130_fd_sc_hd__and2_4
X_07796_ _07796_/A _07796_/B vssd1 vssd1 vccd1 vccd1 _07993_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_64_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09535_ _11576_/A _09536_/B vssd1 vssd1 vccd1 vccd1 _09535_/Y sky130_fd_sc_hd__nor2_2
X_06747_ instruction[41] vssd1 vssd1 vccd1 vccd1 _06747_/Y sky130_fd_sc_hd__inv_2
X_09466_ _09458_/X _09465_/X _10176_/A vssd1 vssd1 vccd1 vccd1 _09466_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_66_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08417_ _08417_/A _08417_/B vssd1 vssd1 vccd1 vccd1 _08460_/A sky130_fd_sc_hd__xor2_4
X_09397_ _10263_/A _09397_/B vssd1 vssd1 vccd1 vccd1 _09401_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08348_ _08260_/A _08260_/C _08260_/B vssd1 vssd1 vccd1 vccd1 _08349_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08279_ _10266_/A _08279_/B vssd1 vssd1 vccd1 vccd1 _08350_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10310_ _10734_/A _07000_/Y _07034_/X _10309_/Y vssd1 vssd1 vccd1 vccd1 _10311_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_116_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11290_ _11290_/A _11290_/B _11290_/C vssd1 vssd1 vccd1 vccd1 _11302_/A sky130_fd_sc_hd__or3_1
X_10241_ _10241_/A _10241_/B vssd1 vssd1 vccd1 vccd1 _10255_/A sky130_fd_sc_hd__xnor2_1
X_10172_ _10176_/A _10172_/B vssd1 vssd1 vccd1 vccd1 _10172_/X sky130_fd_sc_hd__or2_1
Xfanout150 _09748_/A vssd1 vssd1 vccd1 vccd1 _09910_/A1 sky130_fd_sc_hd__buf_6
XANTENNA__10889__B _10889_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout161 _13598_/C vssd1 vssd1 vccd1 vccd1 _13445_/A2 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07544__A _07544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13150__C1 _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout172 _09434_/Y vssd1 vssd1 vccd1 vccd1 _12759_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout183 _07117_/Y vssd1 vssd1 vccd1 vccd1 _13444_/B1 sky130_fd_sc_hd__buf_4
Xfanout194 _09516_/X vssd1 vssd1 vccd1 vccd1 _11587_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12813_ _12990_/B _12813_/B vssd1 vssd1 vccd1 vccd1 _12814_/B sky130_fd_sc_hd__or2_1
XANTENNA__10267__B1 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _13129_/A _12782_/C vssd1 vssd1 vccd1 vccd1 _12744_/X sky130_fd_sc_hd__xor2_1
XANTENNA__08375__A _09659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _12675_/A _12675_/B _12675_/C vssd1 vssd1 vccd1 vccd1 _12676_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11626_ _12092_/A _11626_/B vssd1 vssd1 vccd1 vccd1 _11628_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11767__B1 _10730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08632__B1 _13172_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11557_ _10578_/X _10579_/X _10581_/Y _11107_/Y _11556_/Y vssd1 vssd1 vccd1 vccd1
+ _11557_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_123_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10508_ _10508_/A _10508_/B vssd1 vssd1 vccd1 vccd1 _10510_/B sky130_fd_sc_hd__xnor2_1
X_11488_ curr_PC[14] _11597_/C vssd1 vssd1 vccd1 vccd1 _11488_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10439_ _10434_/X _10435_/X _10438_/Y _10981_/A vssd1 vssd1 vccd1 vccd1 _10441_/A
+ sky130_fd_sc_hd__a31o_1
X_13227_ hold282/A hold118/X vssd1 vssd1 vccd1 vccd1 _13228_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_122_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13158_ _07556_/Y _13196_/A2 hold36/X _13547_/A vssd1 vssd1 vccd1 vccd1 _13615_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _12110_/A _12110_/B _12110_/C vssd1 vssd1 vccd1 vccd1 _12111_/A sky130_fd_sc_hd__o21ai_1
X_13089_ reg1_val[20] _13129_/B _13085_/A vssd1 vssd1 vccd1 vccd1 _13090_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__06769__S _07135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06961__A3 _13029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12495__A1 _12614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13175__B _13191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12495__B2 _07257_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09360__A1 _11732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09360__B2 _10814_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07650_ _07648_/Y _07650_/B vssd1 vssd1 vccd1 vccd1 _07651_/B sky130_fd_sc_hd__and2b_1
X_07581_ _13174_/A1 _07541_/X _07544_/Y _07545_/Y vssd1 vssd1 vccd1 vccd1 _07582_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13444__B1 _13444_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09320_ _09986_/A _10579_/A vssd1 vssd1 vccd1 vccd1 _12780_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_47_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09251_ _09371_/A _09251_/B vssd1 vssd1 vccd1 vccd1 _09261_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__11423__B _11825_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08202_ _07237_/Y _11732_/A _10814_/A1 _07240_/X vssd1 vssd1 vccd1 vccd1 _08203_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09182_ _09182_/A _09182_/B vssd1 vssd1 vccd1 vccd1 _09184_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08133_ _08133_/A _08133_/B vssd1 vssd1 vccd1 vccd1 _08150_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout120_A _07456_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10981__C _10981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08064_ _08064_/A _08064_/B vssd1 vssd1 vccd1 vccd1 _08133_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_114_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07015_ reg1_val[2] _10456_/S vssd1 vssd1 vccd1 vccd1 _07015_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10055__A _12092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08966_ _08967_/B _09013_/A _08929_/X vssd1 vssd1 vccd1 vccd1 _09016_/C sky130_fd_sc_hd__a21o_1
X_07917_ _10050_/A _07917_/B vssd1 vssd1 vccd1 vccd1 _07921_/A sky130_fd_sc_hd__xnor2_1
X_08897_ _08897_/A _08897_/B vssd1 vssd1 vccd1 vccd1 _08970_/A sky130_fd_sc_hd__or2_1
XANTENNA__12486__B2 _12417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07848_ _07848_/A _07848_/B vssd1 vssd1 vccd1 vccd1 _07966_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09512__D_N _13744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07779_ _07653_/A _07653_/B _07659_/B _07657_/Y vssd1 vssd1 vccd1 vccd1 _07782_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09518_ _12598_/C _09517_/X _08197_/A vssd1 vssd1 vccd1 vccd1 _09528_/B sky130_fd_sc_hd__a21o_1
X_10790_ _11286_/A _10790_/B _10790_/C vssd1 vssd1 vccd1 vccd1 _10791_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_78_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07665__A1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _09445_/X _09448_/X _10005_/S vssd1 vssd1 vccd1 vccd1 _09449_/X sky130_fd_sc_hd__mux2_1
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07665__B2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12460_ _12458_/Y _12460_/B vssd1 vssd1 vccd1 vccd1 _12461_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11411_ _07518_/Y fanout7/X _11410_/X _11281_/A vssd1 vssd1 vccd1 vccd1 _11413_/B
+ sky130_fd_sc_hd__a22o_2
XANTENNA__07417__A1 _12421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12391_ _12314_/A _12464_/B hold269/A vssd1 vssd1 vccd1 vccd1 _12391_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11342_ _11342_/A _11452_/A vssd1 vssd1 vccd1 vccd1 _11556_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12164__B _12164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11273_ _11274_/A _11274_/B vssd1 vssd1 vccd1 vccd1 _11388_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_120_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13012_ _13012_/A _13012_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[6] sky130_fd_sc_hd__xnor2_4
X_10224_ _10224_/A _10224_/B vssd1 vssd1 vccd1 vccd1 _10259_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08393__A2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09590__A1 _10814_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09590__B2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10155_ _10155_/A _10155_/B _10155_/C vssd1 vssd1 vccd1 vccd1 _10156_/B sky130_fd_sc_hd__and3_1
XFILLER_0_100_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07274__A _09948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10086_ _11732_/A fanout29/X fanout27/X _07310_/Y vssd1 vssd1 vccd1 vccd1 _10087_/B
+ sky130_fd_sc_hd__o22a_1
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10488__B1 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13426__B1 _13444_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10988_ _10988_/A _10988_/B vssd1 vssd1 vccd1 vccd1 _10988_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12727_ _12727_/A _12727_/B vssd1 vssd1 vccd1 vccd1 _12765_/B sky130_fd_sc_hd__or2_1
XFILLER_0_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12658_ _06821_/Y _09520_/X _12657_/X vssd1 vssd1 vccd1 vccd1 _12658_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__08833__A _09381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11609_ _11610_/A _11610_/B _11610_/C vssd1 vssd1 vccd1 vccd1 _11611_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12589_ _12589_/A _12589_/B vssd1 vssd1 vccd1 vccd1 _12589_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xmax_cap114 _07472_/Y vssd1 vssd1 vccd1 vccd1 _13168_/A1 sky130_fd_sc_hd__buf_6
XFILLER_0_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08384__A2 _10538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _08820_/A _08820_/B vssd1 vssd1 vccd1 vccd1 _08836_/A sky130_fd_sc_hd__xnor2_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12090__A _12253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10191__A2 _11587_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ _09950_/A _08751_/B vssd1 vssd1 vccd1 vccd1 _08777_/B sky130_fd_sc_hd__xnor2_2
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08136__A2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07702_ _09604_/A fanout14/X _07833_/B _09748_/A vssd1 vssd1 vccd1 vccd1 _07703_/B
+ sky130_fd_sc_hd__a22o_1
X_08682_ _08873_/A2 _09216_/B2 _08868_/B1 _08891_/B vssd1 vssd1 vccd1 vccd1 _08683_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07344__B1 _07363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07633_ _07633_/A _07633_/B vssd1 vssd1 vccd1 vccd1 _07647_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_88_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07564_ _07654_/A _07654_/B vssd1 vssd1 vccd1 vccd1 _07655_/A sky130_fd_sc_hd__or2_1
XFILLER_0_76_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09303_ _09303_/A _09303_/B vssd1 vssd1 vccd1 vccd1 _09304_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_75_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07495_ _07184_/D _07448_/Y _07449_/Y _07193_/A vssd1 vssd1 vccd1 vccd1 _07495_/X
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_76_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09234_ _09575_/A _09234_/B vssd1 vssd1 vccd1 vccd1 _09238_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09839__A _09839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09165_ _09288_/A _09165_/B vssd1 vssd1 vccd1 vccd1 _09166_/B sky130_fd_sc_hd__and2_1
XANTENNA__13196__A2 _13196_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12265__A _12764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08116_ _08116_/A _08116_/B vssd1 vssd1 vccd1 vccd1 _08223_/B sky130_fd_sc_hd__xor2_1
XANTENNA__08072__A1 _09216_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09096_ _09094_/B _09094_/C _09094_/A vssd1 vssd1 vccd1 vccd1 _09096_/X sky130_fd_sc_hd__a21o_1
XANTENNA__08072__B2 _08868_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08047_ _10095_/A _08047_/B vssd1 vssd1 vccd1 vccd1 _08054_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09572__A1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09572__B2 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ _09666_/X _09674_/X _10004_/S vssd1 vssd1 vccd1 vccd1 _09998_/X sky130_fd_sc_hd__mux2_1
X_08949_ _09659_/B _08949_/B vssd1 vssd1 vccd1 vccd1 _08954_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08127__A2 _11922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07575__A_N _11076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11960_ _12515_/S _11959_/X _11958_/X vssd1 vssd1 vccd1 vccd1 _11961_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_98_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07822__A _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10911_ _10794_/A _10793_/B _10791_/X vssd1 vssd1 vccd1 vccd1 _10914_/A sky130_fd_sc_hd__a21o_1
X_11891_ _11862_/Y _11863_/X _11864_/X _11866_/Y _11890_/X vssd1 vssd1 vccd1 vccd1
+ _11891_/X sky130_fd_sc_hd__o221a_1
X_13630_ _13731_/CLK hold87/X vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__dfxtp_1
X_10842_ _10711_/A _10711_/B _10709_/Y vssd1 vssd1 vccd1 vccd1 _10843_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13561_ _13561_/A _13561_/B vssd1 vssd1 vccd1 vccd1 _13561_/X sky130_fd_sc_hd__xor2_1
X_10773_ fanout54/X fanout29/X fanout27/X _12268_/A vssd1 vssd1 vccd1 vccd1 _10774_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_82_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12512_ _12513_/A _12635_/B vssd1 vssd1 vccd1 vccd1 _12512_/X sky130_fd_sc_hd__and2_1
X_13492_ _13543_/A hold254/X vssd1 vssd1 vccd1 vccd1 _13714_/D sky130_fd_sc_hd__and2_1
XFILLER_0_35_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12443_ _12441_/Y _12443_/B vssd1 vssd1 vccd1 vccd1 _12443_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_62_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12395__B1 _12795_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12374_ _12374_/A _12733_/A vssd1 vssd1 vccd1 vccd1 _12376_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10945__B2 _07546_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11325_ _11326_/A _11326_/B _11326_/C _11326_/D vssd1 vssd1 vccd1 vccd1 _11440_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_50_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12903__A _13059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12147__B1 _12748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11256_ _11237_/A _12793_/A2 _11586_/B _06943_/A _11255_/Y vssd1 vssd1 vccd1 vccd1
+ _11256_/X sky130_fd_sc_hd__a221o_1
X_10207_ fanout34/X _10915_/A _07471_/Y fanout32/X vssd1 vssd1 vccd1 vccd1 _10208_/B
+ sky130_fd_sc_hd__o22a_1
X_11187_ _11731_/A _11187_/B vssd1 vssd1 vccd1 vccd1 _11191_/A sky130_fd_sc_hd__xnor2_1
X_10138_ _10138_/A _10138_/B vssd1 vssd1 vccd1 vccd1 _10140_/A sky130_fd_sc_hd__xnor2_2
X_10069_ _10070_/A _10070_/B vssd1 vssd1 vccd1 vccd1 _10217_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_82_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09618__A2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08826__B1 _08868_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07280_ _07310_/B _07281_/C _07281_/A vssd1 vssd1 vccd1 vccd1 _07283_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_73_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13178__A2 _13194_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07179__A _10457_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold203 hold203/A vssd1 vssd1 vccd1 vccd1 hold203/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 hold214/A vssd1 vssd1 vccd1 vccd1 hold214/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07801__A1 _08806_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold225 hold225/A vssd1 vssd1 vccd1 vccd1 hold225/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07801__B2 _08806_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12813__A _12990_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold236 hold236/A vssd1 vssd1 vccd1 vccd1 hold236/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold247 hold247/A vssd1 vssd1 vccd1 vccd1 hold247/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold258 hold258/A vssd1 vssd1 vccd1 vccd1 hold258/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09394__A _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09921_ _09922_/A _09922_/B vssd1 vssd1 vccd1 vccd1 _10060_/B sky130_fd_sc_hd__nand2_1
Xhold269 hold269/A vssd1 vssd1 vccd1 vccd1 hold269/X sky130_fd_sc_hd__buf_1
XFILLER_0_111_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06811__A _09254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13350__A2 _13463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09852_ _09849_/X _09851_/X _11575_/S vssd1 vssd1 vccd1 vccd1 _09852_/X sky130_fd_sc_hd__mux2_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08803_ _08820_/A _08802_/Y _08798_/Y vssd1 vssd1 vccd1 vccd1 _08811_/A sky130_fd_sc_hd__o21ai_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _09783_/A _09783_/B vssd1 vssd1 vccd1 vccd1 _09785_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__07345__C _10603_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06995_ reg1_val[5] _06995_/B vssd1 vssd1 vccd1 vccd1 _06996_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_56_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08734_ _08821_/A1 _10522_/A _08868_/B1 _08821_/B2 vssd1 vssd1 vccd1 vccd1 _08735_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08738__A _10542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ _12982_/A _07478_/A _07478_/B _08271_/A _13168_/A1 vssd1 vssd1 vccd1 vccd1
+ _08666_/B sky130_fd_sc_hd__a32o_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ _07616_/A _07616_/B vssd1 vssd1 vccd1 vccd1 _07617_/B sky130_fd_sc_hd__xnor2_2
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08596_ _10236_/A _08596_/B vssd1 vssd1 vccd1 vccd1 _08600_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07547_ _07189_/Y _07297_/Y _07296_/Y _06911_/B vssd1 vssd1 vccd1 vccd1 _07547_/X
+ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__10624__B1 _12867_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07478_ _07478_/A _07478_/B vssd1 vssd1 vccd1 vccd1 _07478_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_64_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09217_ _10050_/A _09217_/B vssd1 vssd1 vccd1 vccd1 _09219_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09288__B _10522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07089__A _09501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09148_ _09949_/A _09148_/B vssd1 vssd1 vccd1 vccd1 _09150_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__09242__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09793__A1 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09079_ _09079_/A _09079_/B vssd1 vssd1 vccd1 vccd1 _09080_/C sky130_fd_sc_hd__or2_1
XANTENNA__09793__B2 _08395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11110_ _10854_/Y _11343_/A _11109_/Y vssd1 vssd1 vccd1 vccd1 _11111_/A sky130_fd_sc_hd__a21o_1
X_12090_ _12253_/A _12090_/B vssd1 vssd1 vccd1 vccd1 _12096_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11041_ _11041_/A _11041_/B vssd1 vssd1 vccd1 vccd1 _11042_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10243__A _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12992_ _12992_/A _12992_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[2] sky130_fd_sc_hd__xor2_4
XFILLER_0_99_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07859__A1 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11943_ _11944_/A _11944_/B _11944_/C vssd1 vssd1 vccd1 vccd1 _11943_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__07859__B2 _08486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11074__A _11281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07271__B _07572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11874_ _11874_/A _11874_/B vssd1 vssd1 vccd1 vccd1 _11876_/A sky130_fd_sc_hd__nand2_1
X_13613_ _13717_/CLK _13613_/D vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08808__B1 _08923_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10825_ _10827_/A _10827_/B vssd1 vssd1 vccd1 vccd1 _10828_/B sky130_fd_sc_hd__and2_1
XANTENNA__12065__C1 _12064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12604__A1 _09529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11802__A wire101/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13544_ _13544_/A _13544_/B vssd1 vssd1 vccd1 vccd1 _13544_/X sky130_fd_sc_hd__xor2_1
XANTENNA__08383__A _10944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10756_ _06971_/Y _10749_/Y _10751_/X _10755_/X vssd1 vssd1 vccd1 vccd1 _10756_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12617__B fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13475_ hold294/A _13474_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13475_/X sky130_fd_sc_hd__mux2_1
X_10687_ _10523_/A _10523_/B _10521_/A vssd1 vssd1 vccd1 vccd1 _10702_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_70_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12426_ _12426_/A _12426_/B _12426_/C vssd1 vssd1 vccd1 vccd1 _12427_/B sky130_fd_sc_hd__and3_1
XANTENNA__09233__B1 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10918__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10918__B2 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12357_ _12358_/A _12358_/B _12358_/C vssd1 vssd1 vccd1 vccd1 _12437_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_10_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11308_ _11308_/A _11308_/B vssd1 vssd1 vccd1 vccd1 _11310_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_10_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12288_ _12288_/A _12288_/B vssd1 vssd1 vccd1 vccd1 _12442_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_120_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13332__A2 _13506_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11239_ _10174_/B _10178_/A _11575_/S vssd1 vssd1 vccd1 vccd1 _11240_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09942__A _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06780_ instruction[0] instruction[1] instruction[2] instruction[41] pred_val vssd1
+ vssd1 vccd1 vccd1 _13082_/A sky130_fd_sc_hd__o311a_4
XANTENNA__13183__B _13191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08450_ _08506_/A _08506_/B _08449_/A vssd1 vssd1 vccd1 vccd1 _08501_/A sky130_fd_sc_hd__o21ai_2
X_07401_ _12485_/A _07401_/B vssd1 vssd1 vccd1 vccd1 _07401_/Y sky130_fd_sc_hd__nand2_1
X_08381_ _08453_/A _08453_/B _08378_/Y vssd1 vssd1 vccd1 vccd1 _08397_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_58_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10606__B1 _12533_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07332_ reg1_val[20] reg1_val[21] vssd1 vssd1 vccd1 vccd1 _07334_/D sky130_fd_sc_hd__nor2_1
XANTENNA__08275__A1 _07239_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08275__B2 _07238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06806__A _09254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07263_ _07264_/A _07264_/B vssd1 vssd1 vccd1 vccd1 _07263_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_116_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09002_ _09318_/A _09002_/B vssd1 vssd1 vccd1 vccd1 _09321_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07194_ _07201_/A _07521_/A vssd1 vssd1 vccd1 vccd1 _07287_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_5_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08578__A2 _07541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11031__B1 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout200_A _08203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10385__A2 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09904_ fanout38/X _07478_/Y _07522_/Y fanout36/X vssd1 vssd1 vccd1 vccd1 _09905_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_1_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07538__B1 _11076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09835_ _10600_/S _09686_/X _10601_/C vssd1 vssd1 vccd1 vccd1 _09835_/X sky130_fd_sc_hd__o21a_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08750__A2 _10049_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09766_ _09766_/A _09766_/B vssd1 vssd1 vccd1 vccd1 _09786_/A sky130_fd_sc_hd__nand2_1
X_06978_ _13015_/A _07492_/A vssd1 vssd1 vccd1 vccd1 _06979_/B sky130_fd_sc_hd__nand2_1
X_08717_ _08717_/A _08717_/B vssd1 vssd1 vccd1 vccd1 _08730_/B sky130_fd_sc_hd__xnor2_2
X_09697_ _12525_/A _09697_/B vssd1 vssd1 vccd1 vccd1 _09697_/Y sky130_fd_sc_hd__nand2_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09998__S _10004_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08648_ _08697_/A _08697_/B vssd1 vssd1 vccd1 vccd1 _08698_/A sky130_fd_sc_hd__or2_1
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12047__C1 _12047_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08579_ _11286_/A _08579_/B vssd1 vssd1 vccd1 vccd1 _08582_/B sky130_fd_sc_hd__xnor2_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12718__A fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ hold287/A _10610_/B vssd1 vssd1 vccd1 vccd1 _10752_/B sky130_fd_sc_hd__or2_1
XFILLER_0_119_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12062__A2 _09520_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11590_ _12748_/B1 _11580_/X _11581_/Y _11589_/X vssd1 vssd1 vccd1 vccd1 _11590_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10541_ _09575_/A _10541_/B _10541_/C vssd1 vssd1 vccd1 vccd1 _10542_/C sky130_fd_sc_hd__nand3b_1
XFILLER_0_106_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13260_ hold280/X hold62/X vssd1 vssd1 vccd1 vccd1 _13498_/B sky130_fd_sc_hd__nand2b_1
X_10472_ _10470_/Y _10472_/B vssd1 vssd1 vccd1 vccd1 _10473_/B sky130_fd_sc_hd__nand2b_1
X_12211_ _12695_/A _12165_/Y _12372_/C vssd1 vssd1 vccd1 vccd1 _12211_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13191_ hold103/X _13191_/B vssd1 vssd1 vccd1 vccd1 hold104/A sky130_fd_sc_hd__or2_1
XFILLER_0_121_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10376__A2 _11047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12142_ _12142_/A _12142_/B vssd1 vssd1 vccd1 vccd1 _12142_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__09518__A1 _12598_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12073_ _11988_/A _12164_/A _12164_/B _11231_/A vssd1 vssd1 vccd1 vccd1 _12129_/A
+ sky130_fd_sc_hd__o31a_1
X_11024_ _10968_/A _10968_/B _10969_/Y vssd1 vssd1 vccd1 vccd1 _11101_/A sky130_fd_sc_hd__a21bo_1
X_12975_ _12968_/B _12970_/B _12968_/A vssd1 vssd1 vccd1 vccd1 _12976_/B sky130_fd_sc_hd__o21ba_2
Xclkbuf_4_2_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13649_/CLK sky130_fd_sc_hd__clkbuf_8
X_11926_ _11821_/A _11821_/B _11833_/A vssd1 vssd1 vccd1 vccd1 _11938_/A sky130_fd_sc_hd__o21a_1
X_11857_ _11857_/A _12037_/A vssd1 vssd1 vccd1 vccd1 _11858_/A sky130_fd_sc_hd__and2_1
X_10808_ _10808_/A _10808_/B vssd1 vssd1 vccd1 vccd1 _10809_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_55_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11788_ hold200/A _11788_/B vssd1 vssd1 vccd1 vccd1 _11788_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13527_ _13527_/A _13527_/B vssd1 vssd1 vccd1 vccd1 _13527_/X sky130_fd_sc_hd__xor2_1
X_10739_ reg1_val[8] curr_PC[8] vssd1 vssd1 vccd1 vccd1 _10739_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09937__A _11281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13458_ hold285/X _13450_/B _13457_/X _13463_/B2 vssd1 vssd1 vccd1 vccd1 hold286/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13459__A _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12409_ _12666_/A _12409_/B vssd1 vssd1 vccd1 vccd1 _12411_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13389_ _09371_/A _13419_/A2 hold102/X vssd1 vssd1 vccd1 vccd1 _13676_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_88_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10367__A2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07950_ _07948_/A _07948_/B _07951_/B vssd1 vssd1 vccd1 vccd1 _07950_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__07176__B _07398_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06901_ reg1_val[17] _07300_/A vssd1 vssd1 vccd1 vccd1 _06902_/B sky130_fd_sc_hd__nand2_1
X_07881_ _07882_/A _07882_/B vssd1 vssd1 vccd1 vccd1 _09113_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_128_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08732__A2 _09910_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09620_ fanout39/X _10915_/A _07471_/Y _08118_/B vssd1 vssd1 vccd1 vccd1 _09621_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11707__A _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06832_ instruction[36] _12981_/C vssd1 vssd1 vccd1 vccd1 _13036_/B sky130_fd_sc_hd__and2_4
XFILLER_0_128_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09551_ _11731_/A _09551_/B vssd1 vssd1 vccd1 vccd1 _09555_/A sky130_fd_sc_hd__xnor2_1
X_06763_ curr_PC[3] vssd1 vssd1 vccd1 vccd1 _10041_/A sky130_fd_sc_hd__inv_2
X_08502_ _08510_/B _08510_/A vssd1 vssd1 vccd1 vccd1 _08512_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_78_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09482_ _09501_/A reg1_val[31] _09839_/A vssd1 vssd1 vccd1 vccd1 _09482_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08433_ _08436_/A _08436_/B vssd1 vssd1 vccd1 vccd1 _08438_/A sky130_fd_sc_hd__and2_1
XFILLER_0_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout150_A _09748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout248_A _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08364_ _08364_/A _08364_/B vssd1 vssd1 vccd1 vccd1 _09077_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07131__S _07135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07315_ _07721_/A _07721_/B vssd1 vssd1 vccd1 vccd1 _07656_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_18_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08295_ _08302_/A _08302_/B _08284_/X vssd1 vssd1 vccd1 vccd1 _08360_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_18_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07246_ _07687_/A _07687_/B _07227_/Y vssd1 vssd1 vccd1 vccd1 _07316_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08751__A _09950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07177_ _11463_/A _07398_/B vssd1 vssd1 vccd1 vccd1 _07177_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12752__B1 _12795_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08184__B1 _08395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09818_ _09819_/B _09819_/A vssd1 vssd1 vccd1 vccd1 _09818_/Y sky130_fd_sc_hd__nand2b_1
X_09749_ _10104_/A fanout9/X fanout4/X _09955_/A vssd1 vssd1 vccd1 vccd1 _09750_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10818__B1 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _12760_/A1 _12745_/X _12753_/Y _12759_/X vssd1 vssd1 vccd1 vccd1 _12760_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _11712_/A _11712_/B vssd1 vssd1 vccd1 vccd1 _11838_/A sky130_fd_sc_hd__or2_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _06821_/Y _12640_/X _06824_/B vssd1 vssd1 vccd1 vccd1 _12691_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09436__A0 _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _11642_/A _11642_/B vssd1 vssd1 vccd1 vccd1 _11654_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09987__A1 _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09987__B2 _09824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11573_ _11471_/A _11471_/B _11469_/B vssd1 vssd1 vccd1 vccd1 _11574_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_107_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13312_ _13579_/B _13579_/C _13579_/A vssd1 vssd1 vccd1 vccd1 _13580_/A sky130_fd_sc_hd__o21a_1
X_10524_ fanout34/X _07478_/Y _07522_/Y fanout32/X vssd1 vssd1 vccd1 vccd1 _10525_/B
+ sky130_fd_sc_hd__o22a_1
X_13243_ hold257/X hold37/X vssd1 vssd1 vccd1 vccd1 _13244_/B sky130_fd_sc_hd__and2b_1
X_10455_ _10453_/X _10454_/X _11575_/S vssd1 vssd1 vccd1 vccd1 _10455_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10349__A2 _10518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13174_ _13174_/A1 _13194_/A2 hold67/X _13543_/A vssd1 vssd1 vccd1 vccd1 _13623_/D
+ sky130_fd_sc_hd__o211a_1
X_10386_ _11709_/A _10386_/B vssd1 vssd1 vccd1 vccd1 _10390_/A sky130_fd_sc_hd__xnor2_1
X_12125_ _12035_/B _12125_/B _12207_/A vssd1 vssd1 vccd1 vccd1 _12125_/X sky130_fd_sc_hd__and3b_1
X_12056_ _12056_/A _12056_/B hold212/A vssd1 vssd1 vccd1 vccd1 _12056_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ hold253/A _11007_/B vssd1 vssd1 vccd1 vccd1 _11251_/C sky130_fd_sc_hd__or2_1
XANTENNA__11527__A _11527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08478__A1 _08933_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12958_ _12961_/D _12958_/B vssd1 vssd1 vccd1 vccd1 new_PC[23] sky130_fd_sc_hd__xnor2_4
XANTENNA__12274__A2 _12764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08478__B2 _07175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07740__A _10542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11482__B1 _09523_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11909_ _12093_/A _11909_/B vssd1 vssd1 vccd1 vccd1 _11915_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12889_ _13048_/B _12890_/B vssd1 vssd1 vccd1 vccd1 _12900_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_23_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07100_ _07099_/X _12778_/A _13744_/A vssd1 vssd1 vccd1 vccd1 _07101_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_15_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08080_ _08080_/A _08080_/B vssd1 vssd1 vccd1 vccd1 _08115_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07031_ _07026_/A _07026_/B _09703_/B _08197_/A vssd1 vssd1 vccd1 vccd1 _09703_/C
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12093__A _12093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06803__B _12981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07205__A2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08982_ _08982_/A _08982_/B _08982_/C vssd1 vssd1 vccd1 vccd1 _09052_/A sky130_fd_sc_hd__and3_1
XFILLER_0_48_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07933_ _11286_/A _07933_/B vssd1 vssd1 vccd1 vccd1 _07937_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09902__A1 _11732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09902__B2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07864_ _07864_/A _07864_/B vssd1 vssd1 vccd1 vccd1 _07870_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07913__B1 _07833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09603_ _09726_/A _09602_/C _09602_/A vssd1 vssd1 vccd1 vccd1 _09611_/B sky130_fd_sc_hd__a21o_1
X_06815_ _06815_/A _06815_/B vssd1 vssd1 vccd1 vccd1 _12693_/A sky130_fd_sc_hd__nor2_2
X_07795_ _10507_/A _07795_/B vssd1 vssd1 vccd1 vccd1 _07993_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09534_ _10601_/B _10601_/C _09534_/C vssd1 vssd1 vccd1 vccd1 _11576_/B sky130_fd_sc_hd__and3_1
X_06746_ instruction[5] vssd1 vssd1 vccd1 vccd1 _09516_/A sky130_fd_sc_hd__inv_2
XANTENNA__08746__A _08746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09465_ _09461_/X _09464_/X _10005_/S vssd1 vssd1 vccd1 vccd1 _09465_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12268__A _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08416_ _08416_/A _08416_/B vssd1 vssd1 vccd1 vccd1 _08463_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09396_ fanout28/X _07522_/Y fanout76/X fanout27/X vssd1 vssd1 vccd1 vccd1 _09397_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_65_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08347_ _08347_/A _08347_/B vssd1 vssd1 vccd1 vccd1 _08349_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_19_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08278_ _08350_/A _08278_/B _08278_/C vssd1 vssd1 vccd1 vccd1 _08350_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_34_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07229_ _07230_/A _07230_/B vssd1 vssd1 vccd1 vccd1 _07229_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_104_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10240_ _10240_/A _10240_/B vssd1 vssd1 vccd1 vccd1 _10241_/B sky130_fd_sc_hd__xnor2_1
X_10171_ _09449_/X _09465_/X _10600_/S vssd1 vssd1 vccd1 vccd1 _10171_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10751__A2 _11793_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout140 _12311_/B1 vssd1 vssd1 vccd1 vccd1 _10606_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout151 _07406_/Y vssd1 vssd1 vccd1 vccd1 _13149_/A sky130_fd_sc_hd__buf_8
Xfanout162 _13196_/A2 vssd1 vssd1 vccd1 vccd1 _13598_/C sky130_fd_sc_hd__buf_4
XANTENNA__11347__A _11554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout184 _13450_/B vssd1 vssd1 vccd1 vccd1 _13506_/A2 sky130_fd_sc_hd__buf_4
Xfanout195 _09508_/Y vssd1 vssd1 vccd1 vccd1 _12793_/A2 sky130_fd_sc_hd__clkbuf_8
X_12812_ _12990_/B _12813_/B vssd1 vssd1 vccd1 vccd1 _12823_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10267__A1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12743_ _12743_/A _12743_/B vssd1 vssd1 vccd1 vccd1 _12743_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10267__B2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ _12675_/A _12675_/B _12675_/C vssd1 vssd1 vccd1 vccd1 _12724_/B sky130_fd_sc_hd__o21a_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10019__A1 _10456_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11625_ _07230_/Y fanout15/X fanout31/X _12331_/A vssd1 vssd1 vccd1 vccd1 _11626_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08632__A1 _08271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11556_ _11556_/A _11763_/A vssd1 vssd1 vccd1 vccd1 _11556_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__08632__B2 _09501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10507_ _10507_/A _10507_/B vssd1 vssd1 vccd1 vccd1 _10508_/B sky130_fd_sc_hd__xnor2_1
X_11487_ _11458_/X _11459_/Y _11461_/Y _11866_/A _11486_/X vssd1 vssd1 vccd1 vccd1
+ _11487_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_123_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13226_ hold118/X hold282/A vssd1 vssd1 vccd1 vccd1 _13226_/X sky130_fd_sc_hd__and2b_1
X_10438_ _10438_/A _10438_/B vssd1 vssd1 vccd1 vccd1 _10438_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_100_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08396__A0 _10263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13157_ hold35/X _13191_/B vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__or2_1
XFILLER_0_20_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10369_ _10369_/A _10369_/B vssd1 vssd1 vccd1 vccd1 _10370_/B sky130_fd_sc_hd__and2_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ _12192_/B _12108_/B vssd1 vssd1 vccd1 vccd1 _12110_/C sky130_fd_sc_hd__nor2_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ _13086_/Y _13088_/B vssd1 vssd1 vccd1 vccd1 _13102_/B sky130_fd_sc_hd__nand2b_2
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12039_ _12207_/A _12368_/A vssd1 vssd1 vccd1 vccd1 _12164_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__12495__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09950__A _09950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09360__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07580_ _07583_/A _07583_/B vssd1 vssd1 vccd1 vccd1 _07584_/A sky130_fd_sc_hd__and2_1
XANTENNA__12247__A2 _12372_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13191__B _13191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12652__C1 _12795_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09250_ _07238_/X _12614_/A _12667_/A _07239_/Y vssd1 vssd1 vccd1 vccd1 _09251_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10301__B1_N _10300_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08201_ _08201_/A _08201_/B _08201_/C vssd1 vssd1 vccd1 vccd1 _08205_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_56_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09181_ _09182_/B _09182_/A vssd1 vssd1 vccd1 vccd1 _09301_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_28_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08132_ _08152_/A _08152_/B vssd1 vssd1 vccd1 vccd1 _08132_/X sky130_fd_sc_hd__and2b_1
XANTENNA__09397__A _10263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10981__D _11106_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08063_ _08064_/A _08064_/B vssd1 vssd1 vccd1 vccd1 _08063_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_fanout113_A _07491_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12707__B1 _12795_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07014_ reg1_val[2] _10176_/A vssd1 vssd1 vccd1 vccd1 _07014_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_12_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08387__B1 _07545_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13380__B1 _13584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12551__A _12551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08965_ _08937_/X _09012_/A _08964_/B vssd1 vssd1 vccd1 vccd1 _09013_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__11167__A _12417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07916_ fanout35/X _13149_/A _08923_/B1 _07699_/B vssd1 vssd1 vccd1 vccd1 _07917_/B
+ sky130_fd_sc_hd__o22a_1
X_08896_ _08897_/A _08896_/B _08896_/C _08896_/D vssd1 vssd1 vccd1 vccd1 _08897_/B
+ sky130_fd_sc_hd__nor4_1
XANTENNA__12486__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07847_ _07844_/A _07844_/B _08037_/A vssd1 vssd1 vccd1 vccd1 _07966_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_79_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07778_ _07709_/A _07709_/B _07708_/A vssd1 vssd1 vccd1 vccd1 _07783_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_79_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09517_ _10866_/B _11587_/A2 _13145_/A vssd1 vssd1 vccd1 vccd1 _09517_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12643__C1 _09507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ _09446_/X _09447_/X _09674_/S vssd1 vssd1 vccd1 vccd1 _09448_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_93_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07665__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout26_A fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09379_ _09379_/A _09379_/B vssd1 vssd1 vccd1 vccd1 _09380_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_62_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11410_ _11410_/A fanout5/X vssd1 vssd1 vccd1 vccd1 _11410_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12390_ hold282/A _12390_/B vssd1 vssd1 vccd1 vccd1 _12464_/B sky130_fd_sc_hd__or2_1
XFILLER_0_22_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11341_ _11341_/A _11341_/B vssd1 vssd1 vccd1 vccd1 _11554_/A sky130_fd_sc_hd__or2_4
XFILLER_0_62_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10246__A _11281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12164__C _12164_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11272_ _11514_/A _11272_/B vssd1 vssd1 vccd1 vccd1 _11274_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13011_ _13009_/Y _13011_/B vssd1 vssd1 vccd1 vccd1 _13012_/B sky130_fd_sc_hd__and2b_1
X_10223_ _10221_/X _10223_/B vssd1 vssd1 vccd1 vccd1 _10224_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_120_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10185__B1 _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07555__A _11709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09590__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ _10155_/B _10155_/C _10155_/A vssd1 vssd1 vccd1 vccd1 _10156_/A sky130_fd_sc_hd__a21oi_1
X_10085_ _10085_/A vssd1 vssd1 vccd1 vccd1 _10093_/A sky130_fd_sc_hd__inv_2
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09770__A _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10488__A1 _07310_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07889__C1 _09254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10488__B2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10987_ _10864_/B _10864_/C _11562_/A vssd1 vssd1 vccd1 vccd1 _10988_/B sky130_fd_sc_hd__a21oi_1
X_12726_ _12724_/A _12724_/B _12724_/C vssd1 vssd1 vccd1 vccd1 _12727_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_45_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12657_ _06824_/B _09516_/X _12657_/B1 reg1_val[28] _12799_/A2 vssd1 vssd1 vccd1
+ vccd1 _12657_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_25_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09929__B _12667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11608_ _11714_/A _11608_/B vssd1 vssd1 vccd1 vccd1 _11610_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_52_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12588_ _12586_/Y _12588_/B vssd1 vssd1 vccd1 vccd1 _12589_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_4_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07449__B _07476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11539_ _11537_/X _11539_/B vssd1 vssd1 vccd1 vccd1 _11540_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_52_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap148 _07420_/Y vssd1 vssd1 vccd1 vccd1 _09955_/A sky130_fd_sc_hd__buf_6
XFILLER_0_111_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13362__B1 _13555_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13209_ hold44/X hold268/X vssd1 vssd1 vccd1 vccd1 _13211_/A sky130_fd_sc_hd__nand2b_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07465__A _11508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _08907_/A _10049_/A2 _09173_/B2 _08197_/A vssd1 vssd1 vccd1 vccd1 _08751_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09869__B1 _12314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07701_ _07704_/B _07704_/A vssd1 vssd1 vccd1 vccd1 _07707_/B sky130_fd_sc_hd__nand2b_1
X_08681_ _08857_/A _08681_/B vssd1 vssd1 vccd1 vccd1 _08712_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07344__A1 _07476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07632_ _07633_/A _07633_/B vssd1 vssd1 vccd1 vccd1 _07632_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13417__A1 _11709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12310__S _12782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06809__A _06928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07563_ _07563_/A _07563_/B vssd1 vssd1 vccd1 vccd1 _07654_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09302_ _09301_/A _09301_/B _09303_/A vssd1 vssd1 vccd1 vccd1 _09302_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11979__A1 _12710_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11979__B2 _12537_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07494_ _07193_/A _07449_/Y _07448_/Y _07184_/D vssd1 vssd1 vccd1 vccd1 _07494_/X
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09233_ fanout40/X fanout68/X fanout66/X fanout56/X vssd1 vssd1 vccd1 vccd1 _09234_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_15_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13742_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_28_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09164_ _09288_/A _09165_/B vssd1 vssd1 vccd1 vccd1 _09289_/A sky130_fd_sc_hd__nor2_1
X_08115_ _08115_/A _08115_/B vssd1 vssd1 vccd1 vccd1 _08223_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08072__A2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09095_ _09094_/B _09094_/C _09094_/A vssd1 vssd1 vccd1 vccd1 _09095_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08046_ _10235_/A1 fanout74/X fanout70/X _10235_/B2 vssd1 vssd1 vccd1 vccd1 _08047_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07280__B1 _07281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07375__A _07634_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09572__A2 _10235_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09997_ _09664_/X _09667_/X _10004_/S vssd1 vssd1 vccd1 vccd1 _09997_/X sky130_fd_sc_hd__mux2_1
X_08948_ _08271_/A _07399_/Y _09910_/A1 _09501_/A vssd1 vssd1 vccd1 vccd1 _08949_/B
+ sky130_fd_sc_hd__a22o_1
X_08879_ _08879_/A _08879_/B vssd1 vssd1 vccd1 vccd1 _08898_/B sky130_fd_sc_hd__xnor2_2
X_10910_ _10910_/A _10910_/B vssd1 vssd1 vccd1 vccd1 _10931_/A sky130_fd_sc_hd__xnor2_1
X_11890_ _09529_/B _11877_/X _11889_/X _11871_/X vssd1 vssd1 vccd1 vccd1 _11890_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11419__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10841_ _10841_/A _10841_/B vssd1 vssd1 vccd1 vccd1 _10843_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13560_ _13591_/A hold270/X vssd1 vssd1 vccd1 vccd1 _13729_/D sky130_fd_sc_hd__and2_1
X_10772_ _11281_/A _10772_/B vssd1 vssd1 vccd1 vccd1 _10776_/A sky130_fd_sc_hd__xnor2_1
X_12511_ _12627_/A _12730_/A vssd1 vssd1 vccd1 vccd1 _12635_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_109_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13491_ hold253/X _13555_/A2 _13490_/X _13542_/B2 vssd1 vssd1 vccd1 vccd1 hold254/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12442_ _12442_/A _12442_/B _12508_/A vssd1 vssd1 vccd1 vccd1 _12443_/B sky130_fd_sc_hd__or3_1
XFILLER_0_35_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13592__B1 _13207_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12373_ _12373_/A _12373_/B vssd1 vssd1 vccd1 vccd1 _12733_/A sky130_fd_sc_hd__nand2_2
XANTENNA__10945__A2 _07891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11324_ _11163_/A _11163_/B _11162_/A vssd1 vssd1 vccd1 vccd1 _11329_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13344__B1 _13506_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11255_ _06943_/B _11587_/A2 _11254_/X vssd1 vssd1 vccd1 vccd1 _11255_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10206_ _12092_/A _10206_/B vssd1 vssd1 vccd1 vccd1 _10215_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11186_ _11638_/A _07643_/B fanout12/X _11527_/A vssd1 vssd1 vccd1 vccd1 _11187_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10137_ _10137_/A _10137_/B vssd1 vssd1 vccd1 vccd1 _10138_/B sky130_fd_sc_hd__xnor2_2
X_10068_ _10068_/A _10068_/B vssd1 vssd1 vccd1 vccd1 _10070_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_89_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10881__A1 _12648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08826__A1 _08866_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08826__B2 _08950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12709_ _12693_/A _12709_/A2 _09515_/Y _06815_/B _12708_/Y vssd1 vssd1 vccd1 vccd1
+ _12709_/X sky130_fd_sc_hd__a221o_1
XANTENNA__09659__B _09659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13689_ _13693_/CLK _13689_/D vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11270__A _11823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07179__B _09496_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold204 hold204/A vssd1 vssd1 vccd1 vccd1 hold204/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold215 hold215/A vssd1 vssd1 vccd1 vccd1 hold215/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07801__A2 _07544_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold226 hold226/A vssd1 vssd1 vccd1 vccd1 hold226/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 hold237/A vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09920_ _09922_/A _09922_/B vssd1 vssd1 vccd1 vccd1 _09923_/A sky130_fd_sc_hd__and2_1
Xhold248 hold248/A vssd1 vssd1 vccd1 vccd1 hold248/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold259 hold259/A vssd1 vssd1 vccd1 vccd1 hold259/X sky130_fd_sc_hd__buf_1
XFILLER_0_0_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09851_ _09712_/X _09850_/X _10176_/A vssd1 vssd1 vccd1 vccd1 _09851_/X sky130_fd_sc_hd__mux2_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08802_ _08820_/B vssd1 vssd1 vccd1 vccd1 _08802_/Y sky130_fd_sc_hd__inv_2
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _09951_/A _07240_/B fanout6/X _09781_/Y vssd1 vssd1 vccd1 vccd1 _09783_/B
+ sky130_fd_sc_hd__a31o_2
X_06994_ _06994_/A vssd1 vssd1 vccd1 vccd1 _06996_/A sky130_fd_sc_hd__inv_2
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08733_ _08857_/A _08733_/B vssd1 vssd1 vccd1 vccd1 _08739_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08664_ _09948_/A _08664_/B vssd1 vssd1 vccd1 vccd1 _08670_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__10321__B1 _12537_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07134__S _07135_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07615_ _07616_/A _07616_/B vssd1 vssd1 vccd1 vccd1 _07615_/Y sky130_fd_sc_hd__nand2_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08595_ _08873_/A2 _10522_/A _09885_/B1 _08891_/B vssd1 vssd1 vccd1 vccd1 _08596_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07546_ _07546_/A _11157_/A vssd1 vssd1 vccd1 vccd1 _07546_/X sky130_fd_sc_hd__or2_4
XFILLER_0_72_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08817__A1 _09671_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07477_ _07478_/A _07478_/B vssd1 vssd1 vccd1 vccd1 _07477_/X sky130_fd_sc_hd__and2_4
XFILLER_0_63_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11180__A _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09216_ _07347_/X fanout35/X _07699_/B _09216_/B2 vssd1 vssd1 vccd1 vccd1 _09217_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_119_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09147_ _08271_/A _12667_/A _10536_/A2 _09501_/A vssd1 vssd1 vccd1 vccd1 _09148_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09242__A1 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07089__B _09703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09242__B2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09585__A _09948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09078_ _09060_/B _09060_/C _09068_/X _09079_/B vssd1 vssd1 vccd1 vccd1 _09080_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__09793__A2 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13326__B1 _13450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08029_ _08028_/A _08108_/A _08028_/B _08026_/A vssd1 vssd1 vccd1 vccd1 _08038_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout93_A _11719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11040_ _11041_/A _11041_/B vssd1 vssd1 vccd1 vccd1 _11161_/B sky130_fd_sc_hd__or2_1
XANTENNA__07833__A _09161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12991_ _12989_/Y _12991_/B vssd1 vssd1 vccd1 vccd1 _12992_/B sky130_fd_sc_hd__nand2b_2
X_11942_ _11942_/A _11942_/B vssd1 vssd1 vccd1 vccd1 _11944_/C sky130_fd_sc_hd__xnor2_2
XANTENNA__07859__A2 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11873_ reg1_val[18] curr_PC[18] vssd1 vssd1 vccd1 vccd1 _11874_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_86_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13612_ _13717_/CLK hold8/X vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfxtp_1
X_10824_ _10937_/B _10824_/B vssd1 vssd1 vccd1 vccd1 _10827_/B sky130_fd_sc_hd__and2_1
XANTENNA__08808__A1 _08873_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08808__B2 _08891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08664__A _09948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11802__B _11802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13543_ _13543_/A _13543_/B vssd1 vssd1 vccd1 vccd1 _13725_/D sky130_fd_sc_hd__and2_1
XFILLER_0_39_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10755_ _06973_/B _11587_/A2 _10753_/Y _10754_/X vssd1 vssd1 vccd1 vccd1 _10755_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13474_ _13474_/A _13474_/B vssd1 vssd1 vccd1 vccd1 _13474_/Y sky130_fd_sc_hd__xnor2_1
X_10686_ _10686_/A _10686_/B vssd1 vssd1 vccd1 vccd1 _10703_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12425_ _12426_/A _12426_/B _12426_/C vssd1 vssd1 vccd1 vccd1 _12502_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__09233__A1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09233__B2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10918__A2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12356_ _12437_/A _12356_/B vssd1 vssd1 vccd1 vccd1 _12358_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_23_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11307_ _11307_/A _11307_/B _11307_/C vssd1 vssd1 vccd1 vccd1 _11308_/B sky130_fd_sc_hd__or3_1
X_12287_ _12287_/A vssd1 vssd1 vccd1 vccd1 _12288_/B sky130_fd_sc_hd__inv_2
X_11238_ _11237_/A _11237_/B _11237_/Y _12047_/C1 vssd1 vssd1 vccd1 vccd1 _11238_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12540__A1 _12518_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11169_ _12253_/A _11169_/B vssd1 vssd1 vccd1 vccd1 _11171_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07400_ _10004_/S _07400_/B vssd1 vssd1 vccd1 vccd1 _13147_/A sky130_fd_sc_hd__xnor2_4
X_08380_ _08380_/A _08380_/B vssd1 vssd1 vccd1 vccd1 _08453_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07331_ reg1_val[18] reg1_val[19] _07435_/B vssd1 vssd1 vccd1 vccd1 _13082_/B sky130_fd_sc_hd__or3_4
XANTENNA__08275__A2 _07300_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07262_ _07264_/A _07264_/B vssd1 vssd1 vccd1 vccd1 _07644_/B sky130_fd_sc_hd__or2_1
XFILLER_0_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09001_ _09001_/A _09001_/B vssd1 vssd1 vccd1 vccd1 _09002_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_115_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07193_ _07193_/A _07193_/B _07192_/C vssd1 vssd1 vccd1 vccd1 _07287_/A sky130_fd_sc_hd__or3b_4
XFILLER_0_14_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11031__A1 wire101/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11031__B2 _11922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09903_ _11507_/A _09903_/B vssd1 vssd1 vccd1 vccd1 _09907_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09527__A2 _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11159__B _11307_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09834_ _12742_/A _09004_/A _09006_/B _11866_/A _09833_/Y vssd1 vssd1 vccd1 vccd1
+ _09834_/X sky130_fd_sc_hd__o311a_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08749__A _09371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _09765_/A _09765_/B vssd1 vssd1 vccd1 vccd1 _09766_/B sky130_fd_sc_hd__nand2_1
X_06977_ _13015_/A _07492_/A vssd1 vssd1 vccd1 vccd1 _06977_/Y sky130_fd_sc_hd__nor2_1
X_08716_ _08761_/A _08761_/B _08713_/X vssd1 vssd1 vccd1 vccd1 _08730_/A sky130_fd_sc_hd__o21a_1
X_09696_ _09696_/A _09696_/B vssd1 vssd1 vccd1 vccd1 _09697_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08647_ _08647_/A _08647_/B vssd1 vssd1 vccd1 vccd1 _08697_/B sky130_fd_sc_hd__xnor2_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11903__A _12421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08578_ _07399_/Y _07541_/X _07545_/Y _09910_/A1 vssd1 vssd1 vccd1 vccd1 _08579_/B
+ sky130_fd_sc_hd__a22o_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07529_ _09591_/A _07529_/B vssd1 vssd1 vccd1 vccd1 _07552_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10540_ _10541_/B _10541_/C _09575_/A vssd1 vssd1 vccd1 vccd1 _10542_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_107_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10471_ reg1_val[6] curr_PC[6] vssd1 vssd1 vccd1 vccd1 _10472_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_91_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12210_ _12440_/B _12210_/B vssd1 vssd1 vccd1 vccd1 _12372_/C sky130_fd_sc_hd__xnor2_4
XFILLER_0_32_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11022__A1 _12825_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13190_ _12189_/A _13196_/A2 hold49/X _13591_/A vssd1 vssd1 vccd1 vccd1 hold50/A
+ sky130_fd_sc_hd__o211a_1
X_12141_ _12052_/A _12052_/B _12050_/B vssd1 vssd1 vccd1 vccd1 _12142_/B sky130_fd_sc_hd__o21a_1
X_12072_ _10342_/A _12068_/X _12071_/X vssd1 vssd1 vccd1 vccd1 dest_val[20] sky130_fd_sc_hd__o21ai_4
X_11023_ _10900_/Y _10984_/X _11864_/A vssd1 vssd1 vccd1 vccd1 _11115_/A sky130_fd_sc_hd__o21ai_1
X_12974_ _12974_/A _12974_/B vssd1 vssd1 vccd1 vccd1 _12976_/A sky130_fd_sc_hd__nor2_2
X_11925_ _11925_/A _11925_/B vssd1 vssd1 vccd1 vccd1 _11940_/A sky130_fd_sc_hd__xor2_2
XANTENNA_clkbuf_4_0_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11856_ _11856_/A _11948_/A vssd1 vssd1 vccd1 vccd1 _12037_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08394__A _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10807_ _10808_/A _10808_/B vssd1 vssd1 vccd1 vccd1 _10809_/A sky130_fd_sc_hd__or2_1
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11787_ hold231/A _11878_/C _12311_/B1 vssd1 vssd1 vccd1 vccd1 _11788_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11261__A1 _12537_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10738_ _10620_/A _10617_/Y _10619_/B vssd1 vssd1 vccd1 vccd1 _10742_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_82_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13526_ _13539_/A hold293/X vssd1 vssd1 vccd1 vccd1 _13721_/D sky130_fd_sc_hd__and2_1
XANTENNA__11261__B2 _12760_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13457_ hold262/X _13456_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13457_/X sky130_fd_sc_hd__mux2_1
X_10669_ _10669_/A _10669_/B vssd1 vssd1 vccd1 vccd1 _10684_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_113_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12408_ _07257_/X fanout8/X fanout3/X _12496_/A vssd1 vssd1 vccd1 vccd1 _12409_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07738__A _10239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13388_ hold76/X _13416_/A2 _13420_/B1 hold101/X _13383_/A vssd1 vssd1 vccd1 vccd1
+ hold102/A sky130_fd_sc_hd__o221a_1
XFILLER_0_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12761__A1 _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12339_ _12496_/A fanout8/X fanout3/X _12413_/A vssd1 vssd1 vccd1 vccd1 _12340_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06991__A2 _07110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06900_ reg1_val[17] _07300_/A vssd1 vssd1 vccd1 vccd1 _06902_/A sky130_fd_sc_hd__or2_1
X_07880_ _11731_/A _07880_/B vssd1 vssd1 vccd1 vccd1 _07882_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10524__B1 _07522_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06831_ _06831_/A _06831_/B vssd1 vssd1 vccd1 vccd1 _12452_/A sky130_fd_sc_hd__nor2_2
X_09550_ _10225_/A _07643_/B fanout13/X _10104_/A vssd1 vssd1 vccd1 vccd1 _09551_/B
+ sky130_fd_sc_hd__a22o_1
X_06762_ _10734_/A vssd1 vssd1 vccd1 vccd1 _06762_/Y sky130_fd_sc_hd__inv_2
X_08501_ _08501_/A _08501_/B vssd1 vssd1 vccd1 vccd1 _08510_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09142__B1 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09481_ _09473_/X _10172_/B _10176_/A vssd1 vssd1 vccd1 vccd1 _09481_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12819__A _12995_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08432_ _09373_/A _08432_/B vssd1 vssd1 vccd1 vccd1 _08436_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06817__A _06886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08363_ _08364_/A _08364_/B vssd1 vssd1 vccd1 vccd1 _08363_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout143_A _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07314_ _10078_/A _07314_/B vssd1 vssd1 vccd1 vccd1 _07721_/B sky130_fd_sc_hd__xnor2_1
X_08294_ _08294_/A _08294_/B vssd1 vssd1 vccd1 vccd1 _08302_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_34_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07245_ _07245_/A _07245_/B vssd1 vssd1 vccd1 vccd1 _07687_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_116_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12554__A _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07176_ _11463_/A _07398_/B vssd1 vssd1 vccd1 vccd1 _07594_/B sky130_fd_sc_hd__and2_4
XFILLER_0_42_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09582__B _10787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08479__A _09948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08184__A1 _13149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08184__B2 _08923_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09817_ _09817_/A _09817_/B vssd1 vssd1 vccd1 vccd1 _09819_/B sky130_fd_sc_hd__xnor2_2
X_09748_ _09748_/A _10518_/A vssd1 vssd1 vccd1 vccd1 _09755_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09133__B1 _07545_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10818__A1 _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _09468_/X _09470_/X _09688_/S vssd1 vssd1 vccd1 vccd1 _09679_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10818__B2 _12103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _11710_/A _11710_/B vssd1 vssd1 vccd1 vccd1 _11712_/B sky130_fd_sc_hd__xnor2_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11491__A1 _12867_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _12733_/C _12688_/X _12689_/Y vssd1 vssd1 vccd1 vccd1 _12690_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09103__A _12421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11641_ _11642_/A _11642_/B vssd1 vssd1 vccd1 vccd1 _11641_/X sky130_fd_sc_hd__and2b_1
XANTENNA__09436__A1 _13129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09987__A2 _09650_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11572_ _11572_/A _11572_/B vssd1 vssd1 vccd1 vccd1 _11574_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08942__A _09659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13311_ _13574_/B _13311_/B vssd1 vssd1 vccd1 vccd1 _13579_/C sky130_fd_sc_hd__and2b_1
X_10523_ _10523_/A _10523_/B vssd1 vssd1 vccd1 vccd1 _10552_/A sky130_fd_sc_hd__xnor2_1
X_13242_ hold37/X hold257/X vssd1 vssd1 vccd1 vccd1 _13244_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_122_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10454_ _09843_/X _09848_/X _10600_/S vssd1 vssd1 vccd1 vccd1 _10454_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13173_ hold66/X _13191_/B vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__or2_1
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10385_ fanout56/X fanout25/X fanout23/X fanout53/X vssd1 vssd1 vccd1 vccd1 _10386_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_103_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10754__B1 _12748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12124_ _11947_/Y _12290_/A _12122_/Y vssd1 vssd1 vccd1 vccd1 _12124_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_102_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12055_ _12056_/B _12056_/A hold212/A vssd1 vssd1 vccd1 vccd1 _12055_/Y sky130_fd_sc_hd__o21bai_1
XANTENNA__10506__B1 _07546_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09372__B1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11006_ _13651_/Q _11693_/A2 _11248_/C _11005_/Y _12533_/B1 vssd1 vssd1 vccd1 vccd1
+ _11014_/A sky130_fd_sc_hd__a311o_1
XANTENNA__11527__B _11802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09124__B1 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09712__S _10004_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12957_ _12949_/B _12954_/B _12947_/X vssd1 vssd1 vccd1 vccd1 _12958_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_59_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11482__A1 _07513_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11908_ fanout20/X fanout10/X fanout5/X fanout18/X vssd1 vssd1 vccd1 vccd1 _11909_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12888_ reg1_val[13] curr_PC[13] _12978_/S vssd1 vssd1 vccd1 vccd1 _12890_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_74_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11839_ _11935_/A _11839_/B vssd1 vssd1 vccd1 vccd1 _11841_/B sky130_fd_sc_hd__and2_1
XFILLER_0_23_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09948__A _09948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13509_ _13509_/A _13509_/B vssd1 vssd1 vccd1 vccd1 _13509_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10993__B1 _12047_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07030_ _09501_/A _13145_/A vssd1 vssd1 vccd1 vccd1 _09701_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_24_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13189__B _13191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08981_ _08981_/A _08981_/B vssd1 vssd1 vccd1 vccd1 _09055_/A sky130_fd_sc_hd__nand2_1
X_07932_ _07300_/Y _07545_/Y _11638_/A _07541_/X vssd1 vssd1 vccd1 vccd1 _07933_/B
+ sky130_fd_sc_hd__a22o_1
X_07863_ _07861_/X _07863_/B vssd1 vssd1 vccd1 vccd1 _07864_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__09902__A2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07634__C _07634_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07913__A1 _10104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07913__B2 _10225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09602_ _09602_/A _09726_/A _09602_/C vssd1 vssd1 vccd1 vccd1 _09726_/B sky130_fd_sc_hd__nand3_1
X_06814_ reg1_val[29] _09254_/B vssd1 vssd1 vccd1 vccd1 _06815_/B sky130_fd_sc_hd__and2_1
X_07794_ _11047_/A fanout75/X _08704_/B fanout85/X vssd1 vssd1 vccd1 vccd1 _07795_/B
+ sky130_fd_sc_hd__o22a_1
X_09533_ _10457_/S _09536_/B vssd1 vssd1 vccd1 vccd1 _09534_/C sky130_fd_sc_hd__or2_4
X_06745_ instruction[3] vssd1 vssd1 vccd1 vccd1 _09524_/A sky130_fd_sc_hd__inv_2
XANTENNA__12549__A _12666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09464_ _09462_/X _09463_/X _09674_/S vssd1 vssd1 vccd1 vccd1 _09464_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12268__B _12666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08415_ _08415_/A _08415_/B vssd1 vssd1 vccd1 vccd1 _08463_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_59_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09395_ _09395_/A vssd1 vssd1 vccd1 vccd1 _09402_/A sky130_fd_sc_hd__inv_2
XFILLER_0_80_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08346_ _08355_/A _08355_/B vssd1 vssd1 vccd1 vccd1 _08357_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_117_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08277_ _08274_/B _08274_/C _08274_/A vssd1 vssd1 vccd1 vccd1 _08278_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07228_ _07212_/B _07213_/A _07212_/C _07521_/A vssd1 vssd1 vccd1 vccd1 _07230_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_0_6_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07159_ reg1_val[4] _07265_/D vssd1 vssd1 vccd1 vccd1 _07160_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_30_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10170_ _10170_/A _10170_/B vssd1 vssd1 vccd1 vccd1 _10170_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout130 _07285_/Y vssd1 vssd1 vccd1 vccd1 _08891_/B sky130_fd_sc_hd__clkbuf_8
Xfanout141 _11231_/A vssd1 vssd1 vccd1 vccd1 _12311_/B1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09354__B1 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout152 _13147_/A vssd1 vssd1 vccd1 vccd1 _08873_/B2 sky130_fd_sc_hd__buf_6
Xfanout163 _13142_/Y vssd1 vssd1 vccd1 vccd1 _13196_/A2 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08002__A _11286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout174 _10236_/A vssd1 vssd1 vccd1 vccd1 _10095_/A sky130_fd_sc_hd__buf_12
Xfanout185 _13550_/A2 vssd1 vssd1 vccd1 vccd1 _13450_/B sky130_fd_sc_hd__buf_4
Xfanout196 _09508_/Y vssd1 vssd1 vccd1 vccd1 _12709_/A2 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13438__C1 _13568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09106__B1 _13151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12811_ reg1_val[2] curr_PC[2] _12825_/S vssd1 vssd1 vccd1 vccd1 _12813_/B sky130_fd_sc_hd__mux2_1
XANTENNA__13453__A2 fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10267__A2 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12742_ _12742_/A _12742_/B vssd1 vssd1 vccd1 vccd1 _12743_/B sky130_fd_sc_hd__nor2_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _12724_/A _12673_/B vssd1 vssd1 vccd1 vccd1 _12675_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_127_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ _11731_/A _11624_/B vssd1 vssd1 vccd1 vccd1 _11628_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09768__A _11508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11767__A2 _12163_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11555_ _11344_/Y _11763_/A _11553_/X vssd1 vssd1 vccd1 vccd1 _11555_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08632__A2 _07477_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06904__B _12981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10506_ fanout51/X _10787_/A _07546_/X _12557_/B vssd1 vssd1 vccd1 vccd1 _10507_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_80_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11486_ _12760_/A1 _11474_/X _11485_/X _11466_/X vssd1 vssd1 vccd1 vccd1 _11486_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12716__A1 _11823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13225_ _13225_/A _13225_/B vssd1 vssd1 vccd1 vccd1 _13561_/A sky130_fd_sc_hd__nor2_1
X_10437_ _09823_/X _09983_/X _09984_/X _10631_/A _10857_/A vssd1 vssd1 vccd1 vccd1
+ _10438_/B sky130_fd_sc_hd__a2111oi_1
XFILLER_0_21_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09593__B1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13156_ _10225_/A _13196_/A2 hold79/X _13547_/A vssd1 vssd1 vccd1 vccd1 hold80/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10368_ _10369_/A _10369_/B vssd1 vssd1 vccd1 vccd1 _10520_/A sky130_fd_sc_hd__nor2_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06946__A2 _06936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ _12107_/A _12107_/B vssd1 vssd1 vccd1 vccd1 _12108_/B sky130_fd_sc_hd__and2_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ reg1_val[21] _13129_/B vssd1 vssd1 vccd1 vccd1 _13088_/B sky130_fd_sc_hd__nand2_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10299_ _09654_/A _09654_/B _10298_/X vssd1 vssd1 vccd1 vccd1 _10302_/A sky130_fd_sc_hd__a21o_1
X_12038_ _11668_/B _12037_/X _12369_/A vssd1 vssd1 vccd1 vccd1 _12368_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__07751__A _10266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13444__A2 _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11455__A1 _10984_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08200_ _08199_/B _08199_/C _09949_/A vssd1 vssd1 vccd1 vccd1 _08201_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_7_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09180_ _09301_/A _09180_/B vssd1 vssd1 vccd1 vccd1 _09182_/B sky130_fd_sc_hd__or2_1
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12404__B1 _12379_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08131_ _10119_/A _08224_/B _08224_/A vssd1 vssd1 vccd1 vccd1 _08152_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_16_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10617__A _13015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06814__B _09254_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08062_ _09949_/A _08062_/B vssd1 vssd1 vccd1 vccd1 _08064_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07831__B1 _13149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07013_ _06928_/A _06936_/B _12995_/B _07011_/X vssd1 vssd1 vccd1 vccd1 _07013_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08387__A1 _10225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout106_A _07557_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08387__B2 _07556_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09584__B1 _09948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10194__A1 _09839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06937__A2 _06980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08964_ _08964_/A _08964_/B vssd1 vssd1 vccd1 vccd1 _09012_/B sky130_fd_sc_hd__nor2_1
X_07915_ _07915_/A vssd1 vssd1 vccd1 vccd1 _07924_/A sky130_fd_sc_hd__inv_2
X_08895_ _10236_/A _08902_/A vssd1 vssd1 vccd1 vccd1 _08896_/D sky130_fd_sc_hd__nor2_1
X_07846_ _08036_/A _08036_/B vssd1 vssd1 vccd1 vccd1 _08037_/A sky130_fd_sc_hd__or2_1
XFILLER_0_98_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07661__A _09575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07777_ _07841_/A _07841_/B _07748_/X vssd1 vssd1 vccd1 vccd1 _07784_/A sky130_fd_sc_hd__a21o_1
XANTENNA__13435__A2 _13598_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09516_ _09516_/A _09516_/B vssd1 vssd1 vccd1 vccd1 _09516_/X sky130_fd_sc_hd__or2_2
XFILLER_0_94_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09447_ reg1_val[4] reg1_val[27] _09463_/S vssd1 vssd1 vccd1 vccd1 _09447_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11911__A _12253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09378_ _09379_/A _09379_/B vssd1 vssd1 vccd1 vccd1 _09378_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_47_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout19_A _07493_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08329_ _09950_/A _08329_/B vssd1 vssd1 vccd1 vccd1 _08333_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10527__A _12421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11340_ _11340_/A _11340_/B _11340_/C vssd1 vssd1 vccd1 vccd1 _11341_/B sky130_fd_sc_hd__and3_1
XFILLER_0_104_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11271_ _12087_/A _07416_/X _07422_/Y _12103_/A vssd1 vssd1 vccd1 vccd1 _11272_/B
+ sky130_fd_sc_hd__o22a_1
X_13010_ reg1_val[6] _13010_/B vssd1 vssd1 vccd1 vccd1 _13011_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_120_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10222_ _10222_/A _10222_/B _10098_/Y vssd1 vssd1 vccd1 vccd1 _10223_/B sky130_fd_sc_hd__or3b_2
X_10153_ _10433_/A _09827_/X _10577_/A _10152_/X vssd1 vssd1 vccd1 vccd1 _10155_/C
+ sky130_fd_sc_hd__o31a_1
X_10084_ _11709_/A _10084_/B vssd1 vssd1 vccd1 vccd1 _10085_/A sky130_fd_sc_hd__xnor2_1
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07889__B1 _07476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10488__A2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12189__A _12189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13426__A2 _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10986_ _11864_/A _10900_/Y _10984_/X _11955_/A vssd1 vssd1 vccd1 vccd1 _10986_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_0_29_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12725_ _12727_/A vssd1 vssd1 vccd1 vccd1 _12725_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12656_ _12656_/A _12656_/B _12754_/C vssd1 vssd1 vccd1 vccd1 _12656_/X sky130_fd_sc_hd__and3_1
XFILLER_0_72_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11607_ _11607_/A _11607_/B vssd1 vssd1 vccd1 vccd1 _11608_/B sky130_fd_sc_hd__or2_1
X_12587_ reg1_val[27] curr_PC[27] vssd1 vssd1 vccd1 vccd1 _12588_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_108_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11538_ _11538_/A _11538_/B _11536_/Y vssd1 vssd1 vccd1 vccd1 _11539_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13748__A _13748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11469_ _11469_/A _11469_/B vssd1 vssd1 vccd1 vccd1 _11471_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_123_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13208_ fanout7/X _13598_/C hold173/X _13605_/A vssd1 vssd1 vccd1 vccd1 _13640_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11268__A _12372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13139_ _13142_/A hold192/X vssd1 vssd1 vccd1 vccd1 _13140_/C sky130_fd_sc_hd__nor2_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07184__C _10889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07700_ _10050_/A _07700_/B vssd1 vssd1 vccd1 vccd1 _07704_/B sky130_fd_sc_hd__xnor2_1
X_08680_ _08806_/B1 _10104_/A _07420_/Y _08806_/A2 vssd1 vssd1 vccd1 vccd1 _08681_/B
+ sky130_fd_sc_hd__a22o_1
X_07631_ _07940_/B _07631_/B vssd1 vssd1 vccd1 vccd1 _07633_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10884__C1 _12533_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06809__B _13054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07562_ _10263_/A _07562_/B vssd1 vssd1 vccd1 vccd1 _07654_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_76_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09301_ _09301_/A _09301_/B vssd1 vssd1 vccd1 vccd1 _09303_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_75_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07493_ _11991_/A _07493_/B vssd1 vssd1 vccd1 vccd1 _07493_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_76_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12827__A _13000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09232_ _10078_/A _09232_/B vssd1 vssd1 vccd1 vccd1 _09239_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__11731__A _11731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09163_ _11731_/A _09163_/B vssd1 vssd1 vccd1 vccd1 _09165_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08114_ _08116_/A _08116_/B vssd1 vssd1 vccd1 vccd1 _08114_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_43_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07804__B1 _10814_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09094_ _09094_/A _09094_/B _09094_/C vssd1 vssd1 vccd1 vccd1 _09097_/A sky130_fd_sc_hd__and3_1
XFILLER_0_4_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11877__S _12525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08045_ _08155_/A _08155_/B _08042_/X vssd1 vssd1 vccd1 vccd1 _08090_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_114_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11178__A _11709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09996_ _09996_/A _09996_/B vssd1 vssd1 vccd1 vccd1 _09996_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_110_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08947_ _08945_/Y _08947_/B vssd1 vssd1 vccd1 vccd1 _09010_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__11116__B1 _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10810__A wire122/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08878_ _08898_/A vssd1 vssd1 vccd1 vccd1 _08878_/Y sky130_fd_sc_hd__inv_2
X_07829_ _07996_/A _07996_/B _07825_/X vssd1 vssd1 vccd1 vccd1 _07836_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_98_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10840_ _10840_/A _10840_/B vssd1 vssd1 vccd1 vccd1 _10841_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11419__A1 _11638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11419__B2 _11527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10890__A2 _11688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10771_ fanout51/X fanout84/X fanout79/X _12557_/B vssd1 vssd1 vccd1 vccd1 _10772_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_66_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_5_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12510_ _12210_/B _12368_/C _12508_/X _12509_/X vssd1 vssd1 vccd1 vccd1 _12730_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13490_ hold295/A _13489_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13490_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12441_ _12288_/A _12361_/Y _12363_/B vssd1 vssd1 vccd1 vccd1 _12441_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__08048__B1 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12372_ _12372_/A _12372_/B _12372_/C _12372_/D vssd1 vssd1 vccd1 vccd1 _12373_/B
+ sky130_fd_sc_hd__nor4_2
XANTENNA__08950__A _09671_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11323_ _11211_/A _11211_/B _11210_/A vssd1 vssd1 vccd1 vccd1 _11331_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13568__A _13568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09548__B1 _07557_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11254_ _07476_/A _11793_/B _12657_/B1 reg1_val[12] vssd1 vssd1 vccd1 vccd1 _11254_/X
+ sky130_fd_sc_hd__o22a_1
X_10205_ fanout14/X _07477_/X _11309_/A _07833_/B vssd1 vssd1 vccd1 vccd1 _10206_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11185_ _11185_/A _11185_/B vssd1 vssd1 vccd1 vccd1 _11193_/A sky130_fd_sc_hd__xor2_1
X_10136_ _10134_/A _10134_/B _10137_/B vssd1 vssd1 vccd1 vccd1 _10136_/X sky130_fd_sc_hd__a21o_1
X_10067_ _10068_/A _10068_/B vssd1 vssd1 vccd1 vccd1 _10217_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_106_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08826__A2 _09216_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10969_ _10970_/B _10970_/A vssd1 vssd1 vccd1 vccd1 _10969_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10094__B1 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12708_ _06815_/A _09520_/X _11688_/B reg1_val[29] _12799_/A2 vssd1 vssd1 vccd1 vccd1
+ _12708_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_0_85_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13688_ _13701_/CLK _13688_/D vssd1 vssd1 vccd1 vccd1 hold136/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12639_ _06801_/Y _06840_/A _06802_/A vssd1 vssd1 vccd1 vccd1 _12639_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_115_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07179__C _10007_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold205 hold229/X vssd1 vssd1 vccd1 vccd1 hold205/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold216 hold216/A vssd1 vssd1 vccd1 vccd1 hold216/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 hold227/A vssd1 vssd1 vccd1 vccd1 hold227/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold238 hold238/A vssd1 vssd1 vccd1 vccd1 hold238/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 hold249/A vssd1 vssd1 vccd1 vccd1 hold249/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13197__B _13207_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09850_ _09487_/X _09491_/X _10007_/S vssd1 vssd1 vccd1 vccd1 _09850_/X sky130_fd_sc_hd__mux2_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ _09371_/A _08801_/B vssd1 vssd1 vccd1 vccd1 _08820_/B sky130_fd_sc_hd__xnor2_2
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _07240_/A fanout6/X _09951_/A vssd1 vssd1 vccd1 vccd1 _09781_/Y sky130_fd_sc_hd__a21oi_1
X_06993_ reg1_val[5] _06995_/B vssd1 vssd1 vccd1 vccd1 _06994_/A sky130_fd_sc_hd__nand2_2
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ _08806_/A2 _09910_/A1 _07420_/Y _08806_/B1 vssd1 vssd1 vccd1 vccd1 _08733_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12846__A0 _13015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ _07175_/X _07492_/Y _10637_/A _08933_/B vssd1 vssd1 vccd1 vccd1 _08664_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10321__A1 _12648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07614_ _10095_/A _07614_/B vssd1 vssd1 vccd1 vccd1 _07616_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08594_ _08746_/A _08594_/B vssd1 vssd1 vccd1 vccd1 _08600_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07545_ _07546_/A _11157_/A vssd1 vssd1 vccd1 vccd1 _07545_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08817__A2 _08778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12557__A _12557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07476_ _07476_/A _07476_/B _07476_/C vssd1 vssd1 vccd1 vccd1 _07478_/B sky130_fd_sc_hd__or3_4
XFILLER_0_29_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09215_ _10119_/A _09215_/B vssd1 vssd1 vccd1 vccd1 _09219_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09146_ _09146_/A _09146_/B vssd1 vssd1 vccd1 vccd1 _09146_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__08770__A _09373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09242__A2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09077_ _09077_/A _09077_/B vssd1 vssd1 vccd1 vccd1 _09079_/B sky130_fd_sc_hd__or2_1
XFILLER_0_71_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10805__A _11719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08028_ _08028_/A _08028_/B vssd1 vssd1 vccd1 vccd1 _08108_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_102_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08202__B1 _10814_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout86_A _11709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ _09979_/A _09979_/B vssd1 vssd1 vccd1 vccd1 _09981_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11636__A _11825_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07833__B _07833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12990_ reg1_val[2] _12990_/B vssd1 vssd1 vccd1 vccd1 _12991_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_99_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11941_ _11942_/A _11942_/B vssd1 vssd1 vccd1 vccd1 _12032_/B sky130_fd_sc_hd__and2_1
XFILLER_0_98_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11872_ reg1_val[18] curr_PC[18] vssd1 vssd1 vccd1 vccd1 _11874_/A sky130_fd_sc_hd__or2_1
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13611_ _13708_/CLK hold10/X vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12065__A1 _12710_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10823_ _10823_/A _10823_/B vssd1 vssd1 vccd1 vccd1 _10824_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08808__A2 _13149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12065__B2 _12537_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13542_ hold275/X _13555_/A2 _13541_/X _13542_/B2 vssd1 vssd1 vccd1 vccd1 _13543_/B
+ sky130_fd_sc_hd__a22o_1
X_10754_ hold295/A _12058_/A _10885_/B _12748_/B1 vssd1 vssd1 vccd1 vccd1 _10754_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10685_ _10685_/A _10685_/B vssd1 vssd1 vccd1 vccd1 _10704_/A sky130_fd_sc_hd__nand2_1
X_13473_ _13269_/X _13473_/B vssd1 vssd1 vccd1 vccd1 _13474_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_35_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09769__B1 _08486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12424_ _12491_/B _12424_/B vssd1 vssd1 vccd1 vccd1 _12426_/C sky130_fd_sc_hd__nand2_1
XANTENNA__09233__A2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12355_ _12355_/A _12355_/B vssd1 vssd1 vccd1 vccd1 _12356_/B sky130_fd_sc_hd__or2_1
XFILLER_0_50_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11306_ _11307_/A _11307_/B _11307_/C vssd1 vssd1 vccd1 vccd1 _11308_/A sky130_fd_sc_hd__o21ai_1
X_12286_ _12286_/A _12286_/B _12286_/C vssd1 vssd1 vccd1 vccd1 _12287_/A sky130_fd_sc_hd__and3_1
XFILLER_0_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11237_ _11237_/A _11237_/B vssd1 vssd1 vccd1 vccd1 _11237_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09941__B1 _08704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12540__A2 _12519_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11168_ _12103_/A fanout38/X fanout36/X fanout54/X vssd1 vssd1 vccd1 vccd1 _11169_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_93_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10119_ _10119_/A _10119_/B vssd1 vssd1 vccd1 vccd1 _10121_/B sky130_fd_sc_hd__xnor2_1
X_11099_ _11099_/A _11099_/B vssd1 vssd1 vccd1 vccd1 _11101_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11500__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08855__A _09950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07330_ reg1_val[18] reg1_val[19] _07435_/B vssd1 vssd1 vccd1 vccd1 _07337_/B sky130_fd_sc_hd__nor3_2
XANTENNA__11281__A _11281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07261_ _07261_/A _07261_/B vssd1 vssd1 vccd1 vccd1 _07264_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08680__B1 _07420_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09000_ _08991_/X _08993_/X _09318_/B _09318_/C _08167_/X vssd1 vssd1 vccd1 vccd1
+ _09001_/B sky130_fd_sc_hd__a2111o_1
XFILLER_0_116_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07192_ _07192_/A _07192_/B _07192_/C vssd1 vssd1 vccd1 vccd1 _07213_/A sky130_fd_sc_hd__and3_4
XANTENNA__08590__A _09371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11031__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10344__B _10727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09902_ _11732_/A fanout27/X fanout70/X fanout29/X vssd1 vssd1 vccd1 vccd1 _09903_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12840__A _13010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09833_ _12742_/A _09006_/B _09005_/Y vssd1 vssd1 vccd1 vccd1 _09833_/Y sky130_fd_sc_hd__o21bai_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09764_ _09765_/A _09765_/B vssd1 vssd1 vccd1 vccd1 _09766_/A sky130_fd_sc_hd__or2_1
X_06976_ _07492_/A _13015_/A vssd1 vssd1 vccd1 vccd1 _06976_/Y sky130_fd_sc_hd__nand2b_1
X_08715_ _08715_/A _08715_/B vssd1 vssd1 vccd1 vccd1 _08761_/B sky130_fd_sc_hd__xnor2_2
X_09695_ _09695_/A _09695_/B vssd1 vssd1 vccd1 vccd1 _09696_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_83_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08646_ _08646_/A _08646_/B vssd1 vssd1 vccd1 vccd1 _08697_/A sky130_fd_sc_hd__xnor2_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08577_ _08577_/A _08577_/B vssd1 vssd1 vccd1 vccd1 _08613_/A sky130_fd_sc_hd__xnor2_1
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07528_ fanout83/X _07522_/Y fanout79/X _11423_/A vssd1 vssd1 vccd1 vccd1 _07529_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07459_ reg1_val[15] _07513_/A vssd1 vssd1 vccd1 vccd1 _11585_/A sky130_fd_sc_hd__xor2_1
XANTENNA__09596__A _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10470_ reg1_val[6] curr_PC[6] vssd1 vssd1 vccd1 vccd1 _10470_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09129_ _09129_/A _09129_/B vssd1 vssd1 vccd1 vccd1 _09130_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_115_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10230__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12140_ _12140_/A _12140_/B vssd1 vssd1 vccd1 vccd1 _12142_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_114_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08005__A _10944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12071_ _12327_/A _12071_/B _12160_/B vssd1 vssd1 vccd1 vccd1 _12071_/X sky130_fd_sc_hd__or3_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11022_ _12825_/S _11018_/X _11019_/X _11021_/Y vssd1 vssd1 vccd1 vccd1 dest_val[10]
+ sky130_fd_sc_hd__a22o_4
XANTENNA__11730__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12973_ _12979_/A _12973_/B vssd1 vssd1 vccd1 vccd1 _12974_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_87_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11924_ _11924_/A _11924_/B vssd1 vssd1 vccd1 vccd1 _11925_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_87_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11855_ _11659_/Y _11757_/Y _11759_/B vssd1 vssd1 vccd1 vccd1 _11855_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_28_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10049__B1 _10915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10806_ _10806_/A _10806_/B vssd1 vssd1 vccd1 vccd1 _10808_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11786_ hold257/A _11786_/B vssd1 vssd1 vccd1 vccd1 _11786_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_82_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13525_ hold292/X _13555_/A2 _13524_/X _13542_/B2 vssd1 vssd1 vccd1 vccd1 hold293/A
+ sky130_fd_sc_hd__a22o_1
X_10737_ _10736_/A _10736_/B _10736_/Y _12047_/C1 vssd1 vssd1 vccd1 vccd1 _10737_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13520__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13538__B2 _13542_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13456_ _13456_/A _13456_/B vssd1 vssd1 vccd1 vccd1 _13456_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10668_ _10668_/A _10668_/B vssd1 vssd1 vccd1 vccd1 _10669_/B sky130_fd_sc_hd__xnor2_1
X_12407_ _12405_/X _12406_/Y _12971_/S _12404_/X vssd1 vssd1 vccd1 vccd1 dest_val[24]
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10599_ _10597_/X _10598_/X _11575_/S vssd1 vssd1 vccd1 vccd1 _10599_/X sky130_fd_sc_hd__mux2_1
X_13387_ _07235_/B _13419_/A2 hold77/X vssd1 vssd1 vccd1 vccd1 _13675_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_106_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12338_ _12668_/A _12338_/B vssd1 vssd1 vccd1 vccd1 _12348_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12269_ _12270_/A _12270_/B vssd1 vssd1 vccd1 vccd1 _12351_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09445__S _09674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10524__A1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10524__B2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06830_ reg1_val[25] _07252_/B vssd1 vssd1 vccd1 vccd1 _06831_/B sky130_fd_sc_hd__and2_1
X_06761_ reg1_val[31] vssd1 vssd1 vccd1 vccd1 _13135_/A sky130_fd_sc_hd__inv_6
XFILLER_0_78_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08500_ _08498_/A _08498_/B _08499_/Y vssd1 vssd1 vccd1 vccd1 _08510_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_78_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09480_ _09476_/X _09479_/X _10005_/S vssd1 vssd1 vccd1 vccd1 _10172_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_78_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08431_ _08821_/B2 fanout85/X fanout82/X _08821_/A1 vssd1 vssd1 vccd1 vccd1 _08432_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_53_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06817__B _13048_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08362_ _08365_/B _08361_/Y _08298_/X vssd1 vssd1 vccd1 vccd1 _08990_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_86_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07313_ _07300_/Y _10536_/A1 wire101/A _10536_/B2 vssd1 vssd1 vccd1 vccd1 _07314_/B
+ sky130_fd_sc_hd__a22o_1
X_08293_ _08293_/A _08367_/A vssd1 vssd1 vccd1 vccd1 _08302_/A sky130_fd_sc_hd__or2_1
XFILLER_0_46_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout136_A _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07244_ _08951_/A _07244_/B vssd1 vssd1 vccd1 vccd1 _07687_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13529__B2 _13542_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06833__A _06928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07175_ _10239_/A _10096_/A _07173_/Y vssd1 vssd1 vccd1 vccd1 _07175_/X sky130_fd_sc_hd__a21o_4
XANTENNA__10355__A _11076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09582__C _10787_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08184__A2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09816_ _09816_/A _09816_/B vssd1 vssd1 vccd1 vccd1 _09817_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_94_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09747_ _09747_/A _09747_/B vssd1 vssd1 vccd1 vccd1 _09789_/A sky130_fd_sc_hd__xnor2_1
X_06959_ _07093_/B vssd1 vssd1 vccd1 vccd1 _10992_/A sky130_fd_sc_hd__inv_2
XANTENNA__09133__A1 _07300_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09133__B2 wire101/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10818__A2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09678_ _09467_/X _09493_/X _09703_/B vssd1 vssd1 vccd1 vccd1 _09678_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_68_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _10944_/A _08640_/B vssd1 vssd1 vccd1 vccd1 _08629_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_68_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08892__B1 _09910_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _11640_/A _11640_/B vssd1 vssd1 vccd1 vccd1 _11642_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_126_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11571_ reg1_val[15] curr_PC[15] vssd1 vssd1 vccd1 vccd1 _11572_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_91_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13310_ _13569_/B _13570_/A _13218_/X vssd1 vssd1 vccd1 vccd1 _13574_/B sky130_fd_sc_hd__a21oi_1
X_10522_ _10522_/A _10522_/B vssd1 vssd1 vccd1 vccd1 _10523_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10453_ _09841_/X _09844_/X _10600_/S vssd1 vssd1 vccd1 vccd1 _10453_/X sky130_fd_sc_hd__mux2_1
X_13241_ hold259/X hold116/X vssd1 vssd1 vccd1 vccd1 _13535_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_32_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10384_ _10215_/A _10214_/Y _10213_/A vssd1 vssd1 vccd1 vccd1 _10395_/A sky130_fd_sc_hd__a21o_1
X_13172_ _13172_/A1 _13194_/A2 hold58/X _13543_/A vssd1 vssd1 vccd1 vccd1 _13622_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12123_ _12035_/B _12207_/A vssd1 vssd1 vccd1 vccd1 _12290_/A sky130_fd_sc_hd__nand2b_1
X_12054_ _13660_/Q _12148_/C vssd1 vssd1 vccd1 vccd1 _12056_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10506__A1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11703__B1 _12695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10506__B2 _12557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11005_ _11693_/A2 _11248_/C _13651_/Q vssd1 vssd1 vccd1 vccd1 _11005_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09124__A1 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09124__B2 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10150__D _10577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13515__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12956_ _12956_/A _12956_/B vssd1 vssd1 vccd1 vccd1 _12961_/D sky130_fd_sc_hd__xnor2_4
XFILLER_0_99_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11907_ _11907_/A _11907_/B vssd1 vssd1 vccd1 vccd1 _11925_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__11482__A2 _12754_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12887_ _12893_/B _12887_/B vssd1 vssd1 vccd1 vccd1 new_PC[12] sky130_fd_sc_hd__and2_4
XFILLER_0_68_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11838_ _11838_/A _11838_/B _11838_/C vssd1 vssd1 vccd1 vccd1 _11839_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_114_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08635__B1 _11047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11769_ _12742_/A _09048_/X _09049_/Y vssd1 vssd1 vccd1 vccd1 _11769_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13508_ _13255_/X _13508_/B vssd1 vssd1 vccd1 vccd1 _13509_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_83_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13439_ _07639_/B _13598_/C hold26/X vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__o21a_1
XFILLER_0_3_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08980_ _08980_/A _08980_/B vssd1 vssd1 vccd1 vccd1 _08980_/X sky130_fd_sc_hd__xor2_1
XANTENNA__10903__A _12551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07931_ _07502_/A _07501_/Y _07500_/A vssd1 vssd1 vccd1 vccd1 _07943_/A sky130_fd_sc_hd__a21bo_2
XFILLER_0_48_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07862_ _07862_/A _07862_/B vssd1 vssd1 vccd1 vccd1 _07863_/B sky130_fd_sc_hd__or2_1
XANTENNA__07634__D _07634_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07913__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09601_ _09753_/B _09600_/B _09600_/C vssd1 vssd1 vccd1 vccd1 _09602_/C sky130_fd_sc_hd__a21o_1
X_06813_ _06815_/A vssd1 vssd1 vccd1 vccd1 _06813_/Y sky130_fd_sc_hd__inv_2
X_07793_ _07796_/A _07796_/B vssd1 vssd1 vccd1 vccd1 _07793_/X sky130_fd_sc_hd__and2_1
XFILLER_0_3_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09532_ _10176_/A _09536_/B vssd1 vssd1 vccd1 vccd1 _10601_/C sky130_fd_sc_hd__or2_1
X_06744_ _13141_/A vssd1 vssd1 vccd1 vccd1 _06744_/Y sky130_fd_sc_hd__inv_2
X_09463_ reg1_val[8] reg1_val[23] _09463_/S vssd1 vssd1 vccd1 vccd1 _09463_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout253_A _13141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08414_ _08353_/A _08353_/C _08353_/B vssd1 vssd1 vccd1 vccd1 _08415_/B sky130_fd_sc_hd__o21ai_1
X_09394_ _12094_/A _09394_/B vssd1 vssd1 vccd1 vccd1 _09395_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08345_ _08345_/A _08345_/B vssd1 vssd1 vccd1 vccd1 _08355_/B sky130_fd_sc_hd__xor2_2
XANTENNA__08626__B1 _10225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08276_ _08951_/A _08276_/B vssd1 vssd1 vccd1 vccd1 _08278_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07227_ _07245_/A _07245_/B vssd1 vssd1 vccd1 vccd1 _07227_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_6_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07158_ _12982_/A _09694_/A reg1_val[2] reg1_val[3] vssd1 vssd1 vccd1 vccd1 _07265_/D
+ sky130_fd_sc_hd__or4_2
XFILLER_0_42_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11909__A _12093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07089_ _09501_/A _09703_/B vssd1 vssd1 vccd1 vccd1 _09659_/A sky130_fd_sc_hd__nand2_2
Xfanout120 _07456_/Y vssd1 vssd1 vccd1 vccd1 _10915_/A sky130_fd_sc_hd__buf_4
Xfanout131 _07285_/Y vssd1 vssd1 vccd1 vccd1 _10235_/B2 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09354__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout142 _12735_/A1 vssd1 vssd1 vccd1 vccd1 _12374_/A sky130_fd_sc_hd__buf_4
XANTENNA__09354__B2 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13150__A2 _13193_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout164 _13193_/B vssd1 vssd1 vccd1 vccd1 _13191_/B sky130_fd_sc_hd__clkbuf_4
Xfanout175 _07267_/X vssd1 vssd1 vccd1 vccd1 _10236_/A sky130_fd_sc_hd__clkbuf_16
Xfanout186 _13550_/A2 vssd1 vssd1 vccd1 vccd1 _13555_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout197 _07210_/Y vssd1 vssd1 vccd1 vccd1 _09659_/B sky130_fd_sc_hd__clkbuf_16
XANTENNA__13438__B1 _13444_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09106__A1 _07347_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09106__B2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12810_ _12816_/B _12810_/B vssd1 vssd1 vccd1 vccd1 new_PC[1] sky130_fd_sc_hd__and2_4
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _12740_/A _12739_/B _12739_/Y _09506_/X vssd1 vssd1 vccd1 vccd1 _12741_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ _12671_/B _12671_/C _12671_/A vssd1 vssd1 vccd1 vccd1 _12673_/B sky130_fd_sc_hd__a21oi_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _11997_/A _07643_/B fanout13/X _11922_/A vssd1 vssd1 vccd1 vccd1 _11624_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07569__A _11508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11554_ _11554_/A _11663_/A vssd1 vssd1 vccd1 vccd1 _11763_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_108_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10505_ _11709_/A _10505_/B vssd1 vssd1 vccd1 vccd1 _10508_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11485_ _12537_/B2 _11473_/X _11484_/X _12710_/B2 _11483_/X vssd1 vssd1 vccd1 vccd1
+ _11485_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_107_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13224_ hold269/X hold39/X vssd1 vssd1 vccd1 vccd1 _13225_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10436_ _10146_/X _10294_/X _10295_/X vssd1 vssd1 vccd1 vccd1 _10438_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_0_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09593__A1 _11732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09593__B2 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13155_ hold78/X _13191_/B vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__or2_1
X_10367_ _07275_/Y fanout6/X _10366_/X _10236_/A vssd1 vssd1 vccd1 vccd1 _10369_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06920__B _06920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06946__A3 _13042_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12106_ _12107_/A _12107_/B vssd1 vssd1 vccd1 vccd1 _12192_/B sky130_fd_sc_hd__nor2_1
X_13086_ reg1_val[21] _13129_/B vssd1 vssd1 vccd1 vccd1 _13086_/Y sky130_fd_sc_hd__nor2_1
X_10298_ _10298_/A _10433_/A _10577_/A _10631_/A vssd1 vssd1 vccd1 vccd1 _10298_/X
+ sky130_fd_sc_hd__or4_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12037_ _12037_/A _12037_/B vssd1 vssd1 vccd1 vccd1 _12037_/X sky130_fd_sc_hd__and2_1
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11554__A _11554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12939_ _12961_/A _12963_/A vssd1 vssd1 vccd1 vccd1 _12941_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_87_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12404__A1 _10730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08130_ _08130_/A _08174_/A vssd1 vssd1 vccd1 vccd1 _08224_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_56_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09281__B1 _08246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08061_ _12982_/A _07203_/Y _08271_/A _07198_/Y vssd1 vssd1 vccd1 vccd1 _08062_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07831__A1 fanout39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07831__B2 _08118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07012_ _06928_/A _06936_/B _12995_/B _07011_/X vssd1 vssd1 vccd1 vccd1 _09496_/S
+ sky130_fd_sc_hd__a31oi_4
XFILLER_0_114_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09694__A _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08387__A2 _07541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11729__A _11802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08963_ _08947_/B _09010_/B _08945_/Y vssd1 vssd1 vccd1 vccd1 _09012_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07914_ _12092_/A _07914_/B vssd1 vssd1 vccd1 vccd1 _07915_/A sky130_fd_sc_hd__xnor2_1
X_08894_ _08902_/B _08902_/A vssd1 vssd1 vccd1 vccd1 _08896_/C sky130_fd_sc_hd__and2b_1
X_07845_ _07845_/A _07845_/B vssd1 vssd1 vccd1 vccd1 _08036_/B sky130_fd_sc_hd__xor2_1
X_07776_ _07776_/A _07776_/B vssd1 vssd1 vccd1 vccd1 _07841_/B sky130_fd_sc_hd__xnor2_2
X_09515_ _09516_/A _09516_/B vssd1 vssd1 vccd1 vccd1 _09515_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_94_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09446_ reg1_val[5] reg1_val[26] _09463_/S vssd1 vssd1 vccd1 vccd1 _09446_/X sky130_fd_sc_hd__mux2_1
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08773__A _10236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09377_ _09377_/A _09377_/B vssd1 vssd1 vccd1 vccd1 _09379_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_47_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08328_ _07219_/Y _11732_/A _10814_/A1 _08328_/B2 vssd1 vssd1 vccd1 vccd1 _08329_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09272__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08259_ _08257_/A _08257_/B _08257_/C vssd1 vssd1 vccd1 vccd1 _08260_/C sky130_fd_sc_hd__a21oi_2
XFILLER_0_62_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11270_ _11823_/A _11270_/B vssd1 vssd1 vccd1 vccd1 _11274_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10221_ _10222_/A _10222_/B _10098_/Y vssd1 vssd1 vccd1 vccd1 _10221_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_120_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10185__A2 _12793_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10152_ _09823_/X _09983_/X _09984_/X vssd1 vssd1 vccd1 vccd1 _10152_/X sky130_fd_sc_hd__a21o_1
XANTENNA__08013__A _10266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10083_ fanout42/X fanout25/X fanout23/X fanout40/X vssd1 vssd1 vccd1 vccd1 _10084_/B
+ sky130_fd_sc_hd__o22a_1
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12189__B _12764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10985_ _11864_/A _10900_/Y _10984_/X vssd1 vssd1 vccd1 vccd1 _10985_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_85_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12724_ _12724_/A _12724_/B _12724_/C vssd1 vssd1 vccd1 vccd1 _12727_/A sky130_fd_sc_hd__nor3_1
XANTENNA__08683__A _10236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12655_ hold247/A _12786_/B1 _12702_/B _12654_/Y _12748_/B1 vssd1 vssd1 vccd1 vccd1
+ _12661_/B sky130_fd_sc_hd__a311o_1
XFILLER_0_127_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07299__A _11793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11606_ _11607_/A _11607_/B vssd1 vssd1 vccd1 vccd1 _11714_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12586_ reg1_val[27] curr_PC[27] vssd1 vssd1 vccd1 vccd1 _12586_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_108_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11537_ _11538_/A _11538_/B _11536_/Y vssd1 vssd1 vccd1 vccd1 _11537_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_52_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11468_ reg1_val[14] curr_PC[14] vssd1 vssd1 vccd1 vccd1 _11469_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_123_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13207_ hold172/X _13207_/B vssd1 vssd1 vccd1 vccd1 hold173/A sky130_fd_sc_hd__or2_1
X_10419_ _10261_/Y _10275_/B _10273_/Y vssd1 vssd1 vccd1 vccd1 _10421_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__13362__A2 _13542_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11399_ _11400_/A _11400_/B vssd1 vssd1 vccd1 vccd1 _11399_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_110_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07238__S _08951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11268__B _11600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13138_ hold143/X hold15/X _13597_/B vssd1 vssd1 vccd1 vccd1 hold192/A sky130_fd_sc_hd__nand3_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _13065_/B _13081_/A vssd1 vssd1 vccd1 vccd1 _13071_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_31_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10900__B _10900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07630_ _07630_/A _07630_/B vssd1 vssd1 vccd1 vccd1 _07631_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_88_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07561_ _10049_/A2 _08395_/B _09885_/B1 fanout28/X vssd1 vssd1 vccd1 vccd1 _07562_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_88_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09300_ _09169_/A _09169_/B _09167_/X vssd1 vssd1 vccd1 vccd1 _09303_/A sky130_fd_sc_hd__a21o_2
X_07492_ _07492_/A _07492_/B vssd1 vssd1 vccd1 vccd1 _07492_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_61_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09231_ _07203_/Y _10536_/A1 _10536_/B2 _07230_/Y vssd1 vssd1 vccd1 vccd1 _09232_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06825__B _12981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09162_ _09910_/A1 _07643_/B fanout13/X _09604_/A vssd1 vssd1 vccd1 vccd1 _09163_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08113_ _08113_/A _08113_/B vssd1 vssd1 vccd1 vccd1 _08116_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07804__A1 _10235_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07804__B2 _10235_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09093_ _09086_/B _09086_/C _09092_/A _09318_/B vssd1 vssd1 vccd1 vccd1 _09094_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_44_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08044_ _08044_/A _08044_/B vssd1 vssd1 vccd1 vccd1 _08155_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07568__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09995_ _12130_/A _09994_/B _09994_/C vssd1 vssd1 vccd1 vccd1 _09996_/B sky130_fd_sc_hd__a21oi_1
X_08946_ _08946_/A _08946_/B vssd1 vssd1 vccd1 vccd1 _08947_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08768__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08877_ _08877_/A _08889_/A vssd1 vssd1 vccd1 vccd1 _08898_/A sky130_fd_sc_hd__nand2_2
XANTENNA__10810__B _11802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07828_ _07828_/A _07828_/B vssd1 vssd1 vccd1 vccd1 _07996_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_79_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11419__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07759_ _07772_/B _07815_/A _07772_/A vssd1 vssd1 vccd1 vccd1 _07774_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11922__A _11922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09493__A0 _13015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10770_ _11708_/A _10770_/B vssd1 vssd1 vccd1 vccd1 _10778_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout31_A _07421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09429_ _09524_/A _13748_/A instruction[5] _13744_/A vssd1 vssd1 vccd1 vccd1 _09429_/X
+ sky130_fd_sc_hd__or4b_4
XFILLER_0_82_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10538__A _10538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08048__A1 _11047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12440_ _12440_/A _12440_/B _12440_/C vssd1 vssd1 vccd1 vccd1 _12682_/B sky130_fd_sc_hd__and3_1
XANTENNA__08048__B2 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11052__B1 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12371_ _12508_/A _12371_/B vssd1 vssd1 vccd1 vccd1 _12480_/A sky130_fd_sc_hd__xor2_4
XANTENNA__08950__B _08950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11322_ _11204_/A _11204_/B _11203_/A vssd1 vssd1 vccd1 vccd1 _11332_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09548__A1 _07699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09548__B2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13344__A2 _13506_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11253_ _11252_/B _11369_/B hold271/A vssd1 vssd1 vccd1 vccd1 _11253_/X sky130_fd_sc_hd__a21o_1
X_10204_ _10100_/A _10100_/B _10103_/A vssd1 vssd1 vccd1 vccd1 _10219_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__07023__A2 _07025_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11184_ _11185_/A _11184_/B vssd1 vssd1 vccd1 vccd1 _11315_/B sky130_fd_sc_hd__nand2_1
X_10135_ _09923_/A _09923_/B _09964_/B _09962_/Y vssd1 vssd1 vccd1 vccd1 _10137_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_100_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07582__A _11286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10066_ _09935_/A _09934_/B _09934_/A vssd1 vssd1 vccd1 vccd1 _10068_/B sky130_fd_sc_hd__o21bai_2
XFILLER_0_89_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10330__A2 _11587_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12607__A1 _12666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10968_ _10968_/A _10968_/B vssd1 vssd1 vccd1 vccd1 _10970_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10094__A1 _10235_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12707_ hold197/A _12374_/A _12750_/B _12795_/A1 vssd1 vssd1 vccd1 vccd1 _12707_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_57_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10094__B2 _10235_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13687_ _13701_/CLK _13687_/D vssd1 vssd1 vccd1 vccd1 hold132/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10899_ _10342_/A _10766_/Y _10898_/X vssd1 vssd1 vccd1 vccd1 dest_val[9] sky130_fd_sc_hd__a21oi_4
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12638_ _12633_/Y _12636_/X _12637_/Y vssd1 vssd1 vccd1 vccd1 _12638_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11043__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12569_ _12567_/X _12569_/B vssd1 vssd1 vccd1 vccd1 _12681_/A sky130_fd_sc_hd__nand2b_2
XANTENNA__07179__D _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11594__A1 _09529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09448__S _09674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12791__B1 _09519_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold206 hold206/A vssd1 vssd1 vccd1 vccd1 hold206/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 hold217/A vssd1 vssd1 vccd1 vccd1 hold217/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 hold228/A vssd1 vssd1 vccd1 vccd1 hold228/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07476__B _07476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold239 hold239/A vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _08950_/B _10522_/A _08868_/B1 _08866_/B2 vssd1 vssd1 vccd1 vccd1 _08801_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _09949_/A _09780_/B vssd1 vssd1 vccd1 vccd1 _09783_/A sky130_fd_sc_hd__xnor2_4
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06992_ reg1_val[5] _07180_/C vssd1 vssd1 vccd1 vccd1 _10447_/B sky130_fd_sc_hd__nand2_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07492__A _07492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ _08758_/A _08758_/B vssd1 vssd1 vccd1 vccd1 _08731_/X sky130_fd_sc_hd__and2_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09711__A1 _09507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08662_ _08662_/A _08662_/B vssd1 vssd1 vccd1 vccd1 _08690_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__10321__A2 _12760_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07613_ fanout56/X _10235_/A1 _10235_/B2 fanout53/X vssd1 vssd1 vccd1 vccd1 _07614_/B
+ sky130_fd_sc_hd__o22a_1
X_08593_ _08923_/B1 _10538_/A _08778_/B _08866_/A2 vssd1 vssd1 vccd1 vccd1 _08594_/B
+ sky130_fd_sc_hd__o22a_1
X_07544_ _07544_/A _07544_/B vssd1 vssd1 vccd1 vccd1 _07544_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_49_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12557__B _12557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07475_ _07476_/B _07476_/C _07476_/A vssd1 vssd1 vccd1 vccd1 _07478_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_91_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09214_ _08118_/B _07451_/X _09885_/B1 fanout39/X vssd1 vssd1 vccd1 vccd1 _09215_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_119_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09145_ _09254_/A _09146_/B vssd1 vssd1 vccd1 vccd1 _09145_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_44_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07789__B1 _08580_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09076_ _08361_/Y _08413_/X _08363_/Y vssd1 vssd1 vccd1 vccd1 _09080_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_31_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08027_ _08027_/A _08027_/B vssd1 vssd1 vccd1 vccd1 _08028_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_4_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13326__A2 _13463_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11189__A _11825_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07005__A2 _06936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08202__A1 _07237_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09978_ _09979_/B _09979_/A vssd1 vssd1 vccd1 vccd1 _09978_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout79_A _08580_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08929_ _08916_/X _08929_/B _08938_/A vssd1 vssd1 vccd1 vccd1 _08929_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_98_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09702__A1 _12515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11940_ _11940_/A _11940_/B vssd1 vssd1 vccd1 vccd1 _11942_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_99_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11871_ _07092_/B _11869_/X _11870_/Y vssd1 vssd1 vccd1 vccd1 _11871_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_67_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13610_ _13708_/CLK hold12/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dfxtp_1
X_10822_ _10823_/A _10823_/B vssd1 vssd1 vccd1 vccd1 _10937_/B sky130_fd_sc_hd__or2_1
XANTENNA__11912__A_N _11913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13541_ hold261/X _13540_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13541_/X sky130_fd_sc_hd__mux2_1
X_10753_ _12058_/A _10885_/B hold295/A vssd1 vssd1 vccd1 vccd1 _10753_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__10268__A _11709_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13472_ _13547_/A _13472_/B vssd1 vssd1 vccd1 vccd1 _13710_/D sky130_fd_sc_hd__and2_1
X_10684_ _10684_/A _10684_/B vssd1 vssd1 vccd1 vccd1 _10685_/B sky130_fd_sc_hd__or2_1
XFILLER_0_82_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09769__A1 _11732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12423_ _12423_/A _12423_/B vssd1 vssd1 vccd1 vccd1 _12424_/B sky130_fd_sc_hd__or2_1
XANTENNA__09769__B2 _10814_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12354_ _12355_/A _12355_/B vssd1 vssd1 vccd1 vccd1 _12437_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06988__D1 _06936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11305_ _11825_/A _11305_/B vssd1 vssd1 vccd1 vccd1 _11307_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12285_ _12286_/A _12286_/B _12286_/C vssd1 vssd1 vccd1 vccd1 _12288_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09792__A _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11236_ _11463_/A _06947_/Y _07041_/X _11235_/Y vssd1 vssd1 vccd1 vccd1 _11237_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09941__A1 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11827__A _12417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09941__B2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11167_ _12417_/A _11167_/B vssd1 vssd1 vccd1 vccd1 _11171_/A sky130_fd_sc_hd__xnor2_1
X_10118_ fanout39/X fanout82/X _11423_/A _08118_/B vssd1 vssd1 vccd1 vccd1 _10119_/B
+ sky130_fd_sc_hd__o22a_1
X_11098_ _11099_/A _11099_/B vssd1 vssd1 vccd1 vccd1 _11222_/A sky130_fd_sc_hd__nand2_1
X_10049_ fanout35/X _10049_/A2 _10915_/A _07699_/B vssd1 vssd1 vccd1 vccd1 _10050_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11500__A1 _11922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11500__B2 wire101/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13739_ _13739_/CLK hold171/X vssd1 vssd1 vccd1 vccd1 hold169/A sky130_fd_sc_hd__dfxtp_1
X_07260_ _07261_/A _07261_/B vssd1 vssd1 vccd1 vccd1 _07644_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08680__A1 _08806_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08871__A _09948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08680__B2 _08806_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07191_ _07281_/A _07309_/A _11793_/A _07297_/A vssd1 vssd1 vccd1 vccd1 _07192_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_0_60_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07487__A _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09901_ _10266_/A _09901_/B vssd1 vssd1 vccd1 vccd1 _09909_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09832_ _09723_/Y _10726_/B _09831_/X vssd1 vssd1 vccd1 vccd1 _09832_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_6_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _09763_/A _09763_/B vssd1 vssd1 vccd1 vccd1 _09765_/B sky130_fd_sc_hd__xnor2_1
X_06975_ _06928_/A _06928_/B _13020_/B _06974_/X vssd1 vssd1 vccd1 vccd1 _07492_/A
+ sky130_fd_sc_hd__a31o_4
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08714_ _08714_/A _08714_/B vssd1 vssd1 vccd1 vccd1 _08761_/A sky130_fd_sc_hd__xnor2_1
X_09694_ _09694_/A curr_PC[1] vssd1 vssd1 vccd1 vccd1 _09695_/B sky130_fd_sc_hd__or2_1
X_08645_ _08645_/A _08645_/B vssd1 vssd1 vccd1 vccd1 _08646_/B sky130_fd_sc_hd__nor2_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08576_ _08576_/A _08576_/B vssd1 vssd1 vccd1 vccd1 _08615_/B sky130_fd_sc_hd__xnor2_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07527_ _07527_/A _07527_/B vssd1 vssd1 vccd1 vccd1 _07527_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07458_ _10263_/A _07458_/B vssd1 vssd1 vccd1 vccd1 _07502_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07389_ _07395_/A _07395_/B vssd1 vssd1 vccd1 vccd1 _12420_/A sky130_fd_sc_hd__nand2_4
XANTENNA__12755__B1 _09519_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09128_ _09129_/A _09129_/B vssd1 vssd1 vccd1 vccd1 _09128_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09620__B1 _07471_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10230__A1 _10374_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09059_ _09055_/B _09055_/C _09057_/A _09055_/A vssd1 vssd1 vccd1 vccd1 _09060_/C
+ sky130_fd_sc_hd__a211o_1
XANTENNA__10230__B2 _10349_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12070_ curr_PC[19] curr_PC[20] _12070_/C vssd1 vssd1 vccd1 vccd1 _12160_/B sky130_fd_sc_hd__and3_1
XFILLER_0_102_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11021_ _12825_/S _11265_/C vssd1 vssd1 vccd1 vccd1 _11021_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07934__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11730__A1 _07198_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11730__B2 _11997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12972_ _12979_/A _12973_/B vssd1 vssd1 vccd1 vccd1 _12974_/A sky130_fd_sc_hd__and2_1
XANTENNA__07860__A _09940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11923_ _11923_/A _11923_/B vssd1 vssd1 vccd1 vccd1 _11924_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_99_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07162__A1 _07535_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11854_ _11852_/Y _11854_/B vssd1 vssd1 vccd1 vccd1 _12035_/A sky130_fd_sc_hd__nand2b_4
XFILLER_0_79_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10049__A1 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10049__B2 _07699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10805_ _11719_/A _10805_/B vssd1 vssd1 vccd1 vccd1 _10806_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11785_ hold292/A hold296/A _11881_/D _12058_/A vssd1 vssd1 vccd1 vccd1 _11786_/B
+ sky130_fd_sc_hd__o31a_1
X_13524_ hold296/A _13523_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13524_/X sky130_fd_sc_hd__mux2_1
X_10736_ _10736_/A _10736_/B vssd1 vssd1 vccd1 vccd1 _10736_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_36_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13455_ _13279_/X _13455_/B vssd1 vssd1 vccd1 vccd1 _13456_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__13538__A2 _13555_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10667_ _10668_/A _10668_/B vssd1 vssd1 vccd1 vccd1 _10667_/X sky130_fd_sc_hd__or2_1
XFILLER_0_125_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12406_ curr_PC[24] _12477_/C _12406_/B1 vssd1 vssd1 vccd1 vccd1 _12406_/Y sky130_fd_sc_hd__o21ai_1
X_13386_ hold1/X _13416_/A2 _13444_/B1 hold76/X _13383_/A vssd1 vssd1 vccd1 vccd1
+ hold77/A sky130_fd_sc_hd__o221a_1
X_10598_ _10000_/X _10005_/X _10600_/S vssd1 vssd1 vccd1 vccd1 _10598_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12337_ _12614_/A fanout16/X fanout12/X _07257_/X vssd1 vssd1 vccd1 vccd1 _12338_/B
+ sky130_fd_sc_hd__a22o_1
X_12268_ _12268_/A _12666_/A vssd1 vssd1 vccd1 vccd1 _12270_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_121_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11219_ _11219_/A _11219_/B vssd1 vssd1 vccd1 vccd1 _11220_/B sky130_fd_sc_hd__or2_1
X_12199_ _12200_/B _12200_/A vssd1 vssd1 vccd1 vccd1 _12286_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__10524__A2 _07478_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06760_ reg1_val[28] vssd1 vssd1 vccd1 vccd1 _12647_/A sky130_fd_sc_hd__inv_2
XANTENNA__09461__S _09674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09142__A2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08430_ _08857_/A _08430_/B vssd1 vssd1 vccd1 vccd1 _08436_/A sky130_fd_sc_hd__xor2_1
X_08361_ _08364_/A _08364_/B vssd1 vssd1 vccd1 vccd1 _08361_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_86_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07312_ _10649_/A _07312_/B vssd1 vssd1 vccd1 vccd1 _08833_/B sky130_fd_sc_hd__or2_2
XFILLER_0_46_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09697__A _12525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08292_ _08293_/A _08292_/B _08292_/C vssd1 vssd1 vccd1 vccd1 _08367_/A sky130_fd_sc_hd__nor3_1
XANTENNA__09385__A_N _09386_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07243_ fanout47/X _08866_/B2 _08950_/B fanout45/X vssd1 vssd1 vccd1 vccd1 _07244_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_73_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13529__A2 _13555_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10636__A _11825_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06833__B _13036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07174_ _10239_/A _10096_/A _07173_/Y vssd1 vssd1 vccd1 vccd1 _09582_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_103_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11960__A1 _12515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07916__B1 _08923_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ _09815_/A _09815_/B vssd1 vssd1 vccd1 vccd1 _09816_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09746_ _09747_/A _09747_/B vssd1 vssd1 vccd1 vccd1 _09896_/B sky130_fd_sc_hd__nand2_1
X_06958_ _06956_/Y _06958_/B vssd1 vssd1 vccd1 vccd1 _07093_/B sky130_fd_sc_hd__nand2b_2
XANTENNA__09133__A2 _07541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _09669_/X _09676_/X _11575_/S vssd1 vssd1 vccd1 vccd1 _09677_/X sky130_fd_sc_hd__mux2_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06889_ reg1_val[18] _07309_/A vssd1 vssd1 vccd1 vccd1 _11958_/B sky130_fd_sc_hd__nand2_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08628_ _08685_/A _08685_/B vssd1 vssd1 vccd1 vccd1 _08640_/B sky130_fd_sc_hd__nand2_2
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08892__A1 _07175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08892__B2 _08933_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08559_ _08559_/A _08621_/A vssd1 vssd1 vccd1 vccd1 _08576_/A sky130_fd_sc_hd__nand2_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11570_ reg1_val[15] curr_PC[15] vssd1 vssd1 vccd1 vccd1 _11572_/A sky130_fd_sc_hd__or2_1
XFILLER_0_64_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10521_ _10521_/A _10521_/B vssd1 vssd1 vccd1 vccd1 _10523_/A sky130_fd_sc_hd__nor2_1
XANTENNA_fanout8_A fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13240_ hold116/X hold259/X vssd1 vssd1 vccd1 vccd1 _13240_/X sky130_fd_sc_hd__and2b_1
X_10452_ _11576_/A _10451_/A _09535_/Y vssd1 vssd1 vccd1 vccd1 _12462_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_122_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13171_ hold57/X _13191_/B vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__or2_1
XFILLER_0_20_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10383_ _10383_/A _10383_/B vssd1 vssd1 vccd1 vccd1 _10397_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_60_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12122_ _11943_/Y _12031_/X _12033_/B vssd1 vssd1 vccd1 vccd1 _12122_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12053_ _11143_/X _12052_/X _12525_/A vssd1 vssd1 vccd1 vccd1 _12053_/X sky130_fd_sc_hd__mux2_1
X_11004_ hold240/A _11004_/B vssd1 vssd1 vccd1 vccd1 _11248_/C sky130_fd_sc_hd__or2_1
XANTENNA__09372__A2 _10787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07590__A _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09124__A2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12955_ reg1_val[23] curr_PC[23] _12978_/S vssd1 vssd1 vccd1 vccd1 _12956_/B sky130_fd_sc_hd__mux2_2
X_11906_ _11906_/A _11906_/B vssd1 vssd1 vccd1 vccd1 _11907_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13208__A1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12886_ _12886_/A _12886_/B _12886_/C vssd1 vssd1 vccd1 vccd1 _12887_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_68_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11837_ _11838_/A _11838_/B _11838_/C vssd1 vssd1 vccd1 vccd1 _11935_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_55_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08635__A1 _08866_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _11703_/X _12163_/B _11767_/Y vssd1 vssd1 vccd1 vccd1 _11768_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__08635__B2 _08950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10719_ _10719_/A _10719_/B _10719_/C vssd1 vssd1 vccd1 vccd1 _10720_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_70_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13507_ _13543_/A hold272/X vssd1 vssd1 vccd1 vccd1 _13717_/D sky130_fd_sc_hd__and2_1
XFILLER_0_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11699_ _07297_/A _11793_/B _07152_/X _11698_/X vssd1 vssd1 vccd1 vccd1 _11699_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_82_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13438_ hold25/X _13142_/A _13444_/B1 hold81/A _13568_/A vssd1 vssd1 vccd1 vccd1
+ hold26/A sky130_fd_sc_hd__o221a_1
XFILLER_0_3_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13369_ _13547_/A hold217/X vssd1 vssd1 vccd1 vccd1 _13666_/D sky130_fd_sc_hd__and2_1
XFILLER_0_23_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07765__A _10119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07930_ _07930_/A _07930_/B vssd1 vssd1 vccd1 vccd1 _07944_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_48_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07861_ _07862_/A _07862_/B vssd1 vssd1 vccd1 vccd1 _07861_/X sky130_fd_sc_hd__and2_1
XFILLER_0_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09600_ _09753_/B _09600_/B _09600_/C vssd1 vssd1 vccd1 vccd1 _09726_/A sky130_fd_sc_hd__nand3_2
X_06812_ reg1_val[29] _09254_/B vssd1 vssd1 vccd1 vccd1 _06815_/A sky130_fd_sc_hd__nor2_1
X_07792_ _09575_/A _07792_/B vssd1 vssd1 vccd1 vccd1 _07796_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08596__A _10236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09531_ _10007_/S _09536_/B _09530_/X vssd1 vssd1 vccd1 vccd1 _10601_/B sky130_fd_sc_hd__o21a_1
X_06743_ hold161/X vssd1 vssd1 vccd1 vccd1 _06743_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12655__C1 _12748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09462_ reg1_val[9] reg1_val[22] _09463_/S vssd1 vssd1 vccd1 vccd1 _09462_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08413_ _08471_/A _08471_/B vssd1 vssd1 vccd1 vccd1 _08413_/X sky130_fd_sc_hd__or2_1
X_09393_ _07471_/Y fanout21/X _08246_/B fanout85/X vssd1 vssd1 vccd1 vccd1 _09394_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout246_A _06928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08344_ _08371_/A _08371_/B _08325_/Y vssd1 vssd1 vccd1 vccd1 _08355_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_46_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08626__A1 _08806_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08626__B2 _08806_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08275_ _07239_/Y _07300_/Y _11638_/A _07238_/X vssd1 vssd1 vccd1 vccd1 _08276_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07226_ _09950_/A _07226_/B vssd1 vssd1 vccd1 vccd1 _07245_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07378__C _07634_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13717_/CLK sky130_fd_sc_hd__clkbuf_8
X_07157_ _12982_/A _09694_/A reg1_val[2] vssd1 vssd1 vccd1 vccd1 _09871_/A sky130_fd_sc_hd__or3_2
XFILLER_0_30_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07088_ instruction[3] _13748_/A vssd1 vssd1 vccd1 vccd1 _09525_/C sky130_fd_sc_hd__nor2_2
XFILLER_0_112_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout110 _07495_/X vssd1 vssd1 vccd1 vccd1 _09885_/B1 sky130_fd_sc_hd__buf_6
XFILLER_0_10_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout132 _07237_/Y vssd1 vssd1 vccd1 vccd1 _08866_/B2 sky130_fd_sc_hd__clkbuf_8
XANTENNA__09354__A2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout143 _11231_/A vssd1 vssd1 vccd1 vccd1 _12735_/A1 sky130_fd_sc_hd__buf_2
Xfanout154 _08857_/A vssd1 vssd1 vccd1 vccd1 _10078_/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__07365__A1 _07476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout165 _13207_/B vssd1 vssd1 vccd1 vccd1 _13193_/B sky130_fd_sc_hd__buf_4
Xfanout187 _07118_/B vssd1 vssd1 vccd1 vccd1 _13550_/A2 sky130_fd_sc_hd__buf_2
Xfanout198 _07210_/Y vssd1 vssd1 vccd1 vccd1 _09949_/A sky130_fd_sc_hd__buf_8
XANTENNA_fanout61_A _10518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09106__A2 _07699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09729_ _10349_/A1 _07643_/B fanout13/X _10225_/A vssd1 vssd1 vccd1 vccd1 _09730_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12740_ _12740_/A _12740_/B vssd1 vssd1 vccd1 vccd1 _12740_/Y sky130_fd_sc_hd__nand2_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _12671_/A _12671_/B _12671_/C vssd1 vssd1 vccd1 vccd1 _12724_/A sky130_fd_sc_hd__and3_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11622_ _11622_/A vssd1 vssd1 vccd1 vccd1 _11631_/A sky130_fd_sc_hd__inv_2
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11553_ _11341_/A _11450_/A _11450_/B vssd1 vssd1 vccd1 vccd1 _11553_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10504_ fanout54/X fanout25/X fanout23/X _12268_/A vssd1 vssd1 vccd1 vccd1 _10505_/B
+ sky130_fd_sc_hd__o22a_1
X_11484_ _10458_/S _09691_/X _09537_/B vssd1 vssd1 vccd1 vccd1 _11484_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13374__B1 _13584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13223_ hold39/X hold269/X vssd1 vssd1 vccd1 vccd1 _13225_/A sky130_fd_sc_hd__and2b_1
X_10435_ _10435_/A _10435_/B _10435_/C vssd1 vssd1 vccd1 vccd1 _10435_/X sky130_fd_sc_hd__or3_1
XANTENNA__10188__B1 _12748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09593__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13154_ _10104_/A _13194_/A2 hold84/X _13547_/A vssd1 vssd1 vccd1 vccd1 _13613_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10366_ _10366_/A fanout5/X vssd1 vssd1 vccd1 vccd1 _10366_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ _12105_/A _12105_/B vssd1 vssd1 vccd1 vccd1 _12107_/B sky130_fd_sc_hd__xnor2_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ _13085_/A _13085_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[20] sky130_fd_sc_hd__nor2_8
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10297_ _10577_/A _10631_/A vssd1 vssd1 vccd1 vccd1 _10297_/X sky130_fd_sc_hd__or2_1
X_12036_ _11855_/X _12037_/B _12207_/B vssd1 vssd1 vccd1 vccd1 _12369_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_18_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13429__A1 _12253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12938_ _12938_/A _12938_/B _12938_/C vssd1 vssd1 vccd1 vccd1 _12963_/A sky130_fd_sc_hd__and3_1
XFILLER_0_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12869_ _13029_/B _12869_/B vssd1 vssd1 vccd1 vccd1 _12870_/B sky130_fd_sc_hd__or2_1
XANTENNA__12666__A _12666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13601__A1 _13207_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11612__B1 _09146_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09281__A1 _10915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09281__B2 _11047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08060_ _10239_/A _08060_/B vssd1 vssd1 vccd1 vccd1 _08064_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07831__A2 _08873_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07011_ reg2_val[2] _07110_/A vssd1 vssd1 vccd1 vccd1 _07011_/X sky130_fd_sc_hd__and2_1
XANTENNA__13497__A _13543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11376__C1 _11375_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08962_ _09005_/A _09008_/A _08961_/Y _08960_/B vssd1 vssd1 vccd1 vccd1 _09010_/B
+ sky130_fd_sc_hd__a22o_1
X_07913_ _10104_/A fanout14/X _07833_/B _10225_/A vssd1 vssd1 vccd1 vccd1 _07914_/B
+ sky130_fd_sc_hd__a22o_1
X_08893_ _09948_/A _08893_/B vssd1 vssd1 vccd1 vccd1 _08902_/B sky130_fd_sc_hd__xnor2_1
X_07844_ _07844_/A _07844_/B vssd1 vssd1 vccd1 vccd1 _08036_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09215__A _10119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07775_ _07845_/A _07773_/Y _07774_/A vssd1 vssd1 vccd1 vccd1 _07841_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_78_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09514_ _09525_/C _09514_/B vssd1 vssd1 vccd1 vccd1 _10866_/B sky130_fd_sc_hd__nand2_8
XFILLER_0_78_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09445_ _09443_/X _09444_/X _09674_/S vssd1 vssd1 vccd1 vccd1 _09445_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09376_ _09376_/A _09376_/B vssd1 vssd1 vccd1 vccd1 _09377_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08327_ _09373_/A _08327_/B vssd1 vssd1 vccd1 vccd1 _08333_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09272__A1 _09955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09272__B2 _09910_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08258_ _08258_/A _08258_/B vssd1 vssd1 vccd1 vccd1 _08260_/B sky130_fd_sc_hd__xor2_2
XANTENNA__12159__A1 _07201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07209_ _09694_/A _07572_/S _07208_/X vssd1 vssd1 vccd1 vccd1 _09779_/A sky130_fd_sc_hd__o21a_2
XANTENNA__13356__B1 _13506_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08189_ _08220_/A _08220_/B vssd1 vssd1 vccd1 vccd1 _08189_/X sky130_fd_sc_hd__and2_1
XANTENNA__12515__S _12515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10220_ _10082_/A _10082_/B _10081_/A vssd1 vssd1 vccd1 vccd1 _10224_/A sky130_fd_sc_hd__o21ai_4
X_10151_ _09325_/A _09325_/B _10150_/X vssd1 vssd1 vccd1 vccd1 _10155_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_100_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10082_ _10082_/A _10082_/B vssd1 vssd1 vccd1 vccd1 _10102_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__06749__A _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09125__A _09575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10984_ _11225_/A _10984_/B vssd1 vssd1 vccd1 vccd1 _10984_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_97_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12723_ _12723_/A _12723_/B vssd1 vssd1 vccd1 vccd1 _12724_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12654_ _12786_/B1 _12702_/B hold247/A vssd1 vssd1 vccd1 vccd1 _12654_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11605_ _12094_/A _11605_/B vssd1 vssd1 vccd1 vccd1 _11607_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12585_ _12524_/A _12521_/Y _12523_/B vssd1 vssd1 vccd1 vccd1 _12589_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_53_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11536_ _11424_/A _11424_/B _11427_/A vssd1 vssd1 vccd1 vccd1 _11536_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_111_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap107 _07556_/Y vssd1 vssd1 vccd1 vccd1 _10349_/A1 sky130_fd_sc_hd__buf_6
X_11467_ reg1_val[14] curr_PC[14] vssd1 vssd1 vccd1 vccd1 _11469_/A sky130_fd_sc_hd__or2_1
XANTENNA__10734__A _10734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13206_ _09145_/Y _13598_/C hold45/X _13605_/A vssd1 vssd1 vccd1 vccd1 _13639_/D
+ sky130_fd_sc_hd__o211a_1
X_10418_ _10259_/A _10258_/B _10256_/Y vssd1 vssd1 vccd1 vccd1 _10421_/A sky130_fd_sc_hd__a21oi_2
X_11398_ _11507_/A _11398_/B vssd1 vssd1 vccd1 vccd1 _11400_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13137_ hold169/X hold3/X hold191/X vssd1 vssd1 vccd1 vccd1 _13597_/B sky130_fd_sc_hd__and3_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ _10349_/A1 _10518_/A _10249_/X _10251_/Y vssd1 vssd1 vccd1 vccd1 _10350_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10581__B1 _10580_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ _13068_/A _13068_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[16] sky130_fd_sc_hd__xor2_4
XANTENNA__12322__A1 _09523_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12019_ _12019_/A _12019_/B vssd1 vssd1 vccd1 vccd1 _12021_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07560_ _07563_/A _07563_/B vssd1 vssd1 vccd1 vccd1 _07566_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08874__A _10236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07491_ _07492_/A _07492_/B vssd1 vssd1 vccd1 vccd1 _07491_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_75_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09230_ _09230_/A _09230_/B vssd1 vssd1 vccd1 vccd1 _09279_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_75_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09161_ _09161_/A fanout9/X vssd1 vssd1 vccd1 vccd1 _09288_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_84_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13004__B _13005_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08112_ _08112_/A _08112_/B vssd1 vssd1 vccd1 vccd1 _08116_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07002__B _10603_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09092_ _09092_/A _09318_/B vssd1 vssd1 vccd1 vccd1 _09092_/X sky130_fd_sc_hd__or2_1
XANTENNA__07804__A2 _11732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13338__B1 _13506_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08043_ _08043_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08155_/A sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout111_A _07494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06841__B _12981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout209_A _09381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07568__A1 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07568__B2 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09994_ _12130_/A _09994_/B _09994_/C vssd1 vssd1 vccd1 vccd1 _09996_/A sky130_fd_sc_hd__and3_1
XFILLER_0_86_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08945_ _08946_/A _08946_/B vssd1 vssd1 vccd1 vccd1 _08945_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09871__C _12235_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11116__A2 _11115_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06791__A2 _06936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08876_ _08877_/A _08876_/B _08876_/C vssd1 vssd1 vccd1 vccd1 _08889_/A sky130_fd_sc_hd__nand3_1
XANTENNA__10324__B1 _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07827_ _10263_/A _07827_/B vssd1 vssd1 vccd1 vccd1 _07996_/A sky130_fd_sc_hd__xnor2_2
X_07758_ _07814_/A _07814_/B vssd1 vssd1 vccd1 vccd1 _07815_/A sky130_fd_sc_hd__or2_1
XANTENNA__12077__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10627__A1 _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11922__B _12764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11824__B1 fanout3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07689_ fanout53/X _08866_/B2 _08950_/B fanout47/X vssd1 vssd1 vccd1 vccd1 _07690_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10819__A _11512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09428_ _13748_/A _13744_/A _09516_/A instruction[3] vssd1 vssd1 vccd1 vccd1 _10730_/B
+ sky130_fd_sc_hd__and4b_4
XFILLER_0_94_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout24_A fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10538__B _10787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09359_ _09359_/A _09359_/B vssd1 vssd1 vccd1 vccd1 _09380_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08048__A2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13692__CLK _13701_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11052__A1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11052__B2 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12370_ _11668_/B _12037_/X _12369_/B _12369_/X _12629_/B vssd1 vssd1 vccd1 vccd1
+ _12371_/B sky130_fd_sc_hd__a311o_2
XFILLER_0_34_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11321_ _11321_/A _11321_/B vssd1 vssd1 vccd1 vccd1 _11334_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_120_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09548__A2 _10522_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11252_ hold271/A _11252_/B _11369_/B vssd1 vssd1 vccd1 vccd1 _11252_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_120_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10203_ _10140_/A _10140_/B _10141_/Y vssd1 vssd1 vccd1 vccd1 _10293_/A sky130_fd_sc_hd__o21ai_4
X_11183_ _11185_/B vssd1 vssd1 vccd1 vccd1 _11184_/B sky130_fd_sc_hd__inv_2
X_10134_ _10134_/A _10134_/B vssd1 vssd1 vccd1 vccd1 _10137_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13584__B _13584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10065_ _09909_/A _09908_/B _09908_/A vssd1 vssd1 vccd1 vccd1 _10068_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10967_ _10967_/A _10967_/B vssd1 vssd1 vccd1 vccd1 _10968_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_15_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10094__A2 _07891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12706_ _12374_/A _12750_/B hold197/A vssd1 vssd1 vccd1 vccd1 _12706_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10898_ _11955_/A _10863_/Y _10866_/X _10897_/X vssd1 vssd1 vccd1 vccd1 _10898_/X
+ sky130_fd_sc_hd__o211a_1
X_13686_ _13701_/CLK hold94/X vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12637_ _12633_/Y _12636_/X _10730_/B vssd1 vssd1 vccd1 vccd1 _12637_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07247__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11043__A1 _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11043__B2 _07477_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12568_ _12568_/A _12568_/B _12568_/C vssd1 vssd1 vccd1 vccd1 _12569_/B sky130_fd_sc_hd__or3_1
XFILLER_0_108_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11519_ _11520_/A _11520_/B vssd1 vssd1 vccd1 vccd1 _11610_/B sky130_fd_sc_hd__nand2b_1
X_12499_ _12499_/A _12499_/B vssd1 vssd1 vccd1 vccd1 _12500_/B sky130_fd_sc_hd__and2_1
Xhold207 hold207/A vssd1 vssd1 vccd1 vccd1 hold207/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold218 hold218/A vssd1 vssd1 vccd1 vccd1 hold218/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 hold229/A vssd1 vssd1 vccd1 vccd1 hold229/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08869__A _09950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09464__S _09674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06991_ reg2_val[5] _07110_/A _12782_/B vssd1 vssd1 vccd1 vccd1 _06995_/B sky130_fd_sc_hd__a21o_2
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ _08730_/A _08730_/B vssd1 vssd1 vccd1 vccd1 _08758_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11295__A _11603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08661_ _08692_/A _08692_/B vssd1 vssd1 vccd1 vccd1 _08661_/X sky130_fd_sc_hd__and2_1
X_07612_ _09575_/A _07612_/B vssd1 vssd1 vccd1 vccd1 _07616_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__12059__B1 _09521_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08592_ _08645_/A _08603_/B vssd1 vssd1 vccd1 vccd1 _08592_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_72_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10609__A1 _07492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07543_ _07544_/A _07544_/B vssd1 vssd1 vccd1 vccd1 _07543_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_49_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10609__B2 _12754_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10639__A _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout159_A _13196_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13015__A _13015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12557__C _12666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07474_ _07474_/A _07474_/B vssd1 vssd1 vccd1 vccd1 _07474_/Y sky130_fd_sc_hd__nand2_1
X_09213_ _12421_/A _09213_/B vssd1 vssd1 vccd1 vccd1 _09221_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_118_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12854__A _13020_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09144_ _07061_/B _07062_/B _07595_/A _07521_/A vssd1 vssd1 vccd1 vccd1 _09146_/B
+ sky130_fd_sc_hd__a31o_4
XANTENNA__06852__A _06928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07789__A1 _10049_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07789__B2 _09173_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09075_ _09073_/A _09073_/B _12299_/A _12213_/B vssd1 vssd1 vccd1 vccd1 _09082_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08026_ _08026_/A _08026_/B vssd1 vssd1 vccd1 vccd1 _08108_/A sky130_fd_sc_hd__nor2_1
Xfanout1 hold234/A vssd1 vssd1 vccd1 vccd1 fanout1/X sky130_fd_sc_hd__buf_6
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08202__A2 _11732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07005__A3 _13000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ _09977_/A _09977_/B vssd1 vssd1 vccd1 vccd1 _09979_/B sky130_fd_sc_hd__xnor2_2
X_08928_ _08929_/B _08928_/B _08928_/C vssd1 vssd1 vccd1 vccd1 _08938_/A sky130_fd_sc_hd__nand3_2
XANTENNA__09702__A2 _09703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08859_ _08881_/A _08881_/B vssd1 vssd1 vccd1 vccd1 _08861_/B sky130_fd_sc_hd__and2_1
X_11870_ _07092_/B _11869_/X _12047_/C1 vssd1 vssd1 vccd1 vccd1 _11870_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10821_ _10821_/A _10821_/B vssd1 vssd1 vccd1 vccd1 _10823_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10226__A1_N wire122/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10752_ hold301/A _10752_/B vssd1 vssd1 vccd1 vccd1 _10885_/B sky130_fd_sc_hd__or2_1
X_13540_ _13540_/A _13540_/B vssd1 vssd1 vccd1 vccd1 _13540_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__12470__B1 _09519_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13471_ hold294/X _13550_/A2 _13470_/X _13563_/B2 vssd1 vssd1 vccd1 vccd1 _13472_/B
+ sky130_fd_sc_hd__a22o_1
X_10683_ _10684_/A _10684_/B vssd1 vssd1 vccd1 vccd1 _10685_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_125_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12764__A fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12422_ _12423_/A _12423_/B vssd1 vssd1 vccd1 vccd1 _12491_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07858__A _10266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09769__A2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06762__A _10734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12353_ _12353_/A _12353_/B vssd1 vssd1 vccd1 vccd1 _12355_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06988__C1 _13010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11304_ _11527_/A fanout9/X fanout4/X _07526_/Y vssd1 vssd1 vccd1 vccd1 _11305_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12284_ _12362_/B _12284_/B vssd1 vssd1 vccd1 vccd1 _12286_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11235_ _11463_/A _11235_/B vssd1 vssd1 vccd1 vccd1 _11235_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10536__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09941__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11166_ _11732_/A fanout34/X fanout32/X _07310_/Y vssd1 vssd1 vccd1 vccd1 _11167_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10117_ _10266_/A _10117_/B vssd1 vssd1 vccd1 vccd1 _10121_/A sky130_fd_sc_hd__xnor2_1
XANTENNA_max_cap73_A _07544_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_14_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13739_/CLK sky130_fd_sc_hd__clkbuf_8
X_11097_ _11097_/A _11097_/B vssd1 vssd1 vccd1 vccd1 _11099_/B sky130_fd_sc_hd__xnor2_1
X_10048_ _09954_/A _09954_/B _09952_/X vssd1 vssd1 vccd1 vccd1 _10063_/A sky130_fd_sc_hd__o21a_2
XANTENNA__11600__C_N _11458_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11500__A2 _07643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11999_ _12000_/A _12000_/B vssd1 vssd1 vccd1 vccd1 _12001_/A sky130_fd_sc_hd__or2_1
XFILLER_0_58_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13738_ _13739_/CLK hold4/X vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13669_ _13736_/CLK hold221/X vssd1 vssd1 vccd1 vccd1 hold219/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08680__A2 _10104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11016__A1 _12537_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07768__A _12421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07190_ _11793_/A _07297_/A vssd1 vssd1 vccd1 vccd1 _07190_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11016__B2 _12710_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09900_ fanout21/X _11423_/A fanout74/X fanout18/X vssd1 vssd1 vccd1 vccd1 _09901_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08599__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09393__B1 _08246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09831_ _09723_/Y _10726_/B _11955_/A vssd1 vssd1 vccd1 vccd1 _09831_/X sky130_fd_sc_hd__a21o_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ _09763_/A _09763_/B vssd1 vssd1 vccd1 vccd1 _09762_/Y sky130_fd_sc_hd__nand2_1
X_06974_ reg2_val[7] _06980_/B vssd1 vssd1 vccd1 vccd1 _06974_/X sky130_fd_sc_hd__and2_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08713_ _08714_/A _08714_/B vssd1 vssd1 vccd1 vccd1 _08713_/X sky130_fd_sc_hd__or2_1
X_09693_ _09694_/A curr_PC[1] vssd1 vssd1 vccd1 vccd1 _09695_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout276_A _13444_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08644_ _08582_/B _08644_/B vssd1 vssd1 vccd1 vccd1 _08645_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08575_ _08575_/A _08575_/B vssd1 vssd1 vccd1 vccd1 _08615_/A sky130_fd_sc_hd__nor2_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07526_ _07526_/A _07527_/B vssd1 vssd1 vccd1 vccd1 _07526_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_64_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07457_ fanout28/X _10049_/A2 _08395_/B _10915_/A vssd1 vssd1 vccd1 vccd1 _07458_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07388_ _07395_/A _07395_/B vssd1 vssd1 vccd1 vccd1 _11514_/A sky130_fd_sc_hd__and2_2
X_09127_ _10095_/A _09127_/B vssd1 vssd1 vccd1 vccd1 _09129_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12755__A1 _13129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09620__A1 fanout39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09620__B2 _08118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09058_ _08566_/X _08981_/B _08570_/X vssd1 vssd1 vccd1 vccd1 _09060_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_32_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10230__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08009_ _08016_/A _08016_/B vssd1 vssd1 vccd1 vccd1 _08009_/X sky130_fd_sc_hd__and2b_1
XANTENNA_fanout91_A _12420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11020_ curr_PC[9] curr_PC[10] _11020_/C vssd1 vssd1 vccd1 vccd1 _11265_/C sky130_fd_sc_hd__and3_1
XANTENNA__13180__A1 _13180_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07934__A1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11730__A2 _07643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07934__B2 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09136__B1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12971_ reg1_val[26] curr_PC[26] _12971_/S vssd1 vssd1 vccd1 vccd1 _12973_/B sky130_fd_sc_hd__mux2_1
X_11922_ _11922_/A _12764_/B vssd1 vssd1 vccd1 vccd1 _11923_/B sky130_fd_sc_hd__nand2_1
X_11853_ _11853_/A _11853_/B _11853_/C vssd1 vssd1 vccd1 vccd1 _11854_/B sky130_fd_sc_hd__nand3_2
XANTENNA__10049__A2 _10049_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10804_ fanout34/X _11423_/A _07543_/X fanout32/X vssd1 vssd1 vccd1 vccd1 _10805_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_95_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11784_ _12710_/B2 _11473_/X _11484_/X _12537_/B2 _11783_/X vssd1 vssd1 vccd1 vccd1
+ _11784_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13523_ _13523_/A _13523_/B vssd1 vssd1 vccd1 vccd1 _13523_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10735_ _10734_/A _06976_/Y _07037_/X _10734_/Y vssd1 vssd1 vccd1 vccd1 _10736_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10666_ _10666_/A _10666_/B vssd1 vssd1 vccd1 vccd1 _10668_/B sky130_fd_sc_hd__xnor2_1
X_13454_ _13450_/X _13453_/X _13459_/A vssd1 vssd1 vccd1 vccd1 hold263/A sky130_fd_sc_hd__o21a_1
XFILLER_0_125_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12405_ curr_PC[24] _12477_/C vssd1 vssd1 vccd1 vccd1 _12405_/X sky130_fd_sc_hd__and2_1
X_13385_ hold1/X _13444_/B1 _13384_/X vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__o21a_1
X_10597_ _09998_/X _10001_/X _10600_/S vssd1 vssd1 vccd1 vccd1 _10597_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12336_ _12336_/A _12336_/B vssd1 vssd1 vccd1 vccd1 _12353_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_23_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12267_ _12668_/A _12267_/B vssd1 vssd1 vccd1 vccd1 _12270_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11218_ _11219_/A _11219_/B vssd1 vssd1 vccd1 vccd1 _11340_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_120_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12198_ _12286_/A _12198_/B vssd1 vssd1 vccd1 vccd1 _12200_/B sky130_fd_sc_hd__nand2_1
X_11149_ _11382_/C _11148_/Y _12825_/S _11146_/X vssd1 vssd1 vccd1 vccd1 dest_val[11]
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_128_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07689__B1 _08950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11485__A1 _12537_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11485__B2 _12710_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08360_ _08360_/A _08360_/B vssd1 vssd1 vccd1 vccd1 _08364_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_58_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07311_ _10649_/A _07312_/B vssd1 vssd1 vccd1 vccd1 _07311_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_86_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08291_ _08291_/A _08291_/B vssd1 vssd1 vccd1 vccd1 _08292_/C sky130_fd_sc_hd__or2_1
XFILLER_0_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07242_ _07252_/D _07220_/Y _07221_/Y _07213_/Y vssd1 vssd1 vccd1 vccd1 _07242_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_27_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07173_ _10239_/A _07200_/B vssd1 vssd1 vccd1 vccd1 _07173_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_103_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07613__B1 _10235_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13162__A1 _07494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08122__A _08907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07916__A1 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07916__B2 _07699_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09814_ _09812_/A _09812_/B _09815_/B vssd1 vssd1 vccd1 vccd1 _09814_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__10920__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09745_ _09745_/A _09745_/B vssd1 vssd1 vccd1 vccd1 _09747_/B sky130_fd_sc_hd__xor2_1
X_06957_ reg1_val[10] _07455_/A vssd1 vssd1 vccd1 vccd1 _06958_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_69_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _09672_/X _09675_/X _10176_/A vssd1 vssd1 vccd1 vccd1 _09676_/X sky130_fd_sc_hd__mux2_1
X_06888_ _06886_/Y _06906_/B1 _06980_/B reg2_val[18] vssd1 vssd1 vccd1 vccd1 _07310_/A
+ sky130_fd_sc_hd__a2bb2o_2
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08627_ _08857_/A _08627_/B vssd1 vssd1 vccd1 vccd1 _08685_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_68_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08892__A2 _07399_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08558_ _08620_/A _08620_/B vssd1 vssd1 vccd1 vccd1 _08621_/A sky130_fd_sc_hd__or2_1
XFILLER_0_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07509_ _11372_/A _11372_/B _07572_/S vssd1 vssd1 vccd1 vccd1 _07517_/B sky130_fd_sc_hd__o21a_2
X_08489_ _09591_/A _08489_/B vssd1 vssd1 vccd1 vccd1 _08495_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10520_ _10520_/A _10520_/B vssd1 vssd1 vccd1 vccd1 _10521_/B sky130_fd_sc_hd__and2_1
XFILLER_0_92_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07201__A _07201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10451_ _10451_/A vssd1 vssd1 vccd1 vccd1 _10451_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_122_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07604__B1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13170_ _07477_/X _13194_/A2 hold52/X _13359_/A vssd1 vssd1 vccd1 vccd1 _13621_/D
+ sky130_fd_sc_hd__o211a_1
X_10382_ _10382_/A _10382_/B vssd1 vssd1 vccd1 vccd1 _10383_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_103_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12121_ _12121_/A _12121_/B vssd1 vssd1 vccd1 vccd1 _12440_/A sky130_fd_sc_hd__and2_2
XFILLER_0_20_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12052_ _12052_/A _12052_/B vssd1 vssd1 vccd1 vccd1 _12052_/X sky130_fd_sc_hd__xor2_1
XANTENNA__11164__B1 _07833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11003_ _12525_/A _11001_/X _11002_/Y _12760_/A1 vssd1 vssd1 vccd1 vccd1 _11003_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11703__A2 _12163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09372__A3 _10787_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12954_ _12961_/B _12954_/B vssd1 vssd1 vccd1 vccd1 new_PC[22] sky130_fd_sc_hd__xnor2_4
XFILLER_0_87_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11905_ _11905_/A _11905_/B vssd1 vssd1 vccd1 vccd1 _11906_/B sky130_fd_sc_hd__or2_1
X_12885_ _12886_/A _12886_/B _12886_/C vssd1 vssd1 vccd1 vccd1 _12893_/B sky130_fd_sc_hd__a21o_1
XANTENNA__13208__A2 _13598_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06853__A2_N _07110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12416__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11836_ _11722_/A _11722_/B _11725_/A vssd1 vssd1 vccd1 vccd1 _11838_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08635__A2 _09173_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11767_ _11703_/X _12163_/B _10730_/B vssd1 vssd1 vccd1 vccd1 _11767_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13506_ hold271/X _13506_/A2 _13505_/X _13506_/B2 vssd1 vssd1 vccd1 vccd1 hold272/A
+ sky130_fd_sc_hd__a22o_1
X_10718_ _10719_/A _10719_/B _10719_/C vssd1 vssd1 vccd1 vccd1 _10852_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_36_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11698_ _11669_/Y _11670_/X _11672_/Y _10866_/B _11697_/Y vssd1 vssd1 vccd1 vccd1
+ _11698_/X sky130_fd_sc_hd__o221a_1
XANTENNA__07111__A _13744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12719__B2 _12764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13437_ _12417_/A _13598_/C hold54/X vssd1 vssd1 vccd1 vccd1 _13700_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_24_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10649_ _10649_/A fanout6/X vssd1 vssd1 vccd1 vccd1 _10649_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_51_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13368_ hold216/X _13563_/B2 _13550_/A2 hold207/X vssd1 vssd1 vccd1 vccd1 hold217/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12319_ _12303_/A _12793_/A2 _09515_/Y _06856_/A _12318_/Y vssd1 vssd1 vccd1 vccd1
+ _12319_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_121_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13299_ _13250_/B _13523_/B _13248_/X vssd1 vssd1 vccd1 vccd1 _13527_/B sky130_fd_sc_hd__a21o_1
XANTENNA__13144__A1 _12764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11155__B1 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07860_ _09940_/A _07860_/B vssd1 vssd1 vccd1 vccd1 _07862_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10902__B1 _07548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06811_ _09254_/B vssd1 vssd1 vccd1 vccd1 _07061_/B sky130_fd_sc_hd__inv_2
X_07791_ fanout82/X fanout68/X fanout66/X fanout76/X vssd1 vssd1 vccd1 vccd1 _07792_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13447__A2 fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09530_ _09482_/X _09536_/B _09703_/B vssd1 vssd1 vccd1 vccd1 _09530_/X sky130_fd_sc_hd__mux2_1
X_09461_ _09459_/X _09460_/X _09674_/S vssd1 vssd1 vccd1 vccd1 _09461_/X sky130_fd_sc_hd__mux2_1
X_08412_ _08471_/A _08471_/B vssd1 vssd1 vccd1 vccd1 _08412_/X sky130_fd_sc_hd__and2_1
XFILLER_0_93_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09392_ _09406_/A vssd1 vssd1 vccd1 vccd1 _09392_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12407__B1 _12971_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08343_ _08343_/A _08343_/B vssd1 vssd1 vccd1 vccd1 _08371_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__09501__A _09501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08626__A2 _10104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout141_A _11231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout239_A _12971_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08274_ _08274_/A _08274_/B _08274_/C vssd1 vssd1 vccd1 vccd1 _08350_/A sky130_fd_sc_hd__or3_2
XFILLER_0_61_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10366__B fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07225_ _08197_/A fanout51/X _08907_/A fanout49/X vssd1 vssd1 vccd1 vccd1 _07226_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12862__A _13025_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07378__D _07378_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07156_ reg1_val[31] _11463_/A vssd1 vssd1 vccd1 vccd1 _07156_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__10197__A1 _11866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07087_ instruction[6] _07086_/Y _07075_/A vssd1 vssd1 vccd1 vccd1 _07087_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout100 _07310_/Y vssd1 vssd1 vccd1 vccd1 _10814_/A1 sky130_fd_sc_hd__buf_8
Xfanout111 _07494_/X vssd1 vssd1 vccd1 vccd1 _10637_/A sky130_fd_sc_hd__buf_6
Xfanout133 _09582_/A vssd1 vssd1 vccd1 vccd1 _08821_/B2 sky130_fd_sc_hd__clkbuf_8
Xfanout144 _07153_/X vssd1 vssd1 vccd1 vccd1 _11231_/A sky130_fd_sc_hd__clkbuf_4
Xfanout155 _08857_/A vssd1 vssd1 vccd1 vccd1 _10537_/A sky130_fd_sc_hd__clkbuf_8
Xfanout166 _13141_/Y vssd1 vssd1 vccd1 vccd1 _13207_/B sky130_fd_sc_hd__buf_4
Xfanout177 _07476_/B vssd1 vssd1 vccd1 vccd1 _07521_/A sky130_fd_sc_hd__buf_6
Xfanout188 _07118_/B vssd1 vssd1 vccd1 vccd1 _13584_/B sky130_fd_sc_hd__buf_4
Xfanout199 _09779_/A vssd1 vssd1 vccd1 vccd1 _09950_/A sky130_fd_sc_hd__buf_12
X_07989_ _07989_/A _07989_/B vssd1 vssd1 vccd1 vccd1 _08071_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__13438__A2 _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09728_ _10050_/A _09728_/B vssd1 vssd1 vccd1 vccd1 _09736_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_97_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09659_ _09659_/A _09659_/B vssd1 vssd1 vccd1 vccd1 _09660_/B sky130_fd_sc_hd__or2_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _12670_/A _12670_/B vssd1 vssd1 vccd1 vccd1 _12671_/C sky130_fd_sc_hd__or2_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _12417_/A _11621_/B vssd1 vssd1 vccd1 vccd1 _11622_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11552_ _11550_/Y _11552_/B vssd1 vssd1 vccd1 vccd1 _11761_/A sky130_fd_sc_hd__nand2b_4
XFILLER_0_80_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10503_ _10503_/A vssd1 vssd1 vccd1 vccd1 _10510_/A sky130_fd_sc_hd__inv_2
X_11483_ _09521_/Y _11476_/Y _11482_/X vssd1 vssd1 vccd1 vccd1 _11483_/X sky130_fd_sc_hd__a21o_1
X_10434_ _09827_/X _09828_/X _10435_/C vssd1 vssd1 vccd1 vccd1 _10434_/X sky130_fd_sc_hd__a21o_1
X_13222_ _13222_/A _13222_/B vssd1 vssd1 vccd1 vccd1 _13565_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_122_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10365_ _10537_/A _10365_/B vssd1 vssd1 vccd1 vccd1 _10369_/A sky130_fd_sc_hd__xor2_1
X_13153_ hold83/X _13193_/B vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__or2_1
XFILLER_0_103_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ _12105_/A _12105_/B vssd1 vssd1 vccd1 vccd1 _12192_/A sky130_fd_sc_hd__and2_1
X_13084_ _13102_/A _13084_/B _13084_/C vssd1 vssd1 vccd1 vccd1 _13085_/B sky130_fd_sc_hd__and3_2
XFILLER_0_20_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10296_ _10296_/A _10296_/B vssd1 vssd1 vccd1 vccd1 _10857_/A sky130_fd_sc_hd__xnor2_4
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12035_ _12035_/A _12035_/B vssd1 vssd1 vccd1 vccd1 _12037_/B sky130_fd_sc_hd__nor2_1
XANTENNA__13429__A2 _13598_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12637__B1 _10730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09502__B1 _12648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12937_ _12937_/A _12937_/B _12937_/C vssd1 vssd1 vccd1 vccd1 _12961_/A sky130_fd_sc_hd__or3_1
XFILLER_0_87_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11860__A1 _10984_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12868_ _13029_/B _12869_/B vssd1 vssd1 vccd1 vccd1 _12879_/A sky130_fd_sc_hd__nand2_1
X_11819_ _11819_/A _11819_/B vssd1 vssd1 vccd1 vccd1 _11820_/B sky130_fd_sc_hd__and2_1
XFILLER_0_7_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _07398_/B _12799_/A2 _12775_/Y _12798_/Y _12971_/S vssd1 vssd1 vccd1 vccd1
+ dest_val[31] sky130_fd_sc_hd__o221a_4
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11612__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11612__B2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09281__A2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07010_ _07008_/Y _07010_/B vssd1 vssd1 vccd1 vccd1 _10026_/A sky130_fd_sc_hd__and2b_1
XANTENNA__09467__S _09493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11376__B1 _11372_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_14_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09991__A _10577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08961_ _08951_/A _08953_/Y _08960_/A vssd1 vssd1 vccd1 vccd1 _08961_/Y sky130_fd_sc_hd__o21ai_1
X_07912_ _07912_/A _07912_/B vssd1 vssd1 vccd1 vccd1 _07927_/A sky130_fd_sc_hd__xnor2_1
X_08892_ _07175_/X _07399_/Y _09910_/A1 _08933_/B vssd1 vssd1 vccd1 vccd1 _08893_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07843_ _07843_/A _07843_/B vssd1 vssd1 vccd1 vccd1 _07844_/B sky130_fd_sc_hd__xnor2_1
X_07774_ _07774_/A _07774_/B vssd1 vssd1 vccd1 vccd1 _07845_/B sky130_fd_sc_hd__or2_1
X_09513_ _13744_/A _09516_/A _09525_/C vssd1 vssd1 vccd1 vccd1 _12781_/A sky130_fd_sc_hd__and3_2
XFILLER_0_94_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09444_ reg1_val[6] reg1_val[25] _09463_/S vssd1 vssd1 vccd1 vccd1 _09444_/X sky130_fd_sc_hd__mux2_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09375_ _09376_/A _09376_/B vssd1 vssd1 vccd1 vccd1 _09375_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10377__A _11719_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08326_ _08821_/B2 fanout82/X fanout76/X _08821_/A1 vssd1 vssd1 vccd1 vccd1 _08327_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12800__A0 _09501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09272__A2 _07643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10096__B fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08257_ _08257_/A _08257_/B _08257_/C vssd1 vssd1 vccd1 vccd1 _08260_/A sky130_fd_sc_hd__and3_1
XFILLER_0_62_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07208_ _07535_/B _07208_/B vssd1 vssd1 vccd1 vccd1 _07208_/X sky130_fd_sc_hd__or2_1
XANTENNA__12159__A2 _11793_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08188_ _08186_/A _08186_/B _08287_/A vssd1 vssd1 vccd1 vccd1 _08220_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07139_ _13744_/A instruction[5] vssd1 vssd1 vccd1 vccd1 _09507_/C sky130_fd_sc_hd__or2_1
XFILLER_0_113_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10150_ _10150_/A _10298_/A _10433_/A _10577_/A vssd1 vssd1 vccd1 vccd1 _10150_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_112_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10081_ _10081_/A _10081_/B vssd1 vssd1 vccd1 vccd1 _10082_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_69_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09840__S _10004_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10983_ _09830_/B _10435_/C _10981_/X _10982_/Y _10980_/Y vssd1 vssd1 vccd1 vccd1
+ _10984_/B sky130_fd_sc_hd__o311a_4
XFILLER_0_97_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12722_ _12723_/A _12722_/B vssd1 vssd1 vccd1 vccd1 _12722_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_38_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09141__A _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12653_ hold249/A _12653_/B vssd1 vssd1 vccd1 vccd1 _12702_/B sky130_fd_sc_hd__or2_1
XFILLER_0_127_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11604_ _12557_/B fanout20/X fanout18/X _07597_/X vssd1 vssd1 vccd1 vccd1 _11605_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12584_ _12584_/A _12584_/B vssd1 vssd1 vccd1 vccd1 _12584_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11535_ _11392_/A _11392_/B _11390_/X vssd1 vssd1 vccd1 vccd1 _11540_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__07596__A _10787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11466_ _11465_/A _11465_/B _11465_/Y _12047_/C1 vssd1 vssd1 vccd1 vccd1 _11466_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13205_ hold44/X _13207_/B vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__or2_1
XFILLER_0_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10417_ _10219_/A _10219_/B _10218_/A vssd1 vssd1 vccd1 vccd1 _10422_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11397_ fanout44/X fanout29/X fanout27/X _07597_/X vssd1 vssd1 vccd1 vccd1 _11398_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_104_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10030__B1 _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13136_ _13136_/A _13136_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[31] sky130_fd_sc_hd__xnor2_4
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _10249_/X _10251_/Y _10349_/A1 _10518_/A vssd1 vssd1 vccd1 vccd1 _10348_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10581__A1 _10300_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13537__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _13068_/A _13068_/B vssd1 vssd1 vccd1 vccd1 _13081_/A sky130_fd_sc_hd__or2_1
X_10279_ _10279_/A _10279_/B vssd1 vssd1 vccd1 vccd1 _10292_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_29_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12018_ _12016_/A _12016_/B _12019_/B vssd1 vssd1 vccd1 vccd1 _12110_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07490_ _07557_/A _07180_/C _07363_/B _07186_/B _07476_/B vssd1 vssd1 vccd1 vccd1
+ _07492_/B sky130_fd_sc_hd__a41o_4
XFILLER_0_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_504 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09160_ _12668_/A _09160_/B vssd1 vssd1 vccd1 vccd1 fanout9/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_56_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08111_ _08111_/A _08111_/B vssd1 vssd1 vccd1 vccd1 _08162_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09091_ _08105_/Y _08994_/B _08996_/Y vssd1 vssd1 vccd1 vccd1 _09094_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_114_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08042_ _08043_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08042_/X sky130_fd_sc_hd__or2_1
XFILLER_0_31_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11349__B1 _11600_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13020__B _13020_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout104_A _07276_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07568__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09993_ _12130_/A _10044_/A _10726_/C _11955_/A vssd1 vssd1 vccd1 vccd1 _09993_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_110_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08944_ _08944_/A _08944_/B vssd1 vssd1 vccd1 vccd1 _08946_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10660__A _11603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08875_ _08901_/A _08901_/B _08872_/C vssd1 vssd1 vccd1 vccd1 _08876_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07826_ _09216_/B2 fanout28/X _08395_/B _08868_/B1 vssd1 vssd1 vccd1 vccd1 _07827_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12077__A1 _07230_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07757_ _07757_/A _07757_/B vssd1 vssd1 vccd1 vccd1 _07814_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12077__B2 _12189_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10088__B1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11824__A1 _11997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07688_ _10050_/A _07694_/B vssd1 vssd1 vccd1 vccd1 _07688_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11824__B2 _11922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09427_ _09427_/A _10150_/A vssd1 vssd1 vccd1 vccd1 _10726_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10538__C _10787_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09358_ _09358_/A _09358_/B vssd1 vssd1 vccd1 vccd1 _09359_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08309_ _08309_/A _08309_/B vssd1 vssd1 vccd1 vccd1 _08311_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07256__A1 _07594_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11052__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09289_ _09289_/A _09289_/B _09289_/C vssd1 vssd1 vccd1 vccd1 _09414_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_35_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11320_ _11319_/A _11319_/B _11319_/C vssd1 vssd1 vccd1 vccd1 _11321_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08305__A _10236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11251_ hold291/A hold280/A _11251_/C vssd1 vssd1 vccd1 vccd1 _11369_/B sky130_fd_sc_hd__or3_1
XFILLER_0_105_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_515 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10202_ _10145_/A _10145_/B _10143_/X vssd1 vssd1 vccd1 vccd1 _10296_/A sky130_fd_sc_hd__a21oi_4
X_11182_ _11182_/A _11182_/B vssd1 vssd1 vccd1 vccd1 _11185_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10133_ _09898_/A _09897_/B _09897_/A vssd1 vssd1 vccd1 vccd1 _10138_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_100_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10064_ _09946_/A _09946_/B _09945_/A vssd1 vssd1 vccd1 vccd1 _10070_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__13501__B2 _13506_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12068__B2 _10866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10966_ _10966_/A _10966_/B vssd1 vssd1 vccd1 vccd1 _10967_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10729__B _11151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12705_ hold219/A _12705_/B vssd1 vssd1 vccd1 vccd1 _12750_/B sky130_fd_sc_hd__or2_1
X_13685_ _13701_/CLK hold122/X vssd1 vssd1 vccd1 vccd1 _13685_/Q sky130_fd_sc_hd__dfxtp_1
X_10897_ _10897_/A _10897_/B _10897_/C vssd1 vssd1 vccd1 vccd1 _10897_/X sky130_fd_sc_hd__and3_1
XFILLER_0_85_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12636_ _12373_/A _12373_/B _12635_/Y _12056_/B vssd1 vssd1 vccd1 vccd1 _12636_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_38_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07247__A1 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07247__B2 _08866_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12240__A1 _12710_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11043__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12567_ _12568_/A _12568_/B _12568_/C vssd1 vssd1 vccd1 vccd1 _12567_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_53_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12791__A2 _07398_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11518_ _12253_/A _11518_/B vssd1 vssd1 vccd1 vccd1 _11520_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_25_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12498_ _12499_/A _12499_/B vssd1 vssd1 vccd1 vccd1 _12568_/A sky130_fd_sc_hd__nor2_1
Xhold208 hold208/A vssd1 vssd1 vccd1 vccd1 hold208/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold219 hold219/A vssd1 vssd1 vccd1 vccd1 hold219/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11449_ _11449_/A _11449_/B _11449_/C vssd1 vssd1 vccd1 vccd1 _11450_/B sky130_fd_sc_hd__and3_1
XFILLER_0_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ reg1_val[28] _13136_/A vssd1 vssd1 vccd1 vccd1 _13120_/B sky130_fd_sc_hd__nand2_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06990_ reg2_val[5] _07110_/A _12782_/B vssd1 vssd1 vccd1 vccd1 _07180_/C sky130_fd_sc_hd__a21oi_4
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08660_ _08660_/A _08660_/B vssd1 vssd1 vccd1 vccd1 _08692_/B sky130_fd_sc_hd__xnor2_2
X_07611_ _11732_/A fanout68/X fanout66/X _10814_/A1 vssd1 vssd1 vccd1 vccd1 _07612_/B
+ sky130_fd_sc_hd__o22a_1
X_08591_ _08643_/A _08643_/B _08587_/Y vssd1 vssd1 vccd1 vccd1 _08603_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_49_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07542_ _07526_/A _07523_/A _07521_/B _07521_/A vssd1 vssd1 vccd1 vccd1 _07544_/B
+ sky130_fd_sc_hd__a31o_4
XANTENNA__10609__A2 _10889_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13015__B _13015_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07473_ _07473_/A _07473_/B vssd1 vssd1 vccd1 vccd1 _11283_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09212_ _07833_/B _10374_/B2 _10349_/A1 fanout14/X vssd1 vssd1 vccd1 vccd1 _09213_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10490__B1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09143_ _10239_/A _09143_/B vssd1 vssd1 vccd1 vccd1 _09150_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_8_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout221_A _10603_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06852__B _13020_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07789__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10242__B1 _08704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09074_ _09077_/A _09074_/B vssd1 vssd1 vccd1 vccd1 _12299_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08025_ _08024_/A _08024_/C _08024_/B vssd1 vssd1 vccd1 vccd1 _08026_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout2 hold234/A vssd1 vssd1 vccd1 vccd1 fanout2/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09976_ _09816_/A _09816_/B _09814_/X vssd1 vssd1 vccd1 vccd1 _09977_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_110_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08927_ _08920_/A _08920_/B _08920_/C vssd1 vssd1 vccd1 vccd1 _08928_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_99_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08858_ _08864_/A _08864_/B _08851_/Y vssd1 vssd1 vccd1 vccd1 _08881_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__08795__A _09373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07809_ _08021_/B _08021_/C _08021_/A vssd1 vssd1 vccd1 vccd1 _08022_/A sky130_fd_sc_hd__o21ai_1
X_08789_ _08789_/A _08789_/B vssd1 vssd1 vccd1 vccd1 _08814_/A sky130_fd_sc_hd__xnor2_1
X_10820_ _10821_/A _10821_/B vssd1 vssd1 vccd1 vccd1 _10937_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_94_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10751_ _07449_/A _11793_/B _12657_/B1 reg1_val[8] _10750_/Y vssd1 vssd1 vccd1 vccd1
+ _10751_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_55_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13470_ hold283/X _13469_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13470_/X sky130_fd_sc_hd__mux2_1
X_10682_ _10682_/A _10682_/B vssd1 vssd1 vccd1 vccd1 _10684_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12764__B _12764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12421_ _12421_/A _12421_/B vssd1 vssd1 vccd1 vccd1 _12423_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12352_ _12352_/A _12352_/B vssd1 vssd1 vccd1 vccd1 _12353_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_23_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11303_ _11302_/A _11302_/B _11302_/C vssd1 vssd1 vccd1 vccd1 _11311_/B sky130_fd_sc_hd__a21oi_1
X_12283_ _12283_/A _12283_/B _12283_/C vssd1 vssd1 vccd1 vccd1 _12284_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_105_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09926__B1 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11234_ _07093_/A _11120_/B _06950_/B vssd1 vssd1 vccd1 vccd1 _11235_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_31_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10536__A1 _10536_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10536__B2 _10536_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11396__A _11603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11165_ _12092_/A _11165_/B vssd1 vssd1 vccd1 vccd1 _11174_/A sky130_fd_sc_hd__xnor2_1
X_10116_ fanout20/X fanout74/X fanout70/X fanout18/X vssd1 vssd1 vccd1 vccd1 _10117_/B
+ sky130_fd_sc_hd__o22a_1
X_11096_ _11097_/A _11097_/B vssd1 vssd1 vccd1 vccd1 _11153_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_117_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10047_ _09977_/A _09977_/B _09978_/Y vssd1 vssd1 vccd1 vccd1 _10145_/A sky130_fd_sc_hd__o21ai_4
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_310 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11998_ _12087_/C _11998_/B vssd1 vssd1 vccd1 vccd1 _12000_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07114__A _13748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13737_ _13739_/CLK _13737_/D vssd1 vssd1 vccd1 vccd1 hold218/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08665__B1 _08271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10949_ _10950_/A _10950_/B vssd1 vssd1 vccd1 vccd1 _11029_/A sky130_fd_sc_hd__and2_1
XFILLER_0_42_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13668_ _13736_/CLK hold168/X vssd1 vssd1 vccd1 vccd1 _13668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12619_ _12620_/A _12671_/A vssd1 vssd1 vccd1 vccd1 _12677_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_109_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13599_ hold169/X hold3/X hold218/X _13599_/D vssd1 vssd1 vccd1 vccd1 _13599_/X sky130_fd_sc_hd__and4b_1
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09475__S _09493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13174__C1 _13543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09393__A1 _07471_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09830_ _10433_/A _09830_/B vssd1 vssd1 vccd1 vccd1 _10726_/B sky130_fd_sc_hd__xor2_2
XANTENNA__09393__B2 fanout85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ _10095_/A _09761_/B vssd1 vssd1 vccd1 vccd1 _09763_/B sky130_fd_sc_hd__xnor2_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06973_ _06971_/Y _06973_/B vssd1 vssd1 vccd1 vccd1 _10736_/A sky130_fd_sc_hd__and2b_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08712_ _08712_/A _08712_/B vssd1 vssd1 vccd1 vccd1 _08714_/B sky130_fd_sc_hd__xnor2_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09692_ _09677_/X _09691_/X _10458_/S vssd1 vssd1 vccd1 vccd1 _09692_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_83_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09504__A _10734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08643_ _08643_/A _08643_/B vssd1 vssd1 vccd1 vccd1 _08646_/A sky130_fd_sc_hd__xor2_1
XANTENNA_fanout171_A _12759_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout269_A _06920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08574_ _08574_/A _08574_/B vssd1 vssd1 vccd1 vccd1 _08575_/B sky130_fd_sc_hd__and2_1
XFILLER_0_89_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07024__A _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07525_ _07523_/A _07521_/B _07476_/B vssd1 vssd1 vccd1 vccd1 _07527_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_49_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11255__A2 _11587_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07456_ _07456_/A _07456_/B vssd1 vssd1 vccd1 vccd1 _07456_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_64_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07387_ _07386_/A _07386_/B _07865_/B vssd1 vssd1 vccd1 vccd1 _07395_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09126_ fanout47/X _10235_/A1 _10235_/B2 fanout45/X vssd1 vssd1 vccd1 vccd1 _09127_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_60_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12755__A2 _09254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09620__A2 _10915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09057_ _09057_/A _09057_/B vssd1 vssd1 vccd1 vccd1 _11957_/C sky130_fd_sc_hd__xor2_4
XANTENNA__12804__S _12825_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08008_ _08008_/A _08008_/B vssd1 vssd1 vccd1 vccd1 _08016_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07694__A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11715__B1 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13180__A2 _13194_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07934__A2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ _09960_/A _09960_/B vssd1 vssd1 vccd1 vccd1 _09959_/X sky130_fd_sc_hd__and2b_1
XANTENNA__09136__A1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09136__B2 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12970_ _12970_/A _12970_/B vssd1 vssd1 vccd1 vccd1 new_PC[25] sky130_fd_sc_hd__xnor2_4
XANTENNA__07147__B1 _06928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11921_ _11921_/A _11921_/B vssd1 vssd1 vccd1 vccd1 _11923_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_86_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11852_ _11853_/A _11853_/B _11853_/C vssd1 vssd1 vccd1 vccd1 _11852_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_67_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10803_ _11825_/A _10803_/B vssd1 vssd1 vccd1 vccd1 _10806_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11783_ _07435_/X _07436_/Y _12235_/C _11782_/X vssd1 vssd1 vccd1 vccd1 _11783_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13522_ _13539_/A _13522_/B vssd1 vssd1 vccd1 vccd1 _13720_/D sky130_fd_sc_hd__and2_1
X_10734_ _10734_/A _10734_/B vssd1 vssd1 vccd1 vccd1 _10734_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_27_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13453_ hold245/X fanout2/X _13452_/Y _13463_/B2 vssd1 vssd1 vccd1 vccd1 _13453_/X
+ sky130_fd_sc_hd__o211a_1
X_10665_ _10665_/A _10665_/B vssd1 vssd1 vccd1 vccd1 _10666_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_35_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10726__C _10726_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12404_ _10730_/B _12375_/Y _12376_/X _12379_/Y _12403_/X vssd1 vssd1 vccd1 vccd1
+ _12404_/X sky130_fd_sc_hd__a311o_1
X_13384_ hold149/X _13416_/A2 _09950_/A _13419_/A2 _13383_/A vssd1 vssd1 vccd1 vccd1
+ _13384_/X sky130_fd_sc_hd__o221a_1
X_10596_ _11576_/A _10595_/A _09535_/Y vssd1 vssd1 vccd1 vccd1 _10596_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__10757__A1 _09523_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12335_ _12335_/A _12335_/B vssd1 vssd1 vccd1 vccd1 _12355_/A sky130_fd_sc_hd__and2_1
X_12266_ _07257_/X fanout16/X fanout12/X _12496_/A vssd1 vssd1 vccd1 vccd1 _12267_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11706__B1 _07891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11217_ _11217_/A _11217_/B vssd1 vssd1 vccd1 vccd1 _11219_/B sky130_fd_sc_hd__xor2_1
X_12197_ _12197_/A _12197_/B vssd1 vssd1 vccd1 vccd1 _12198_/B sky130_fd_sc_hd__nand2_1
X_11148_ curr_PC[11] _11265_/C _10342_/A vssd1 vssd1 vccd1 vccd1 _11148_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13545__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11079_ _11079_/A _11079_/B vssd1 vssd1 vccd1 vccd1 _11082_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07689__A1 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07689__B2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10693__B1 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07310_ _07310_/A _07310_/B vssd1 vssd1 vccd1 vccd1 _07310_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_73_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08290_ _08290_/A _08290_/B _08290_/C vssd1 vssd1 vccd1 vccd1 _08291_/B sky130_fd_sc_hd__and3_1
XFILLER_0_128_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07241_ _07213_/Y _07221_/Y _07220_/Y _07252_/D vssd1 vssd1 vccd1 vccd1 _12331_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_116_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07172_ _08203_/A _07172_/B vssd1 vssd1 vccd1 vccd1 _07200_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_54_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07613__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07613__B2 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13162__A2 _13194_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09813_ _09617_/Y _09631_/B _09629_/Y vssd1 vssd1 vccd1 vccd1 _09815_/B sky130_fd_sc_hd__o21a_1
XANTENNA__07916__A2 _13149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10920__A1 _07282_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10920__B2 _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ _09745_/A _09745_/B vssd1 vssd1 vccd1 vccd1 _09896_/A sky130_fd_sc_hd__or2_1
X_06956_ reg1_val[10] _07455_/A vssd1 vssd1 vccd1 vccd1 _06956_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__06858__A _06928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09234__A _09575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09675_ _09673_/X _09674_/X _10005_/S vssd1 vssd1 vccd1 vccd1 _09675_/X sky130_fd_sc_hd__mux2_1
X_06887_ reg2_val[18] _06980_/B _06906_/B1 _06886_/Y vssd1 vssd1 vccd1 vccd1 _07309_/A
+ sky130_fd_sc_hd__o2bb2a_4
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08626_ _08806_/A2 _10104_/A _10225_/A _08806_/B1 vssd1 vssd1 vccd1 vccd1 _08627_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ _08557_/A _08557_/B vssd1 vssd1 vccd1 vccd1 _08620_/B sky130_fd_sc_hd__nand2_1
X_07508_ _11126_/A reg1_val[12] _07328_/B reg1_val[13] vssd1 vssd1 vccd1 vccd1 _11372_/B
+ sky130_fd_sc_hd__o31a_1
X_08488_ _08873_/B2 fanout84/X _08580_/B _13149_/A vssd1 vssd1 vccd1 vccd1 _08489_/B
+ sky130_fd_sc_hd__o22a_1
X_07439_ _07445_/A _07445_/B vssd1 vssd1 vccd1 vccd1 _11708_/A sky130_fd_sc_hd__nand2_8
XANTENNA__13203__B _13207_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10319__S _10457_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10450_ _11472_/S _09690_/X _09534_/C vssd1 vssd1 vccd1 vccd1 _10451_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__07201__B _07201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09109_ _09110_/A _09110_/B vssd1 vssd1 vccd1 vccd1 _09111_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_60_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07604__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07604__B2 _10235_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10381_ _10382_/A _10382_/B vssd1 vssd1 vccd1 vccd1 _10381_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_103_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12120_ _12120_/A _12120_/B _12120_/C vssd1 vssd1 vccd1 vccd1 _12121_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_102_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12051_ _11967_/A _11967_/B _11965_/B vssd1 vssd1 vccd1 vccd1 _12052_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11164__A1 _11922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11164__B2 _11997_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09843__S _10004_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11002_ _10998_/Y _10999_/X _12525_/A vssd1 vssd1 vccd1 vccd1 _11002_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11674__A _12515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12953_ _12940_/Y _12961_/C _12963_/B vssd1 vssd1 vccd1 vccd1 _12954_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__08868__B1 _08868_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11904_ _11905_/A _11905_/B vssd1 vssd1 vccd1 vccd1 _11906_/A sky130_fd_sc_hd__nand2_1
X_12884_ _12893_/A _12884_/B vssd1 vssd1 vccd1 vccd1 _12886_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12416__A1 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11835_ _11733_/A _11733_/B _11736_/A vssd1 vssd1 vccd1 vccd1 _11841_/A sky130_fd_sc_hd__a21o_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07599__A _09950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11766_ _11948_/A _11766_/B vssd1 vssd1 vccd1 vccd1 _12163_/B sky130_fd_sc_hd__xnor2_4
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13505_ hold291/A _13504_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13505_/X sky130_fd_sc_hd__mux2_1
X_10717_ _10717_/A _10717_/B vssd1 vssd1 vccd1 vccd1 _10719_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11697_ _11676_/Y _11677_/X _11696_/X vssd1 vssd1 vccd1 vccd1 _11697_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13436_ hold53/X _13142_/A _13444_/B1 hold25/X _13568_/A vssd1 vssd1 vccd1 vccd1
+ hold54/A sky130_fd_sc_hd__o221a_1
XFILLER_0_24_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10648_ _11076_/A _10648_/B vssd1 vssd1 vccd1 vccd1 _10652_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13367_ _13547_/A hold230/X vssd1 vssd1 vccd1 vccd1 _13665_/D sky130_fd_sc_hd__and2_1
XFILLER_0_106_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10579_ _10579_/A _10579_/B _10579_/C vssd1 vssd1 vccd1 vccd1 _10579_/X sky130_fd_sc_hd__or3_1
XFILLER_0_2_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12318_ _06856_/B _09520_/X _12317_/X vssd1 vssd1 vccd1 vccd1 _12318_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13298_ _13518_/B _13519_/A _13251_/X vssd1 vssd1 vccd1 vccd1 _13523_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_121_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13144__A2 _13598_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12249_ _12420_/A _12249_/B vssd1 vssd1 vccd1 vccd1 _12255_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11155__A1 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10902__A1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10902__B2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06810_ _06809_/Y _06872_/B1 _06873_/B1 reg2_val[29] vssd1 vssd1 vccd1 vccd1 _09254_/B
+ sky130_fd_sc_hd__a2bb2o_4
X_07790_ _09591_/A _07790_/B vssd1 vssd1 vccd1 vccd1 _07796_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09460_ reg1_val[10] reg1_val[21] _09463_/S vssd1 vssd1 vccd1 vccd1 _09460_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08893__A _09948_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08411_ _08411_/A _08411_/B vssd1 vssd1 vccd1 vccd1 _08471_/B sky130_fd_sc_hd__xnor2_2
X_09391_ _09221_/A _09221_/B _09220_/A vssd1 vssd1 vccd1 vccd1 _09406_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08342_ _08406_/A _08341_/B _08337_/X vssd1 vssd1 vccd1 vccd1 _08371_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_46_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08273_ _08272_/B _08272_/C _09659_/B vssd1 vssd1 vccd1 vccd1 _08274_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__07834__A1 _12421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07021__B _07025_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07224_ _07252_/B _07224_/B vssd1 vssd1 vccd1 vccd1 _12413_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_73_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07155_ reg1_val[31] _11463_/A vssd1 vssd1 vccd1 vccd1 _07155_/X sky130_fd_sc_hd__and2_1
XANTENNA__07598__B1 _07597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07086_ _12778_/A _07085_/Y _06794_/A vssd1 vssd1 vccd1 vccd1 _07086_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_112_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11146__B2 _11866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07972__A _09575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09663__S _09703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout123 _07451_/X vssd1 vssd1 vccd1 vccd1 _10049_/A2 sky130_fd_sc_hd__buf_6
XFILLER_0_100_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout134 _12742_/A vssd1 vssd1 vccd1 vccd1 _11562_/A sky130_fd_sc_hd__buf_4
Xfanout145 _09575_/A vssd1 vssd1 vccd1 vccd1 _11076_/A sky130_fd_sc_hd__buf_8
Xfanout156 _07295_/X vssd1 vssd1 vccd1 vccd1 _08857_/A sky130_fd_sc_hd__buf_12
Xfanout167 _09504_/Y vssd1 vssd1 vccd1 vccd1 _12537_/B2 sky130_fd_sc_hd__buf_4
XANTENNA__11494__A _11825_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout178 _07177_/Y vssd1 vssd1 vccd1 vccd1 _07476_/B sky130_fd_sc_hd__buf_8
X_07988_ _07989_/A _07989_/B vssd1 vssd1 vccd1 vccd1 _07988_/X sky130_fd_sc_hd__or2_1
Xfanout189 _09524_/Y vssd1 vssd1 vccd1 vccd1 _12533_/B1 sky130_fd_sc_hd__clkbuf_8
X_09727_ fanout35/X _10522_/A _09885_/B1 _07699_/B vssd1 vssd1 vccd1 vccd1 _09728_/B
+ sky130_fd_sc_hd__o22a_2
X_06939_ reg1_val[12] _07476_/A vssd1 vssd1 vccd1 vccd1 _06939_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_69_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10657__B1 _11638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09658_ _10730_/B _09658_/B _09658_/C vssd1 vssd1 vccd1 vccd1 _09658_/X sky130_fd_sc_hd__and3_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08609_ _08609_/A _08609_/B vssd1 vssd1 vccd1 vccd1 _08658_/A sky130_fd_sc_hd__xnor2_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _09753_/A _09588_/C _09588_/A vssd1 vssd1 vccd1 vccd1 _09600_/B sky130_fd_sc_hd__a21o_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _12103_/A fanout34/X fanout32/X fanout54/X vssd1 vssd1 vccd1 vccd1 _11621_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_92_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07212__A _07230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11551_ _11551_/A _11551_/B _11551_/C vssd1 vssd1 vccd1 vccd1 _11552_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_108_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10502_ _11281_/A _10502_/B vssd1 vssd1 vccd1 vccd1 _10503_/A sky130_fd_sc_hd__xnor2_1
X_11482_ _07513_/X _12754_/C _09523_/Y _11478_/Y _11481_/Y vssd1 vssd1 vccd1 vccd1
+ _11482_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_123_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13221_ hold278/A hold46/X vssd1 vssd1 vccd1 vccd1 _13222_/B sky130_fd_sc_hd__and2b_1
X_10433_ _10433_/A _10577_/A _10631_/A _10857_/A vssd1 vssd1 vccd1 vccd1 _10435_/C
+ sky130_fd_sc_hd__or4_2
XFILLER_0_21_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10188__A2 _12314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07589__B1 _08950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13152_ hold7/X _13193_/B _13151_/Y _13543_/A vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__o211a_1
X_10364_ _10536_/A1 _12667_/A _10536_/A2 _10536_/B2 vssd1 vssd1 vccd1 vccd1 _10365_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10593__C1 _12047_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12103_ _12103_/A _12666_/A vssd1 vssd1 vccd1 vccd1 _12105_/B sky130_fd_sc_hd__nor2_1
X_13083_ _13084_/B _13084_/C _13102_/A vssd1 vssd1 vccd1 vccd1 _13085_/A sky130_fd_sc_hd__a21oi_4
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10295_ _10296_/A _10296_/B vssd1 vssd1 vccd1 vccd1 _10295_/X sky130_fd_sc_hd__and2_1
X_12034_ _11852_/Y _11943_/Y _11945_/B vssd1 vssd1 vccd1 vccd1 _12207_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_88_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12936_ _12936_/A _12936_/B vssd1 vssd1 vccd1 vccd1 _12951_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_88_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12867_ reg1_val[10] curr_PC[10] _12867_/S vssd1 vssd1 vccd1 vccd1 _12869_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_56_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11818_ _11819_/A _11819_/B vssd1 vssd1 vccd1 vccd1 _11929_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_68_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09266__B1 _13135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12798_ _09507_/X _12778_/X _12797_/X vssd1 vssd1 vccd1 vccd1 _12798_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11073__B1 _07891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11612__A2 _07891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11749_ _11749_/A _11749_/B vssd1 vssd1 vccd1 vccd1 _11751_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09569__A1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09569__B2 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13419_ _07443_/X _13419_/A2 hold152/X vssd1 vssd1 vccd1 vccd1 hold153/A sky130_fd_sc_hd__o21a_1
XFILLER_0_59_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08960_ _08960_/A _08960_/B vssd1 vssd1 vccd1 vccd1 _09008_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09483__S _09839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07911_ _07911_/A _07911_/B vssd1 vssd1 vccd1 vccd1 _07912_/B sky130_fd_sc_hd__xor2_2
XANTENNA__07792__A _09575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08891_ _09674_/S _08891_/B vssd1 vssd1 vccd1 vccd1 _08902_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_75_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07842_ _07842_/A _07842_/B vssd1 vssd1 vccd1 vccd1 _07844_/A sky130_fd_sc_hd__xor2_1
XANTENNA__10887__B1 _12748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07752__B1 _09885_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07773_ _07774_/A _07774_/B vssd1 vssd1 vccd1 vccd1 _07773_/Y sky130_fd_sc_hd__nor2_1
X_09512_ _09524_/A _09516_/A instruction[4] _13744_/A vssd1 vssd1 vccd1 vccd1 _12598_/C
+ sky130_fd_sc_hd__or4b_4
XANTENNA__07016__B _10456_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11150__B1_N _10984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09443_ _13015_/A reg1_val[24] _09463_/S vssd1 vssd1 vccd1 vccd1 _09443_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_94_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10658__A _12421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout251_A _13141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06855__B _07230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09257__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09374_ _08271_/A fanout6/X _09949_/A vssd1 vssd1 vccd1 vccd1 _09376_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_47_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08128__A _09951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08325_ _08343_/A _08343_/B vssd1 vssd1 vccd1 vccd1 _08325_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_62_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08256_ _08256_/A _08256_/B vssd1 vssd1 vccd1 vccd1 _08257_/C sky130_fd_sc_hd__and2_1
XFILLER_0_7_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06871__A _06886_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07207_ _12982_/A _09694_/A vssd1 vssd1 vccd1 vccd1 _07208_/B sky130_fd_sc_hd__xor2_1
XANTENNA__13356__A2 _13506_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08187_ _08286_/A _08286_/B vssd1 vssd1 vccd1 vccd1 _08287_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07138_ instruction[5] _09516_/B vssd1 vssd1 vccd1 vccd1 _09529_/B sky130_fd_sc_hd__or2_4
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07069_ _12581_/A _07068_/X _07082_/A vssd1 vssd1 vccd1 vccd1 _07069_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_100_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10080_ _10080_/A _10080_/B vssd1 vssd1 vccd1 vccd1 _10081_/B sky130_fd_sc_hd__or2_1
XANTENNA__07207__A _12982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10982_ _10438_/A _10438_/B _10981_/X vssd1 vssd1 vccd1 vccd1 _10982_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_0_97_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12721_ _12723_/B vssd1 vssd1 vccd1 vccd1 _12722_/B sky130_fd_sc_hd__inv_2
XFILLER_0_38_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12652_ hold219/A _12735_/A1 _12705_/B _12651_/Y _12795_/A1 vssd1 vssd1 vccd1 vccd1
+ _12661_/C sky130_fd_sc_hd__a311o_1
XFILLER_0_127_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11603_ _11603_/A _11603_/B vssd1 vssd1 vccd1 vccd1 _11607_/A sky130_fd_sc_hd__xnor2_1
X_12583_ _12695_/A _12583_/B vssd1 vssd1 vccd1 vccd1 _12584_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_93_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10802__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11534_ _11428_/A _11428_/B _11431_/A vssd1 vssd1 vccd1 vccd1 _11544_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_108_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07596__B _10787_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11465_ _11465_/A _11465_/B vssd1 vssd1 vccd1 vccd1 _11465_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13204_ _12667_/A _13598_/C hold31/X _13605_/A vssd1 vssd1 vccd1 vccd1 _13638_/D
+ sky130_fd_sc_hd__o211a_1
X_10416_ _10279_/A _10279_/B _10278_/A vssd1 vssd1 vccd1 vccd1 _10426_/A sky130_fd_sc_hd__a21o_1
X_11396_ _11603_/A _11396_/B vssd1 vssd1 vccd1 vccd1 _11400_/A sky130_fd_sc_hd__xnor2_1
X_13135_ _13135_/A _13135_/B vssd1 vssd1 vccd1 vccd1 _13136_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10347_ _10241_/A _10241_/B _10239_/Y vssd1 vssd1 vccd1 vccd1 _10351_/A sky130_fd_sc_hd__a21o_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ reg1_val[15] _13059_/B _13062_/A vssd1 vssd1 vccd1 vccd1 _13068_/B sky130_fd_sc_hd__a21oi_2
X_10278_ _10278_/A _10278_/B vssd1 vssd1 vccd1 vccd1 _10279_/B sky130_fd_sc_hd__nor2_2
X_12017_ _11923_/A _11923_/B _11921_/A vssd1 vssd1 vccd1 vccd1 _12019_/B sky130_fd_sc_hd__o21a_1
XANTENNA__07117__A _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10097__B2 _10239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11294__B1 _07368_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12919_ _12956_/A _12920_/B vssd1 vssd1 vccd1 vccd1 _12938_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08110_ _08164_/A _08164_/B vssd1 vssd1 vccd1 vccd1 _08167_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09478__S _09493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09090_ _12583_/B _12584_/A vssd1 vssd1 vccd1 vccd1 _09090_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_16_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08041_ _08041_/A _08041_/B vssd1 vssd1 vccd1 vccd1 _08043_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__13338__A2 _13506_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09992_ _12130_/A _10044_/A _10726_/C vssd1 vssd1 vccd1 vccd1 _09992_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07973__B1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08943_ _08959_/A _08959_/B vssd1 vssd1 vccd1 vccd1 _08946_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08874_ _10236_/A _08874_/B vssd1 vssd1 vccd1 vccd1 _08876_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07725__B1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10324__A2 _12793_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07825_ _07828_/A _07828_/B vssd1 vssd1 vccd1 vccd1 _07825_/X sky130_fd_sc_hd__and2_1
XANTENNA__12868__A _13029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07756_ _10263_/A _07756_/B vssd1 vssd1 vccd1 vccd1 _07814_/A sky130_fd_sc_hd__xor2_1
XANTENNA__12077__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10088__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10088__B2 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07687_ _07687_/A _07687_/B vssd1 vssd1 vccd1 vccd1 _07694_/B sky130_fd_sc_hd__xor2_2
XANTENNA__10388__A _11913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11824__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09426_ _09426_/A _09426_/B vssd1 vssd1 vccd1 vccd1 _10150_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_66_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09357_ _09357_/A _09357_/B vssd1 vssd1 vccd1 vccd1 _09358_/B sky130_fd_sc_hd__or2_1
XANTENNA__13577__A2 _13584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08308_ _08377_/A _08377_/B vssd1 vssd1 vccd1 vccd1 _08311_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_74_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09288_ _09288_/A _10522_/B vssd1 vssd1 vccd1 vccd1 _09289_/C sky130_fd_sc_hd__and2_1
XFILLER_0_7_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08239_ _08239_/A _08239_/B vssd1 vssd1 vccd1 vccd1 _08242_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_34_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11250_ hold214/A _11693_/A2 _11366_/B _12533_/B1 vssd1 vssd1 vccd1 vccd1 _11250_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_0_120_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10201_ _12130_/A _10344_/A vssd1 vssd1 vccd1 vccd1 _10201_/X sky130_fd_sc_hd__and2_1
X_11181_ _11182_/A _11182_/B vssd1 vssd1 vccd1 vccd1 _11315_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11760__A1 _11550_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10132_ _09968_/A _09968_/B _09967_/A vssd1 vssd1 vccd1 vccd1 _10142_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13501__A2 _13506_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10063_ _10063_/A _10063_/B vssd1 vssd1 vccd1 vccd1 _10131_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_15_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11276__B1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10965_ _10964_/A _10964_/B _10966_/A vssd1 vssd1 vccd1 vccd1 _10965_/X sky130_fd_sc_hd__a21bo_1
X_12704_ hold299/A _12786_/B1 _12746_/B _12748_/B1 vssd1 vssd1 vccd1 vccd1 _12704_/X
+ sky130_fd_sc_hd__a31o_1
X_13684_ _13684_/CLK _13684_/D vssd1 vssd1 vccd1 vccd1 hold120/A sky130_fd_sc_hd__dfxtp_1
X_10896_ _09860_/A _10879_/Y _12225_/B _09839_/A _10893_/X vssd1 vssd1 vccd1 vccd1
+ _10897_/C sky130_fd_sc_hd__o221a_1
X_12635_ _12635_/A _12635_/B _12635_/C vssd1 vssd1 vccd1 vccd1 _12635_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12776__B1 _10734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap11_A _09145_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07247__A2 _08950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12566_ _12625_/B _12566_/B vssd1 vssd1 vccd1 vccd1 _12568_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07400__A _10004_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11517_ fanout46/X fanout38/X fanout36/X fanout50/X vssd1 vssd1 vccd1 vccd1 _11518_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_108_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12497_ _12557_/D _12497_/B vssd1 vssd1 vccd1 vccd1 _12499_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold209 hold209/A vssd1 vssd1 vccd1 vccd1 hold209/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11448_ _11449_/A _11449_/B _11449_/C vssd1 vssd1 vccd1 vccd1 _11450_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_111_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11379_ _12537_/B2 _11364_/X _11365_/X _12760_/A1 _11378_/Y vssd1 vssd1 vccd1 vccd1
+ _11379_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13118_ reg1_val[28] _13136_/A vssd1 vssd1 vccd1 vccd1 _13120_/A sky130_fd_sc_hd__or2_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ _13049_/A _13057_/A vssd1 vssd1 vccd1 vccd1 _13051_/C sky130_fd_sc_hd__nand2_1
XANTENNA__12700__B1 _12782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07610_ _10078_/A _07610_/B vssd1 vssd1 vccd1 vccd1 _07617_/A sky130_fd_sc_hd__xnor2_2
X_08590_ _09371_/A _08590_/B vssd1 vssd1 vccd1 vccd1 _08643_/B sky130_fd_sc_hd__xnor2_2
X_07541_ _10507_/A _11157_/A _07538_/X vssd1 vssd1 vccd1 vccd1 _07541_/X sky130_fd_sc_hd__a21o_4
XFILLER_0_72_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07472_ _07472_/A _07472_/B vssd1 vssd1 vccd1 vccd1 _07472_/Y sky130_fd_sc_hd__xnor2_4
X_09211_ _09154_/A _09154_/B _09152_/Y vssd1 vssd1 vccd1 vccd1 _09225_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__10490__A1 _07299_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13559__A2 _13584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10490__B2 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09142_ _07200_/Y fanout51/X fanout49/X _09582_/A vssd1 vssd1 vccd1 vccd1 _09143_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_16_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10242__A1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09073_ _09073_/A _09073_/B vssd1 vssd1 vccd1 vccd1 _12214_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10242__B2 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12519__B1 _10866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08024_ _08024_/A _08024_/B _08024_/C vssd1 vssd1 vccd1 vccd1 _08026_/A sky130_fd_sc_hd__and3_1
XFILLER_0_71_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout3 fanout4/X vssd1 vssd1 vccd1 vccd1 fanout3/X sky130_fd_sc_hd__buf_6
XFILLER_0_114_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09975_ _09975_/A _09975_/B vssd1 vssd1 vccd1 vccd1 _09977_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_110_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08926_ _08926_/A vssd1 vssd1 vccd1 vccd1 _08928_/B sky130_fd_sc_hd__inv_2
XANTENNA__09671__S _09671_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08857_ _08857_/A _08857_/B vssd1 vssd1 vccd1 vccd1 _08864_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07174__A1 _10239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07808_ _07808_/A _08008_/B vssd1 vssd1 vccd1 vccd1 _08021_/C sky130_fd_sc_hd__nor2_1
X_08788_ _08788_/A _08788_/B vssd1 vssd1 vccd1 vccd1 _09033_/A sky130_fd_sc_hd__xor2_2
XANTENNA__06921__A1 _06936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11258__B1 _11257_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07739_ fanout42/X _10235_/B2 _10814_/A1 _10235_/A1 vssd1 vssd1 vccd1 vccd1 _07740_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_94_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10750_ _10750_/A _10750_/B _12235_/C vssd1 vssd1 vccd1 vccd1 _10750_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_67_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09409_ _09409_/A _09409_/B vssd1 vssd1 vccd1 vccd1 _09410_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_54_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10681_ _10682_/B _10682_/A vssd1 vssd1 vccd1 vccd1 _10838_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_109_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12420_ _12420_/A _12421_/B vssd1 vssd1 vccd1 vccd1 _12491_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08316__A _09591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12351_ _12351_/A _12351_/B _12351_/C vssd1 vssd1 vccd1 vccd1 _12352_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_62_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11302_ _11302_/A _11302_/B _11302_/C vssd1 vssd1 vccd1 vccd1 _11311_/A sky130_fd_sc_hd__and3_1
XANTENNA__11981__A1 _09521_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12282_ _12283_/A _12283_/B _12283_/C vssd1 vssd1 vccd1 vccd1 _12362_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_105_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11233_ _11233_/A _11233_/B vssd1 vssd1 vccd1 vccd1 _11233_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__09926__A1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09926__B2 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10536__A2 _10536_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11164_ _11922_/A fanout14/X _07833_/B _11997_/A vssd1 vssd1 vccd1 vccd1 _11165_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10115_ _10115_/A vssd1 vssd1 vccd1 vccd1 _10127_/A sky130_fd_sc_hd__inv_2
X_11095_ _11095_/A _11095_/B vssd1 vssd1 vccd1 vccd1 _11097_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13486__B2 _13542_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10046_ _09982_/A _09982_/B _09980_/X vssd1 vssd1 vccd1 vccd1 _10148_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_117_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
X_11997_ _11997_/A _12666_/A vssd1 vssd1 vccd1 vccd1 _11998_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_85_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08665__A1 _12982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10948_ _11709_/A _10948_/B vssd1 vssd1 vccd1 vccd1 _10950_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13736_ _13736_/CLK hold142/X vssd1 vssd1 vccd1 vccd1 hold140/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08665__B2 _13168_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10879_ _10879_/A vssd1 vssd1 vccd1 vccd1 _10879_/Y sky130_fd_sc_hd__inv_2
X_13667_ _13705_/CLK _13667_/D vssd1 vssd1 vccd1 vccd1 hold166/A sky130_fd_sc_hd__dfxtp_1
X_12618_ _07876_/Y fanout7/X _12617_/Y _11823_/A vssd1 vssd1 vccd1 vccd1 _12671_/A
+ sky130_fd_sc_hd__a22o_1
X_13598_ _13597_/X hold169/X _13598_/C vssd1 vssd1 vccd1 vccd1 hold170/A sky130_fd_sc_hd__and3b_1
XFILLER_0_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12549_ _12666_/A _12549_/B vssd1 vssd1 vccd1 vccd1 _12551_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11421__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_1 _07548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10491__A _11603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09393__A2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09760_ _10235_/B2 _10787_/B _10787_/C _10235_/A1 fanout44/X vssd1 vssd1 vccd1 vccd1
+ _09761_/B sky130_fd_sc_hd__o32a_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06972_ reg1_val[8] _07184_/D vssd1 vssd1 vccd1 vccd1 _06973_/B sky130_fd_sc_hd__nand2_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08711_ _08744_/A _08744_/B vssd1 vssd1 vccd1 vccd1 _08714_/A sky130_fd_sc_hd__nand2b_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09691_ _09684_/X _09690_/X _11472_/S vssd1 vssd1 vccd1 vccd1 _09691_/X sky130_fd_sc_hd__mux2_1
X_08642_ _08642_/A _08642_/B vssd1 vssd1 vccd1 vccd1 _08650_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07305__A _10095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08573_ _08573_/A _08573_/B vssd1 vssd1 vccd1 vccd1 _08980_/A sky130_fd_sc_hd__xnor2_2
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout164_A _13193_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07524_ _07524_/A _11410_/A vssd1 vssd1 vccd1 vccd1 _07524_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_76_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07024__B _10004_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07455_ _07455_/A _07456_/B vssd1 vssd1 vccd1 vccd1 _07455_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_9_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07386_ _07386_/A _07386_/B vssd1 vssd1 vccd1 vccd1 _07386_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_106_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09125_ _09575_/A _09125_/B vssd1 vssd1 vccd1 vccd1 _09129_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09666__S _09703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09056_ _11864_/C _11864_/D _11864_/B vssd1 vssd1 vccd1 vccd1 _11957_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08007_ _08044_/A _08044_/B _08003_/X vssd1 vssd1 vccd1 vccd1 _08016_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_4_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11715__A1 _12331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11715__B2 _12413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09958_ _10522_/B _09958_/B vssd1 vssd1 vccd1 vccd1 _09960_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09136__A2 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08909_ _08908_/B _08908_/C _09659_/B vssd1 vssd1 vccd1 vccd1 _08910_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__11479__B1 _11586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07147__A1 _12578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09889_ _11731_/A _09889_/B vssd1 vssd1 vccd1 vccd1 _09893_/A sky130_fd_sc_hd__xnor2_1
X_11920_ _11920_/A _11920_/B vssd1 vssd1 vccd1 vccd1 _11921_/B sky130_fd_sc_hd__or2_1
X_11851_ _11851_/A _11851_/B vssd1 vssd1 vccd1 vccd1 _11853_/C sky130_fd_sc_hd__xor2_2
X_10802_ _07472_/Y fanout8/X fanout4/X _07455_/Y vssd1 vssd1 vccd1 vccd1 _10803_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11045__A2_N fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11782_ _11774_/A _12793_/A2 _11586_/B _06902_/A _11781_/Y vssd1 vssd1 vccd1 vccd1
+ _11782_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_28_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10733_ _06977_/Y _10590_/A _10590_/B _06979_/B vssd1 vssd1 vccd1 vccd1 _10734_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_67_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13521_ hold296/X _13555_/A2 _13520_/X _13542_/B2 vssd1 vssd1 vccd1 vccd1 _13522_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07869__B _11731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10576__A _10857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13452_ fanout2/X _13452_/B vssd1 vssd1 vccd1 vccd1 _13452_/Y sky130_fd_sc_hd__nand2_1
X_10664_ _10664_/A _10664_/B vssd1 vssd1 vccd1 vccd1 _10665_/B sky130_fd_sc_hd__or2_1
XFILLER_0_36_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12403_ _12760_/A1 _12389_/X _12402_/Y _12383_/X vssd1 vssd1 vccd1 vccd1 _12403_/X
+ sky130_fd_sc_hd__a211o_1
X_13383_ _13383_/A hold150/X vssd1 vssd1 vccd1 vccd1 _13673_/D sky130_fd_sc_hd__and2_1
XANTENNA__12600__C1 _12971_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10595_ _10595_/A vssd1 vssd1 vccd1 vccd1 _10595_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_105_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12334_ _12334_/A _12334_/B _12334_/C vssd1 vssd1 vccd1 vccd1 _12335_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_23_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12265_ _12764_/B _12265_/B vssd1 vssd1 vccd1 vccd1 _12272_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11706__A1 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11706__B2 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11216_ _11217_/A _11217_/B vssd1 vssd1 vccd1 vccd1 _11340_/A sky130_fd_sc_hd__nand2_1
X_12196_ _12197_/A _12197_/B vssd1 vssd1 vccd1 vccd1 _12286_/A sky130_fd_sc_hd__or2_1
XANTENNA__08583__B1 _09173_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11147_ curr_PC[11] _11265_/C vssd1 vssd1 vccd1 vccd1 _11382_/C sky130_fd_sc_hd__and2_1
XFILLER_0_101_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11078_ _11078_/A _11078_/B vssd1 vssd1 vccd1 vccd1 _11079_/B sky130_fd_sc_hd__or2_1
XANTENNA__08335__B1 _08486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10029_ hold226/A _11693_/A2 _10027_/X _12533_/B1 vssd1 vssd1 vccd1 vccd1 _10029_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__07689__A2 _08866_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06897__B1 _06906_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10693__A1 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10693__B2 _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13719_ _13719_/CLK _13719_/D vssd1 vssd1 vccd1 vccd1 hold300/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07240_ _07240_/A _07240_/B vssd1 vssd1 vccd1 vccd1 _07240_/X sky130_fd_sc_hd__or2_2
XFILLER_0_27_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07171_ _08203_/A _07172_/B vssd1 vssd1 vccd1 vccd1 _07200_/A sky130_fd_sc_hd__or2_1
XFILLER_0_54_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07795__A _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09486__S _09493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07613__A2 _10235_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09812_ _09812_/A _09812_/B vssd1 vssd1 vccd1 vccd1 _09815_/A sky130_fd_sc_hd__or2_1
XFILLER_0_94_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10920__A2 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09743_ _09571_/Y _09579_/B _09578_/A vssd1 vssd1 vccd1 vccd1 _09745_/B sky130_fd_sc_hd__o21a_1
X_06955_ reg1_val[10] _07456_/A vssd1 vssd1 vccd1 vccd1 _06955_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08326__B1 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout281_A _13444_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06858__B _13015_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09674_ _09460_/X _09462_/X _09674_/S vssd1 vssd1 vccd1 vccd1 _09674_/X sky130_fd_sc_hd__mux2_1
X_06886_ _06886_/A _12995_/B vssd1 vssd1 vccd1 vccd1 _06886_/Y sky130_fd_sc_hd__nor2_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08625_ _10236_/A _08625_/B vssd1 vssd1 vccd1 vccd1 _08685_/A sky130_fd_sc_hd__xnor2_2
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06888__B1 _06980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12876__A _13036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ _08556_/A _08556_/B vssd1 vssd1 vccd1 vccd1 _08557_/B sky130_fd_sc_hd__nand2_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09826__B1 _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07507_ reg1_val[13] _07572_/S vssd1 vssd1 vccd1 vccd1 _07517_/A sky130_fd_sc_hd__nor2_1
X_08487_ _09940_/A _08553_/A _08553_/B vssd1 vssd1 vccd1 vccd1 _08498_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_119_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07438_ _07445_/A _07445_/B vssd1 vssd1 vccd1 vccd1 _07438_/X sky130_fd_sc_hd__and2_1
XFILLER_0_107_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13386__B1 _13444_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07369_ _08866_/A2 fanout39/X _07366_/X _08118_/B vssd1 vssd1 vccd1 vccd1 _07370_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_91_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09108_ _09108_/A _09108_/B vssd1 vssd1 vccd1 vccd1 _09110_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07604__A2 _10235_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10380_ _10380_/A _10380_/B vssd1 vssd1 vccd1 vccd1 _10382_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09039_ _09039_/A _09039_/B vssd1 vssd1 vccd1 vccd1 _11461_/A sky130_fd_sc_hd__or2_1
XFILLER_0_20_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12050_ _12050_/A _12050_/B vssd1 vssd1 vccd1 vccd1 _12052_/A sky130_fd_sc_hd__nand2_1
X_11001_ _10313_/Y _11000_/X _11576_/A vssd1 vssd1 vccd1 vccd1 _11001_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11164__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11955__A _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10372__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12649__C1 _09529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08317__B1 _08778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08868__A1 _08907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12952_ _12952_/A vssd1 vssd1 vccd1 vccd1 _12961_/C sky130_fd_sc_hd__inv_2
XANTENNA__08868__B2 _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11903_ _12421_/A _11903_/B vssd1 vssd1 vccd1 vccd1 _11905_/B sky130_fd_sc_hd__xnor2_1
X_12883_ _13042_/B _12883_/B vssd1 vssd1 vccd1 vccd1 _12884_/B sky130_fd_sc_hd__or2_1
XANTENNA__07540__A1 _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11834_ _11727_/A _11727_/B _11739_/A vssd1 vssd1 vccd1 vccd1 _11845_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12416__A2 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09160__A _12668_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11765_ _10860_/B _11343_/Y _11763_/Y _11764_/Y vssd1 vssd1 vccd1 vccd1 _11766_/B
+ sky130_fd_sc_hd__o31ai_4
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10716_ _10717_/A _10717_/B vssd1 vssd1 vccd1 vccd1 _10852_/A sky130_fd_sc_hd__nand2_1
X_13504_ _13504_/A _13504_/B vssd1 vssd1 vccd1 vccd1 _13504_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11696_ _11696_/A _11696_/B _11696_/C _11696_/D vssd1 vssd1 vccd1 vccd1 _11696_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_24_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10647_ _10538_/A _07891_/X fanout10/X _07577_/X vssd1 vssd1 vccd1 vccd1 _10648_/B
+ sky130_fd_sc_hd__o22a_1
X_13435_ _07393_/X _13598_/C hold110/X vssd1 vssd1 vccd1 vccd1 _13699_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_3_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13366_ hold205/X _13542_/B2 _13550_/A2 hold216/X vssd1 vssd1 vccd1 vccd1 hold230/A
+ sky130_fd_sc_hd__a22o_1
X_10578_ _09988_/X _09989_/X _10579_/C vssd1 vssd1 vccd1 vccd1 _10578_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_11_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06915__A_N _07544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12317_ _07230_/A _12799_/A2 _11688_/B reg1_val[23] vssd1 vssd1 vccd1 vccd1 _12317_/X
+ sky130_fd_sc_hd__o22a_1
X_13297_ _13513_/B _13514_/A _13253_/X vssd1 vssd1 vccd1 vccd1 _13519_/A sky130_fd_sc_hd__a21o_1
X_12248_ fanout15/X _09145_/Y fanout7/X fanout31/X vssd1 vssd1 vccd1 vccd1 _12249_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11155__A2 _07891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12179_ _12180_/A _12180_/B vssd1 vssd1 vccd1 vccd1 _12258_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10902__A2 _07543_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09335__A _12092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11863__B1 _11955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08410_ _08466_/A _08466_/B _08369_/X vssd1 vssd1 vccd1 vccd1 _08471_/A sky130_fd_sc_hd__a21oi_2
X_09390_ _09390_/A _09390_/B vssd1 vssd1 vccd1 vccd1 _09408_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_59_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08341_ _08337_/X _08341_/B vssd1 vssd1 vccd1 vccd1 _08406_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_80_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08272_ _09659_/B _08272_/B _08272_/C vssd1 vssd1 vccd1 vccd1 _08274_/B sky130_fd_sc_hd__and3_1
XFILLER_0_73_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07223_ _07223_/A _07224_/B vssd1 vssd1 vccd1 vccd1 _07223_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_15_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10944__A _10944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12040__B1 _12164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07154_ _12578_/A _12778_/A vssd1 vssd1 vccd1 vccd1 _12056_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_6_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07598__A1 _08907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07598__B2 _08328_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07085_ _12740_/A _07084_/X _07060_/Y vssd1 vssd1 vccd1 vccd1 _07085_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13466__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout113 _07491_/X vssd1 vssd1 vccd1 vccd1 _10522_/A sky130_fd_sc_hd__buf_8
Xfanout124 _07366_/X vssd1 vssd1 vccd1 vccd1 _09216_/B2 sky130_fd_sc_hd__buf_6
Xfanout135 _12056_/B vssd1 vssd1 vccd1 vccd1 _12742_/A sky130_fd_sc_hd__buf_4
XANTENNA__10354__B1 _10538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout146 _08746_/A vssd1 vssd1 vccd1 vccd1 _09575_/A sky130_fd_sc_hd__buf_12
XANTENNA__09245__A _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout157 _07240_/X vssd1 vssd1 vccd1 vccd1 _08950_/B sky130_fd_sc_hd__clkbuf_8
Xfanout168 _09435_/X vssd1 vssd1 vccd1 vccd1 _09493_/S sky130_fd_sc_hd__clkbuf_8
X_07987_ _09371_/A _07987_/B vssd1 vssd1 vccd1 vccd1 _08071_/A sky130_fd_sc_hd__xnor2_4
Xfanout179 _09373_/A vssd1 vssd1 vccd1 vccd1 _10239_/A sky130_fd_sc_hd__buf_12
X_09726_ _09726_/A _09726_/B vssd1 vssd1 vccd1 vccd1 _09740_/A sky130_fd_sc_hd__nand2_2
X_06938_ reg2_val[12] _06980_/B _06936_/X vssd1 vssd1 vccd1 vccd1 _07476_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__10106__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10657__A1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09657_ _12742_/A _09656_/B _09656_/C vssd1 vssd1 vccd1 vccd1 _09658_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__10657__B2 fanout31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06869_ _06869_/A _06869_/B vssd1 vssd1 vccd1 vccd1 _12046_/A sky130_fd_sc_hd__nor2_2
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ _08608_/A _08608_/B vssd1 vssd1 vccd1 vccd1 _08609_/B sky130_fd_sc_hd__nand2_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ _09588_/A _09753_/A _09588_/C vssd1 vssd1 vccd1 vccd1 _09753_/B sky130_fd_sc_hd__nand3_2
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _08891_/B _10049_/A2 _09885_/B1 _08873_/A2 vssd1 vssd1 vccd1 vccd1 _08540_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07286__B1 _07201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11550_ _11551_/A _11551_/B _11551_/C vssd1 vssd1 vccd1 vccd1 _11550_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_9_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10501_ fanout46/X fanout84/X _08580_/B fanout49/X vssd1 vssd1 vccd1 vccd1 _10502_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_80_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11481_ _07094_/B _09509_/X _11587_/A2 _06927_/B _11480_/X vssd1 vssd1 vccd1 vccd1
+ _11481_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_0_107_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13220_ hold46/X hold278/A vssd1 vssd1 vccd1 vccd1 _13222_/A sky130_fd_sc_hd__and2b_1
X_10432_ _10432_/A _10432_/B vssd1 vssd1 vccd1 vccd1 _10981_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_33_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07589__A1 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07589__B2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11385__A2 _11600_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13151_ _13151_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13151_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_0_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10363_ _10363_/A _10363_/B vssd1 vssd1 vccd1 vccd1 _10371_/A sky130_fd_sc_hd__xnor2_4
X_12102_ _12011_/A _12011_/B _12009_/Y vssd1 vssd1 vccd1 vccd1 _12105_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13082_ _13082_/A _13082_/B vssd1 vssd1 vccd1 vccd1 _13084_/C sky130_fd_sc_hd__nand2_2
X_10294_ _10296_/A _10296_/B vssd1 vssd1 vccd1 vccd1 _10294_/X sky130_fd_sc_hd__or2_1
X_12033_ _12031_/X _12033_/B vssd1 vssd1 vccd1 vccd1 _12207_/A sky130_fd_sc_hd__and2b_2
XFILLER_0_18_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10896__B2 _09839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12935_ _12956_/A _12935_/B vssd1 vssd1 vccd1 vccd1 _12936_/B sky130_fd_sc_hd__or2_1
XFILLER_0_125_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12866_ _12872_/B _12866_/B vssd1 vssd1 vccd1 vccd1 new_PC[9] sky130_fd_sc_hd__and2_4
XANTENNA__10748__B _12056_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07403__A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11817_ _11929_/A _11817_/B vssd1 vssd1 vccd1 vccd1 _11819_/B sky130_fd_sc_hd__or2_1
XFILLER_0_55_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ _09529_/B _12783_/X _12796_/X _12781_/Y vssd1 vssd1 vccd1 vccd1 _12797_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11073__A1 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11073__B2 _08580_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ _11749_/A _11749_/B vssd1 vssd1 vccd1 vccd1 _11849_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_56_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10764__A _12825_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11679_ reg1_val[16] curr_PC[16] vssd1 vssd1 vccd1 vccd1 _11679_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13418_ _13690_/Q _13142_/A _13444_/B1 hold151/X _13383_/A vssd1 vssd1 vccd1 vccd1
+ hold152/A sky130_fd_sc_hd__o221a_1
XFILLER_0_107_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13349_ _13359_/A hold196/X vssd1 vssd1 vccd1 vccd1 _13656_/D sky130_fd_sc_hd__and2_1
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10584__B1 _10730_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08529__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07910_ _07911_/A _07911_/B vssd1 vssd1 vccd1 vccd1 _07910_/Y sky130_fd_sc_hd__nor2_1
X_08890_ _08889_/A _08889_/C _08889_/B vssd1 vssd1 vccd1 vccd1 _08896_/B sky130_fd_sc_hd__a21oi_1
X_07841_ _07841_/A _07841_/B vssd1 vssd1 vccd1 vccd1 _07848_/B sky130_fd_sc_hd__xor2_2
XANTENNA__07752__A1 _10049_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07752__B2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07772_ _07772_/A _07772_/B _07815_/A vssd1 vssd1 vccd1 vccd1 _07774_/B sky130_fd_sc_hd__and3_1
XANTENNA__12089__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09511_ _13748_/A _13744_/A instruction[5] instruction[3] vssd1 vssd1 vccd1 vccd1
+ _09511_/X sky130_fd_sc_hd__and4b_1
X_09442_ _09440_/X _09441_/X _09688_/S vssd1 vssd1 vccd1 vccd1 _09442_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09373_ _09373_/A _09373_/B vssd1 vssd1 vccd1 vccd1 _09376_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_59_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09257__A1 _08271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09257__B2 _12982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout244_A _12782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08324_ _08322_/A _08322_/B _08402_/A vssd1 vssd1 vccd1 vccd1 _08343_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_46_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08255_ _08255_/A _08255_/B vssd1 vssd1 vccd1 vccd1 _08256_/B sky130_fd_sc_hd__or2_1
XFILLER_0_117_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10674__A _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06871__B _13010_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07206_ _10239_/A _07206_/B vssd1 vssd1 vccd1 vccd1 _07245_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08186_ _08186_/A _08186_/B vssd1 vssd1 vccd1 vccd1 _08286_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10024__C1 _10734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07137_ instruction[5] _09516_/B vssd1 vssd1 vccd1 vccd1 _07137_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_15_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09674__S _09674_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07068_ _06849_/C _07067_/X _12578_/B vssd1 vssd1 vccd1 vccd1 _07068_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_30_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10327__B1 _12796_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07207__B _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09709_ _10007_/S _11793_/B _09706_/Y _09707_/X _09708_/X vssd1 vssd1 vccd1 vccd1
+ _09709_/X sky130_fd_sc_hd__o221a_1
XANTENNA__09703__A _12515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10981_ _10981_/A _10981_/B _10981_/C _11106_/A vssd1 vssd1 vccd1 vccd1 _10981_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12720_ fanout10/X _12666_/A _12718_/Y _12769_/S vssd1 vssd1 vccd1 vccd1 _12723_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_97_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12651_ _12735_/A1 _12705_/B hold219/A vssd1 vssd1 vccd1 vccd1 _12651_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11602_ fanout50/X fanout38/X fanout36/X _12557_/A vssd1 vssd1 vccd1 vccd1 _11603_/B
+ sky130_fd_sc_hd__o22a_1
X_12582_ _12581_/A _12581_/B _12581_/Y _09506_/X vssd1 vssd1 vccd1 vccd1 _12582_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10802__A1 _07472_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10802__B2 _07455_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11533_ _11533_/A _11533_/B vssd1 vssd1 vccd1 vccd1 _11546_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_92_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13598__C _13598_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11464_ _11463_/A _06931_/Y _07043_/X _11463_/Y vssd1 vssd1 vccd1 vccd1 _11465_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_61_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10415_ _10415_/A _10415_/B vssd1 vssd1 vccd1 vccd1 _10428_/A sky130_fd_sc_hd__xor2_4
X_13203_ hold30/X _13207_/B vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__or2_1
X_11395_ _12268_/A fanout38/X fanout36/X fanout46/X vssd1 vssd1 vccd1 vccd1 _11396_/B
+ sky130_fd_sc_hd__o22a_1
X_13134_ _13131_/A _13133_/B _13131_/B vssd1 vssd1 vccd1 vccd1 _13135_/B sky130_fd_sc_hd__a21boi_2
X_10346_ _10288_/A _10288_/B _10289_/Y vssd1 vssd1 vccd1 vccd1 _10429_/A sky130_fd_sc_hd__a21bo_2
XANTENNA__10030__A2 _12793_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ _13065_/A _13065_/B vssd1 vssd1 vccd1 vccd1 _13068_/A sky130_fd_sc_hd__or2_2
X_10277_ _10277_/A _10277_/B vssd1 vssd1 vccd1 vccd1 _10278_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_29_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10750__C _12235_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12016_ _12016_/A _12016_/B vssd1 vssd1 vccd1 vccd1 _12019_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10869__A1 _10734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07195__C1 _06875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11862__B _12163_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13659_/CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA__10097__A2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13135__A _13135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11294__A1 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12918_ reg1_val[18] curr_PC[18] _12978_/S vssd1 vssd1 vccd1 vccd1 _12920_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_88_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11294__B2 _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12849_ _12858_/A _12849_/B vssd1 vssd1 vccd1 vccd1 _12851_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_28_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13440__C1 _13568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12794__A1 _09839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08040_ _08040_/A _08040_/B vssd1 vssd1 vccd1 vccd1 _08043_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09991_ _10577_/A _09991_/B vssd1 vssd1 vccd1 vccd1 _10726_/C sky130_fd_sc_hd__xor2_4
XANTENNA__07973__A1 _10235_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07973__B2 _08873_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08942_ _09659_/B _08942_/B vssd1 vssd1 vccd1 vccd1 _08959_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10309__B1 _10734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09507__B _13748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13029__B _13029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08873_ _09674_/S _08873_/A2 _08891_/B _08873_/B2 vssd1 vssd1 vccd1 vccd1 _08874_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07725__A1 _09173_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07725__B2 _07471_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07824_ _10266_/A _07824_/B vssd1 vssd1 vccd1 vccd1 _07828_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07027__B _07110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07755_ _08395_/B _10522_/A _07557_/Y fanout28/X vssd1 vssd1 vccd1 vccd1 _07756_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07489__B1 _07476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10088__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07686_ _07686_/A _07686_/B vssd1 vssd1 vccd1 vccd1 _07710_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08139__A _10078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09425_ _09426_/A _09426_/B vssd1 vssd1 vccd1 vccd1 _09989_/A sky130_fd_sc_hd__and2_1
XFILLER_0_19_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09356_ _09357_/A _09357_/B vssd1 vssd1 vccd1 vccd1 _09358_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08307_ _08857_/A _08307_/B vssd1 vssd1 vccd1 vccd1 _08377_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_90_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09287_ _09346_/A _09287_/B vssd1 vssd1 vccd1 vccd1 _09289_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_35_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08238_ _08236_/X _08993_/A vssd1 vssd1 vccd1 vccd1 _09003_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_50_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12537__B2 _12537_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08169_ _08169_/A _08169_/B vssd1 vssd1 vccd1 vccd1 _08232_/B sky130_fd_sc_hd__xor2_1
X_10200_ _10200_/A _10200_/B vssd1 vssd1 vccd1 vccd1 _10344_/A sky130_fd_sc_hd__nand2_1
X_11180_ _12094_/A _11180_/B vssd1 vssd1 vccd1 vccd1 _11182_/B sky130_fd_sc_hd__xnor2_2
X_10131_ _10131_/A _10131_/B vssd1 vssd1 vccd1 vccd1 _10144_/A sky130_fd_sc_hd__xor2_4
XANTENNA__07218__A _12982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10062_ _10063_/A _10063_/B vssd1 vssd1 vccd1 vccd1 _10282_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_100_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11276__A1 _07310_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09152__B _09153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11276__B2 _07282_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10964_ _10964_/A _10964_/B vssd1 vssd1 vccd1 vccd1 _10966_/B sky130_fd_sc_hd__and2_1
XANTENNA__08049__A _09575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12703_ _12786_/B1 _12746_/B hold299/A vssd1 vssd1 vccd1 vccd1 _12703_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13683_ _13701_/CLK hold21/X vssd1 vssd1 vccd1 vccd1 hold157/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10895_ _12225_/B vssd1 vssd1 vccd1 vccd1 _10895_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07888__A _10239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12634_ _12635_/B _12635_/C vssd1 vssd1 vccd1 vccd1 _12634_/X sky130_fd_sc_hd__or2_1
XANTENNA__06792__A _13135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12776__A1 _13129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12565_ _12565_/A _12565_/B _12565_/C vssd1 vssd1 vccd1 vccd1 _12566_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_80_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11516_ _11516_/A _11516_/B vssd1 vssd1 vccd1 vccd1 _11520_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_41_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12496_ _12496_/A _12666_/A vssd1 vssd1 vccd1 vccd1 _12497_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_34_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11447_ _11447_/A _11447_/B vssd1 vssd1 vccd1 vccd1 _11449_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11378_ _11367_/Y _11368_/X _11377_/Y _09493_/S _11376_/X vssd1 vssd1 vccd1 vccd1
+ _11378_/Y sky130_fd_sc_hd__o221ai_2
XFILLER_0_21_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13117_ _13117_/A _13121_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[27] sky130_fd_sc_hd__xnor2_4
X_10329_ _07180_/C _11793_/B _10326_/Y _10327_/X _10328_/X vssd1 vssd1 vccd1 vccd1
+ _10329_/X sky130_fd_sc_hd__o221a_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ reg1_val[13] _13048_/B vssd1 vssd1 vccd1 vccd1 _13057_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_56_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08904__B1 _07420_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10489__A _12093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06930__A2 _06980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11267__A1 _12867_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07540_ _10507_/A _11157_/A _07538_/X vssd1 vssd1 vccd1 vccd1 _10787_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07471_ _07471_/A _07472_/B vssd1 vssd1 vccd1 vccd1 _07471_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__09880__A1 _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09210_ _09195_/A _09195_/B _09196_/Y vssd1 vssd1 vccd1 vccd1 _09311_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__09489__S _09493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10490__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09141_ _09951_/A _09141_/B vssd1 vssd1 vccd1 vccd1 _09151_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_8_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11113__A _11342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09072_ _09071_/B _09079_/A _09077_/B vssd1 vssd1 vccd1 vccd1 _09073_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_44_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10242__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08023_ _07817_/A _07817_/C _07817_/B vssd1 vssd1 vccd1 vccd1 _08024_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout4 fanout4/A vssd1 vssd1 vccd1 vccd1 fanout4/X sky130_fd_sc_hd__buf_8
XANTENNA__09396__B1 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13192__A1 _07230_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09974_ _09974_/A _09974_/B vssd1 vssd1 vccd1 vccd1 _09975_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08925_ _08931_/A _08931_/B vssd1 vssd1 vccd1 vccd1 _08926_/A sky130_fd_sc_hd__nand2b_1
X_08856_ _08887_/A _08887_/B vssd1 vssd1 vccd1 vccd1 _08864_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09253__A _10239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07807_ _07807_/A _07807_/B vssd1 vssd1 vccd1 vccd1 _08008_/B sky130_fd_sc_hd__xnor2_1
X_08787_ _08788_/A _08788_/B vssd1 vssd1 vccd1 vccd1 _09044_/C sky130_fd_sc_hd__or2_2
XANTENNA__06921__A2 _06936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11258__A1 _09521_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07738_ _10239_/A _07738_/B vssd1 vssd1 vccd1 vccd1 _07741_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12455__B1 _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07669_ _07749_/B vssd1 vssd1 vccd1 vccd1 _07669_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12818__S _12825_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09408_ _09408_/A _09408_/B vssd1 vssd1 vccd1 vccd1 _09409_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_48_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10680_ _10838_/A _10680_/B vssd1 vssd1 vccd1 vccd1 _10682_/B sky130_fd_sc_hd__or2_1
XANTENNA_fanout22_A fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09339_ _09228_/A _09228_/B _09229_/Y vssd1 vssd1 vccd1 vccd1 _09340_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_62_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10769__B1 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12350_ _12351_/A _12351_/B _12351_/C vssd1 vssd1 vccd1 vccd1 _12352_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_22_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11301_ _11301_/A _11301_/B vssd1 vssd1 vccd1 vccd1 _11302_/C sky130_fd_sc_hd__xor2_2
X_12281_ _12362_/A _12281_/B vssd1 vssd1 vccd1 vccd1 _12283_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_15_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11232_ _11117_/B _11118_/A _11562_/A vssd1 vssd1 vccd1 vccd1 _11233_/B sky130_fd_sc_hd__a21o_1
XANTENNA__09926__A2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08332__A _09371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11163_ _11163_/A _11163_/B vssd1 vssd1 vccd1 vccd1 _11204_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10114_ _09894_/A _09894_/B _09892_/Y vssd1 vssd1 vccd1 vccd1 _10115_/A sky130_fd_sc_hd__o21ai_1
X_11094_ _11095_/A _11095_/B vssd1 vssd1 vccd1 vccd1 _11153_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__13486__A2 _13555_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10045_ _12742_/A _10200_/A vssd1 vssd1 vccd1 vccd1 _10045_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09163__A _11731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11996_ _12189_/A fanout8/X fanout3/X _07198_/Y vssd1 vssd1 vccd1 vccd1 _12087_/C
+ sky130_fd_sc_hd__a22o_1
X_13735_ _13735_/CLK _13735_/D vssd1 vssd1 vccd1 vccd1 hold233/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10947_ fanout49/X fanout25/X fanout23/X _12557_/A vssd1 vssd1 vccd1 vccd1 _10948_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_128_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13666_ _13736_/CLK _13666_/D vssd1 vssd1 vccd1 vccd1 hold207/A sky130_fd_sc_hd__dfxtp_1
X_10878_ _10451_/Y _10877_/X _11576_/A vssd1 vssd1 vccd1 vccd1 _10879_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_85_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12617_ _12617_/A fanout7/X vssd1 vssd1 vccd1 vccd1 _12617_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_109_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13597_ _13599_/D _13597_/B vssd1 vssd1 vccd1 vccd1 _13597_/X sky130_fd_sc_hd__and2_1
XFILLER_0_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07625__B1 _08118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11421__A1 wire101/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12548_ _12667_/A fanout8/X fanout3/X _12614_/A vssd1 vssd1 vccd1 vccd1 _12549_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11421__B2 _13180_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_2 _09707_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ _12543_/B _12478_/Y _12971_/S _12476_/X vssd1 vssd1 vccd1 vccd1 dest_val[25]
+ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__10772__A _11281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13174__A1 _13174_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06971_ reg1_val[8] _07184_/D vssd1 vssd1 vccd1 vccd1 _06971_/Y sky130_fd_sc_hd__nor2_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08710_ _09950_/A _08710_/B vssd1 vssd1 vccd1 vccd1 _08744_/B sky130_fd_sc_hd__xnor2_2
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09690_ _09686_/X _09689_/X _10176_/A vssd1 vssd1 vccd1 vccd1 _09690_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_83_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09550__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08641_ _08662_/A _08639_/Y _08629_/Y vssd1 vssd1 vccd1 vccd1 _08650_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_89_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08572_ _09068_/B _09057_/A vssd1 vssd1 vccd1 vccd1 _08572_/Y sky130_fd_sc_hd__nor2_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07523_ _07523_/A _07523_/B vssd1 vssd1 vccd1 vccd1 _11309_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_119_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13323__A _13459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07454_ _07186_/B _07186_/C _07183_/Y _07476_/B vssd1 vssd1 vccd1 vccd1 _07456_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_9_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07321__A _11126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13042__B _13042_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07385_ reg1_val[24] _07634_/B _07634_/C reg1_val[25] vssd1 vssd1 vccd1 vccd1 _07386_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_123_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09124_ fanout42/X fanout68/X fanout66/X fanout40/X vssd1 vssd1 vccd1 vccd1 _09125_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09055_ _09055_/A _09055_/B _09055_/C vssd1 vssd1 vccd1 vccd1 _11864_/D sky130_fd_sc_hd__nand3_2
XFILLER_0_114_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08006_ _08006_/A _08006_/B vssd1 vssd1 vccd1 vccd1 _08044_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11715__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09957_ _10225_/A fanout9/X fanout4/X _10104_/A vssd1 vssd1 vccd1 vccd1 _09958_/B
+ sky130_fd_sc_hd__a22o_1
X_08908_ _09659_/B _08908_/B _08908_/C vssd1 vssd1 vccd1 vccd1 _08910_/B sky130_fd_sc_hd__and3_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _10374_/B2 _07643_/B fanout13/X _10349_/A1 vssd1 vssd1 vccd1 vccd1 _09889_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08839_ _08860_/B _08860_/A vssd1 vssd1 vccd1 vccd1 _08843_/C sky130_fd_sc_hd__and2b_1
X_11850_ _11851_/A _11851_/B vssd1 vssd1 vccd1 vccd1 _11944_/B sky130_fd_sc_hd__nand2b_1
X_10801_ _10801_/A vssd1 vssd1 vccd1 vccd1 _10808_/A sky130_fd_sc_hd__inv_2
XANTENNA__10857__A _10857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11781_ _06902_/B _09516_/X _09525_/Y reg1_val[17] vssd1 vssd1 vccd1 vccd1 _11781_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_0_79_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13520_ hold251/X _13519_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13520_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07855__B1 _11047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10732_ _11562_/A _10731_/B _10731_/C vssd1 vssd1 vccd1 vccd1 _10732_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__08327__A _09373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10576__B _10981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13451_ _13451_/A _13451_/B vssd1 vssd1 vccd1 vccd1 _13452_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10663_ _10664_/A _10664_/B vssd1 vssd1 vccd1 vccd1 _10665_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_82_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12402_ _12391_/Y _12392_/X _12401_/X vssd1 vssd1 vccd1 vccd1 _12402_/Y sky130_fd_sc_hd__o21ai_1
X_10594_ _11472_/S _09496_/X _09534_/C vssd1 vssd1 vccd1 vccd1 _10595_/A sky130_fd_sc_hd__o21ai_2
X_13382_ hold149/X _07118_/B _13207_/B _12982_/A vssd1 vssd1 vccd1 vccd1 hold150/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12600__B1 _12657_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12333_ _12334_/A _12334_/B _12334_/C vssd1 vssd1 vccd1 vccd1 _12335_/A sky130_fd_sc_hd__a21o_1
XANTENNA__13156__A1 _10225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12264_ _12413_/A fanout8/X fanout3/X _12331_/A vssd1 vssd1 vccd1 vccd1 _12265_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08062__A _09949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11706__A2 _07597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11215_ _11215_/A _11215_/B vssd1 vssd1 vccd1 vccd1 _11217_/B sky130_fd_sc_hd__xnor2_1
X_12195_ _12195_/A _12195_/B vssd1 vssd1 vccd1 vccd1 _12197_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08583__A1 _08821_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08583__B2 _08821_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11146_ _11115_/X _11116_/Y _11118_/Y _11866_/A _11145_/X vssd1 vssd1 vccd1 vccd1
+ _11146_/X sky130_fd_sc_hd__a221o_1
X_11077_ _11078_/A _11078_/B vssd1 vssd1 vccd1 vccd1 _11079_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08335__A1 _13149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08335__B2 _08923_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07406__A _10456_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10028_ _10606_/A2 _10027_/X hold226/A vssd1 vssd1 vccd1 vccd1 _10028_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07125__B _07129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10693__A2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11890__A1 _09529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09621__A _10119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10767__A _11151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11979_ _12710_/B2 _11241_/X _11259_/X _12537_/B2 _11978_/X vssd1 vssd1 vccd1 vccd1
+ _11980_/C sky130_fd_sc_hd__a221o_1
XANTENNA__06964__B _10889_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13718_ _13719_/CLK _13718_/D vssd1 vssd1 vccd1 vccd1 hold289/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13649_ _13649_/CLK _13649_/D vssd1 vssd1 vccd1 vccd1 hold163/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12982__A _12982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07170_ _08203_/A _07172_/B vssd1 vssd1 vccd1 vccd1 _10096_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07363__C_N _07398_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09811_ _09811_/A _09811_/B vssd1 vssd1 vccd1 vccd1 _09816_/A sky130_fd_sc_hd__or2_2
XANTENNA__09771__B1 _08704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09742_ _09627_/A _09626_/B _09624_/X vssd1 vssd1 vccd1 vccd1 _09745_/A sky130_fd_sc_hd__a21oi_2
X_06954_ _06928_/A _06936_/B _13036_/B _06952_/X vssd1 vssd1 vccd1 vccd1 _07456_/A
+ sky130_fd_sc_hd__a31oi_4
XFILLER_0_94_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08326__A1 _08821_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08326__B2 _08821_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ _09456_/X _09459_/X _09674_/S vssd1 vssd1 vccd1 vccd1 _09673_/X sky130_fd_sc_hd__mux2_1
X_06885_ instruction[28] _12981_/C vssd1 vssd1 vccd1 vccd1 _12995_/B sky130_fd_sc_hd__and2_4
XANTENNA_fanout274_A _13444_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _08891_/B _10522_/A _08868_/B1 _08873_/A2 vssd1 vssd1 vccd1 vccd1 _08625_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ _08555_/A _08555_/B vssd1 vssd1 vccd1 vccd1 _08620_/A sky130_fd_sc_hd__xor2_1
XANTENNA__09826__B2 _09650_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06874__B _07201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07506_ _07506_/A _07506_/B vssd1 vssd1 vccd1 vccd1 _07651_/A sky130_fd_sc_hd__xor2_4
X_08486_ _09671_/S _08486_/B vssd1 vssd1 vccd1 vccd1 _08553_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08147__A _09591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07437_ _07435_/X _07436_/Y _07637_/B vssd1 vssd1 vccd1 vccd1 _07445_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_18_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_13_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13735_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07368_ _12177_/A _07368_/B vssd1 vssd1 vccd1 vccd1 _07368_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_32_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11397__B1 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09107_ _10050_/A _09107_/B vssd1 vssd1 vccd1 vccd1 _09108_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07299_ _11793_/A _07300_/B vssd1 vssd1 vccd1 vccd1 _07299_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_115_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09038_ _09044_/B _09044_/C _09044_/D vssd1 vssd1 vccd1 vccd1 _09039_/B sky130_fd_sc_hd__and3_1
XFILLER_0_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11149__B1 _12825_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11000_ _09845_/X _09849_/X _11575_/S vssd1 vssd1 vccd1 vccd1 _11000_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10372__A1 _07455_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10372__B2 wire122/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09425__B _09426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08317__A1 _09885_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08317__B2 _10049_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07226__A _09950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12951_ _12951_/A _12951_/B vssd1 vssd1 vccd1 vccd1 _12952_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08868__A2 _09216_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11902_ _12557_/A _07416_/X _07422_/Y _12557_/B vssd1 vssd1 vccd1 vccd1 _11903_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_99_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12882_ _13042_/B _12883_/B vssd1 vssd1 vccd1 vccd1 _12893_/A sky130_fd_sc_hd__nand2_1
X_11833_ _11833_/A _11833_/B vssd1 vssd1 vccd1 vccd1 _11847_/A sky130_fd_sc_hd__and2_1
XFILLER_0_68_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _11345_/X _11763_/A _11950_/A _11762_/X vssd1 vssd1 vccd1 vccd1 _11764_/Y
+ sky130_fd_sc_hd__a31oi_2
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08057__A _10119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13503_ _13257_/X _13503_/B vssd1 vssd1 vccd1 vccd1 _13504_/B sky130_fd_sc_hd__nand2b_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _10715_/A _10715_/B vssd1 vssd1 vccd1 vccd1 _10717_/B sky130_fd_sc_hd__xnor2_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11695_ _09493_/S _11577_/Y _11694_/X vssd1 vssd1 vccd1 vccd1 _11696_/D sky130_fd_sc_hd__o21ai_1
XFILLER_0_126_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13434_ hold95/X _13142_/A _13444_/B1 hold53/X _13568_/A vssd1 vssd1 vccd1 vccd1
+ hold110/A sky130_fd_sc_hd__o221a_1
XFILLER_0_24_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10646_ _10544_/A _10544_/C _10544_/B vssd1 vssd1 vccd1 vccd1 _10654_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_70_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13365_ _13543_/A hold206/X vssd1 vssd1 vccd1 vccd1 _13664_/D sky130_fd_sc_hd__and2_1
XFILLER_0_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10577_ _10577_/A _10631_/A _10857_/A _10981_/A vssd1 vssd1 vccd1 vccd1 _10579_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_0_51_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09450__C1 _10456_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12316_ hold282/A _12314_/X _12315_/Y vssd1 vssd1 vccd1 vccd1 _12316_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13296_ _13508_/B _13509_/A _13255_/X vssd1 vssd1 vccd1 vccd1 _13514_/A sky130_fd_sc_hd__a21o_1
X_12247_ _12165_/Y _12372_/C _11231_/A vssd1 vssd1 vccd1 vccd1 _12296_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_121_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12178_ _07361_/Y fanout7/X _12177_/X _12253_/A vssd1 vssd1 vccd1 vccd1 _12180_/B
+ sky130_fd_sc_hd__a22o_1
X_11129_ _12648_/A _11129_/B vssd1 vssd1 vccd1 vccd1 _11129_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09351__A _10078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08340_ _08340_/A _08340_/B vssd1 vssd1 vccd1 vccd1 _08341_/B sky130_fd_sc_hd__or2_2
XFILLER_0_80_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11615__A1 _11708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08271_ _08271_/A wire101/A vssd1 vssd1 vccd1 vccd1 _08272_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08492__B1 _08704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07222_ _07221_/A _07213_/A _07213_/B _07521_/A vssd1 vssd1 vccd1 vccd1 _07224_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_0_27_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07153_ _12578_/A _12778_/A vssd1 vssd1 vccd1 vccd1 _07153_/X sky130_fd_sc_hd__and2_1
XANTENNA__08244__B1 _08486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12040__A1 _12695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07598__A2 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09992__B1 _10726_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07084_ _12693_/A _07083_/Y _07061_/Y vssd1 vssd1 vccd1 vccd1 _07084_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_2_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout103 _07299_/Y vssd1 vssd1 vccd1 vccd1 _11732_/A sky130_fd_sc_hd__buf_8
Xfanout125 _07347_/X vssd1 vssd1 vccd1 vccd1 _08866_/A2 sky130_fd_sc_hd__buf_6
XANTENNA__08430__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout136 _11231_/A vssd1 vssd1 vccd1 vccd1 _11864_/A sky130_fd_sc_hd__buf_4
XANTENNA__10354__B2 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout147 _07532_/Y vssd1 vssd1 vccd1 vccd1 _08746_/A sky130_fd_sc_hd__clkbuf_16
Xfanout158 _07200_/Y vssd1 vssd1 vccd1 vccd1 _08821_/A1 sky130_fd_sc_hd__buf_6
X_07986_ fanout56/X _07240_/X fanout40/X _08866_/B2 vssd1 vssd1 vccd1 vccd1 _07987_/B
+ sky130_fd_sc_hd__o22a_2
Xfanout169 _09435_/X vssd1 vssd1 vccd1 vccd1 _09839_/A sky130_fd_sc_hd__clkbuf_4
X_09725_ _09644_/A _09644_/B _09645_/Y vssd1 vssd1 vccd1 vccd1 _09822_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__10106__A1 _10349_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06937_ reg2_val[12] _06980_/B _06936_/X vssd1 vssd1 vccd1 vccd1 _07188_/B sky130_fd_sc_hd__a21o_1
XANTENNA__10106__B2 _10225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09656_ _12742_/A _09656_/B _09656_/C vssd1 vssd1 vccd1 vccd1 _09658_/B sky130_fd_sc_hd__or3_1
XANTENNA__10657__A2 _11527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06868_ _07483_/A _07201_/A vssd1 vssd1 vccd1 vccd1 _06869_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_97_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08607_ _08607_/A _08607_/B vssd1 vssd1 vccd1 vccd1 _08608_/B sky130_fd_sc_hd__or2_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ _09586_/B _09586_/C _09779_/A vssd1 vssd1 vccd1 vccd1 _09588_/C sky130_fd_sc_hd__a21o_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06799_ reg1_val[27] _07252_/A vssd1 vssd1 vccd1 vccd1 _06802_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_49_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _08746_/A _08538_/B vssd1 vssd1 vccd1 vccd1 _08544_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07286__A1 _07521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08469_ _08470_/A _08470_/B vssd1 vssd1 vccd1 vccd1 _08469_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_37_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10500_ _10500_/A _10500_/B vssd1 vssd1 vccd1 vccd1 _10557_/A sky130_fd_sc_hd__xnor2_4
X_11480_ _07526_/A _12799_/A2 _12657_/B1 reg1_val[14] _11479_/Y vssd1 vssd1 vccd1
+ vccd1 _11480_/X sky130_fd_sc_hd__o221a_1
X_10431_ _10432_/A _10432_/B vssd1 vssd1 vccd1 vccd1 _10431_/X sky130_fd_sc_hd__and2_1
XFILLER_0_123_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07589__A2 _08866_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10042__B1 _12825_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13150_ hold9/X _13193_/B _13149_/Y _13459_/A vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__o211a_1
X_10362_ _10363_/A _10363_/B vssd1 vssd1 vccd1 vccd1 _10362_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12101_ _12012_/A _12012_/B _12001_/A vssd1 vssd1 vccd1 vccd1 _12112_/A sky130_fd_sc_hd__o21a_1
X_13081_ _13081_/A _13081_/B _13081_/C _13081_/D vssd1 vssd1 vccd1 vccd1 _13084_/B
+ sky130_fd_sc_hd__or4_2
X_10293_ _10293_/A _10293_/B vssd1 vssd1 vccd1 vccd1 _10296_/B sky130_fd_sc_hd__xnor2_4
X_12032_ _12032_/A _12032_/B _12032_/C vssd1 vssd1 vccd1 vccd1 _12033_/B sky130_fd_sc_hd__or3_1
Xhold190 hold190/A vssd1 vssd1 vccd1 vccd1 hold190/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07210__A1 _09694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09155__B _13129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12934_ _12956_/A _12935_/B vssd1 vssd1 vccd1 vccd1 _12936_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_125_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12865_ _12865_/A _12865_/B _12865_/C vssd1 vssd1 vccd1 vccd1 _12866_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_96_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11816_ _11816_/A _11816_/B vssd1 vssd1 vccd1 vccd1 _11817_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _12796_/A1 _12787_/Y _12795_/X vssd1 vssd1 vccd1 vccd1 _12796_/X sky130_fd_sc_hd__o21a_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07277__A1 _10542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11073__A2 _07597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _11648_/A _11647_/B _11647_/A vssd1 vssd1 vccd1 vccd1 _11749_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_126_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11678_ _11574_/A _11574_/B _11572_/B vssd1 vssd1 vccd1 vccd1 _11682_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_114_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_718 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13417_ _11709_/A _13419_/A2 hold23/X vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__o21a_1
XANTENNA__13140__B _13584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10629_ _10981_/A _10981_/B vssd1 vssd1 vccd1 vccd1 _10629_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_113_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10033__B1 _12796_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13348_ hold193/X _13506_/B2 _13506_/A2 hold195/X vssd1 vssd1 vccd1 vccd1 hold196/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13279_ hold9/X hold262/X vssd1 vssd1 vccd1 vccd1 _13279_/X sky130_fd_sc_hd__and2b_1
XANTENNA__08529__A1 _08907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08529__B2 _08197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08250__A _10263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10336__A1 _12525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07840_ _07838_/A _07838_/B _07969_/A vssd1 vssd1 vccd1 vccd1 _07848_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__07752__A2 _08486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12089__A1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07771_ _07770_/A _07813_/A vssd1 vssd1 vccd1 vccd1 _07845_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__12089__B2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09510_ _09507_/X _09509_/X _07091_/Y vssd1 vssd1 vccd1 vccd1 _09528_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09441_ reg1_val[2] reg1_val[29] _09463_/S vssd1 vssd1 vccd1 vccd1 _09441_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09372_ _07200_/Y _10787_/B _10787_/C fanout44/X _09582_/A vssd1 vssd1 vccd1 vccd1
+ _09373_/B sky130_fd_sc_hd__o32a_1
XFILLER_0_87_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09257__A2 _10536_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08323_ _08401_/A _08401_/B vssd1 vssd1 vccd1 vccd1 _08402_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_117_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09662__C1 _11866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout237_A _12867_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08254_ _08205_/A _08205_/C _08205_/B vssd1 vssd1 vccd1 vccd1 _08257_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_62_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08425__A _09659_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07205_ _08821_/B2 fanout56/X _08821_/A1 fanout53/X vssd1 vssd1 vccd1 vccd1 _07206_/B
+ sky130_fd_sc_hd__o22a_1
X_08185_ _10263_/A _08185_/B vssd1 vssd1 vccd1 vccd1 _08286_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_104_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07136_ _09524_/A _13748_/A _13744_/A vssd1 vssd1 vccd1 vccd1 _09516_/B sky130_fd_sc_hd__or3_2
XFILLER_0_30_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07067_ _12452_/A _07077_/A _07079_/A vssd1 vssd1 vccd1 vccd1 _07067_/X sky130_fd_sc_hd__o21a_1
XANTENNA__12381__S _12515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07969_ _07969_/A _07969_/B vssd1 vssd1 vccd1 vccd1 _08030_/A sky130_fd_sc_hd__nand2_2
X_09708_ _07208_/B _12235_/C _12657_/B1 reg1_val[1] vssd1 vssd1 vccd1 vccd1 _09708_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09703__B _09703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10980_ _10628_/Y _11227_/A _10978_/Y vssd1 vssd1 vccd1 vccd1 _10980_/Y sky130_fd_sc_hd__a21oi_1
X_09639_ _09392_/Y _09406_/B _09404_/Y vssd1 vssd1 vccd1 vccd1 _09641_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_69_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11026__A _11027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12650_ _13668_/Q _12650_/B vssd1 vssd1 vccd1 vccd1 _12705_/B sky130_fd_sc_hd__or2_1
X_11601_ _12372_/A _12372_/B vssd1 vssd1 vccd1 vccd1 _11601_/X sky130_fd_sc_hd__or2_1
X_12581_ _12581_/A _12581_/B vssd1 vssd1 vccd1 vccd1 _12581_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_65_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11532_ _11533_/A _11533_/B vssd1 vssd1 vccd1 vccd1 _11532_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__10802__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11463_ _11463_/A _11463_/B vssd1 vssd1 vccd1 vccd1 _11463_/Y sky130_fd_sc_hd__nor2_1
X_13202_ _12614_/A _13598_/C hold29/X _13605_/A vssd1 vssd1 vccd1 vccd1 _13637_/D
+ sky130_fd_sc_hd__o211a_1
X_10414_ _10414_/A _10414_/B vssd1 vssd1 vccd1 vccd1 _10415_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_21_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11394_ _12093_/A _11394_/B vssd1 vssd1 vccd1 vccd1 _11401_/A sky130_fd_sc_hd__xnor2_1
X_13133_ _13133_/A _13133_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[30] sky130_fd_sc_hd__xnor2_4
XFILLER_0_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10345_ _10293_/A _10293_/B _10291_/X vssd1 vssd1 vccd1 vccd1 _10432_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09708__B1 _12657_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ reg1_val[16] _13129_/B vssd1 vssd1 vccd1 vccd1 _13065_/B sky130_fd_sc_hd__and2_1
X_10276_ _10277_/A _10277_/B vssd1 vssd1 vccd1 vccd1 _10278_/A sky130_fd_sc_hd__and2_1
X_12015_ _11907_/A _11906_/B _11906_/A vssd1 vssd1 vccd1 vccd1 _12021_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__07195__B1 _07521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12917_ _12922_/B _12917_/B vssd1 vssd1 vccd1 vccd1 new_PC[17] sky130_fd_sc_hd__xnor2_4
XANTENNA__11294__A2 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12848_ _13015_/B _12848_/B vssd1 vssd1 vccd1 vccd1 _12849_/B sky130_fd_sc_hd__or2_1
XFILLER_0_61_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12779_ _12742_/B _12743_/A _12742_/A vssd1 vssd1 vccd1 vccd1 _12780_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_56_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12243__B2 _10866_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13440__B1 _13444_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13151__A _13151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08245__A _11708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09947__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09990_ _10579_/A _10579_/B _09988_/X _09989_/X vssd1 vssd1 vccd1 vccd1 _09991_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_122_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07295__S _07572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07973__A2 _11732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08941_ _08271_/A _09910_/A1 _07420_/Y _09501_/A vssd1 vssd1 vccd1 vccd1 _08942_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11506__B1 _07891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08872_ _08901_/A _08901_/B _08872_/C vssd1 vssd1 vccd1 vccd1 _08877_/A sky130_fd_sc_hd__nand3_2
XANTENNA__13685__CLK _13701_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07725__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07823_ _08923_/B1 fanout21/X _08246_/B _07347_/X vssd1 vssd1 vccd1 vccd1 _07824_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10190__C1 _10189_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout187_A _07118_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07754_ _07757_/A _07757_/B vssd1 vssd1 vccd1 vccd1 _07772_/B sky130_fd_sc_hd__nand2_1
X_07685_ _07686_/B _07686_/A vssd1 vssd1 vccd1 vccd1 _07780_/B sky130_fd_sc_hd__and2b_1
X_09424_ _09424_/A _09424_/B vssd1 vssd1 vccd1 vccd1 _09426_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_87_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09355_ _09575_/A _09355_/B vssd1 vssd1 vccd1 vccd1 _09357_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06882__B _07281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08306_ _08806_/A2 wire122/A _13166_/A1 _08806_/B1 vssd1 vssd1 vccd1 vccd1 _08307_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10245__B1 fanout79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09286_ _09286_/A _09286_/B vssd1 vssd1 vccd1 vccd1 _09287_/B sky130_fd_sc_hd__or2_1
XFILLER_0_47_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08237_ _08236_/A _08236_/B _08236_/C vssd1 vssd1 vccd1 vccd1 _08993_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_7_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09685__S _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12537__A2 _12793_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08168_ _08168_/A _08168_/B vssd1 vssd1 vccd1 vccd1 _08232_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07119_ instruction[2] instruction[1] pred_val instruction[0] vssd1 vssd1 vccd1 vccd1
+ _07122_/B sky130_fd_sc_hd__and4b_1
X_08099_ _08109_/B _08109_/A vssd1 vssd1 vccd1 vccd1 _08099_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_30_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10130_ _10130_/A _10130_/B vssd1 vssd1 vccd1 vccd1 _10131_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_101_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10061_ _10282_/A _10061_/B vssd1 vssd1 vccd1 vccd1 _10063_/B sky130_fd_sc_hd__nor2_2
XANTENNA__09433__B _13748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07234__A _09950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10963_ _10796_/A _10796_/B _10830_/A vssd1 vssd1 vccd1 vccd1 _10966_/A sky130_fd_sc_hd__o21bai_1
XANTENNA__11276__A2 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12473__B2 _12710_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10298__C _10577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12702_ hold247/A _12702_/B vssd1 vssd1 vccd1 vccd1 _12746_/B sky130_fd_sc_hd__or2_1
X_13682_ _13693_/CLK _13682_/D vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dfxtp_1
X_10894_ _10458_/S _10457_/X _09537_/B vssd1 vssd1 vccd1 vccd1 _12225_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_128_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12633_ _12733_/B vssd1 vssd1 vccd1 vccd1 _12633_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08429__B1 _10637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13422__B1 _13444_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06792__B _07398_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12776__A2 _09254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12564_ _12565_/A _12565_/B _12565_/C vssd1 vssd1 vccd1 vccd1 _12625_/B sky130_fd_sc_hd__o21a_1
X_11515_ _11516_/A _11516_/B vssd1 vssd1 vccd1 vccd1 _11610_/A sky130_fd_sc_hd__nand2_1
X_12495_ _12614_/A fanout8/X fanout3/X _07257_/X vssd1 vssd1 vccd1 vccd1 _12557_/D
+ sky130_fd_sc_hd__a22o_1
X_11446_ _11447_/B _11447_/A vssd1 vssd1 vccd1 vccd1 _11551_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_1_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11377_ _10458_/S _09852_/X _09537_/B vssd1 vssd1 vccd1 vccd1 _11377_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13116_ reg1_val[27] _13136_/A vssd1 vssd1 vccd1 vccd1 _13121_/B sky130_fd_sc_hd__xnor2_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10328_ _07160_/Y _12235_/C _12657_/B1 reg1_val[5] vssd1 vssd1 vccd1 vccd1 _10328_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ reg1_val[13] _13048_/B vssd1 vssd1 vccd1 vccd1 _13049_/A sky130_fd_sc_hd__or2_1
XANTENNA__07128__B _07129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10259_ _10259_/A _10259_/B vssd1 vssd1 vccd1 vccd1 _10277_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_56_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12161__B1 _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08904__A1 _07238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08904__B2 _07239_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06967__B _06980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08668__B1 _09173_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07470_ _07456_/A _07186_/B _07186_/C _07183_/Y _07476_/B vssd1 vssd1 vccd1 vccd1
+ _07472_/B sky130_fd_sc_hd__a41o_4
XFILLER_0_88_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09140_ _07237_/Y fanout44/X _07597_/X _08950_/B vssd1 vssd1 vccd1 vccd1 _09141_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09071_ _09077_/B _09071_/B _09079_/A vssd1 vssd1 vccd1 vccd1 _09073_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_16_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08022_ _08022_/A _08022_/B vssd1 vssd1 vccd1 vccd1 _08024_/B sky130_fd_sc_hd__and2_1
XFILLER_0_4_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08703__A _08746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09396__A1 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout5 fanout5/A vssd1 vssd1 vccd1 vccd1 fanout5/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__09396__B2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13192__A2 _13194_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07319__A _13015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09973_ _09974_/A _09974_/B vssd1 vssd1 vccd1 vccd1 _09973_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_110_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08924_ _09659_/B _08924_/B vssd1 vssd1 vccd1 vccd1 _08931_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12152__B1 _11688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08855_ _09950_/A _08855_/B vssd1 vssd1 vccd1 vccd1 _08887_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06906__B1 _06906_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07806_ _08008_/A vssd1 vssd1 vccd1 vccd1 _07808_/A sky130_fd_sc_hd__inv_2
XANTENNA__12598__C _12598_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08786_ _08786_/A _08786_/B vssd1 vssd1 vccd1 vccd1 _09044_/B sky130_fd_sc_hd__xor2_2
XANTENNA__06921__A3 _13059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07737_ fanout56/X _08821_/A1 fanout40/X _08821_/B2 vssd1 vssd1 vccd1 vccd1 _07738_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13490__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10466__B1 _12657_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07668_ _07668_/A _07668_/B vssd1 vssd1 vccd1 vccd1 _07749_/B sky130_fd_sc_hd__or2_1
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09407_ _09408_/A _09408_/B vssd1 vssd1 vccd1 vccd1 _09409_/A sky130_fd_sc_hd__and2_1
XFILLER_0_109_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07599_ _09950_/A _07599_/B vssd1 vssd1 vccd1 vccd1 _07601_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09338_ _09338_/A _09338_/B vssd1 vssd1 vccd1 vccd1 _09340_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_75_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12758__A2 _12793_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10769__A1 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10769__B2 fanout50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout15_A _07417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08831__B1 _13149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09269_ _09604_/A fanout9/X fanout4/X _09161_/A vssd1 vssd1 vccd1 vccd1 _09270_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11300_ _11300_/A _11300_/B vssd1 vssd1 vccd1 vccd1 _11301_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13168__C1 _13543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12280_ _12280_/A _12280_/B vssd1 vssd1 vccd1 vccd1 _12281_/B sky130_fd_sc_hd__or2_1
XFILLER_0_16_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11718__B1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11231_ _11231_/A _12372_/A _11600_/A vssd1 vssd1 vccd1 vccd1 _11231_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__09428__B _13744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07229__A _07230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11162_ _11162_/A _11162_/B vssd1 vssd1 vccd1 vccd1 _11163_/B sky130_fd_sc_hd__nor2_1
X_10113_ _10113_/A _10113_/B vssd1 vssd1 vccd1 vccd1 _10130_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_101_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11093_ _10967_/A _10967_/B _10965_/X vssd1 vssd1 vccd1 vccd1 _11095_/B sky130_fd_sc_hd__a21bo_1
X_10044_ _10044_/A _10726_/C vssd1 vssd1 vccd1 vccd1 _10200_/A sky130_fd_sc_hd__nor2_1
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11995_ _12107_/A _11995_/B vssd1 vssd1 vccd1 vccd1 _12000_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_58_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13734_ _13735_/CLK _13734_/D vssd1 vssd1 vccd1 vccd1 hold299/A sky130_fd_sc_hd__dfxtp_1
X_10946_ _11072_/A _10946_/B vssd1 vssd1 vccd1 vccd1 _10950_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13665_ _13719_/CLK _13665_/D vssd1 vssd1 vccd1 vccd1 hold216/A sky130_fd_sc_hd__dfxtp_1
X_10877_ _09676_/X _09684_/X _11472_/S vssd1 vssd1 vccd1 vccd1 _10877_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_85_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10209__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12616_ _12675_/B _12616_/B vssd1 vssd1 vccd1 vccd1 _12620_/A sky130_fd_sc_hd__or2_1
XFILLER_0_38_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13596_ hold3/X _13592_/X _13595_/Y rst vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__a211oi_1
XFILLER_0_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07625__A1 fanout39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12547_ curr_PC[27] _12546_/B _12971_/S vssd1 vssd1 vccd1 vccd1 _12547_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07625__B2 _07557_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11421__A2 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09619__A _12094_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12478_ curr_PC[25] _12405_/X _07108_/D vssd1 vssd1 vccd1 vccd1 _12478_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__08523__A _11286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_3 _10170_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13174__A2 _13194_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11429_ _11430_/A _11430_/B vssd1 vssd1 vccd1 vccd1 _11431_/A sky130_fd_sc_hd__or2_1
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07139__A _13744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06970_ reg1_val[8] _07449_/A vssd1 vssd1 vccd1 vccd1 _10867_/B sky130_fd_sc_hd__and2_1
XFILLER_0_67_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06978__A _13015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09550__A1 _10225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08640_ _10944_/A _08640_/B vssd1 vssd1 vccd1 vccd1 _08662_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09550__B2 _10104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07561__B1 _09885_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08571_ _08571_/A _08571_/B vssd1 vssd1 vccd1 vccd1 _09057_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_89_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07522_ _07522_/A _07523_/B vssd1 vssd1 vccd1 vccd1 _07522_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__07313__B1 wire101/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07453_ _11800_/A _07453_/B vssd1 vssd1 vccd1 vccd1 _07453_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_64_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11124__A _11126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07384_ reg1_val[24] _07634_/B _07634_/C vssd1 vssd1 vccd1 vccd1 _07384_/X sky130_fd_sc_hd__or3_1
X_09123_ _10078_/A _09123_/B vssd1 vssd1 vccd1 vccd1 _09130_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09054_ _09055_/B _09055_/C _09055_/A vssd1 vssd1 vccd1 vccd1 _11864_/C sky130_fd_sc_hd__a21o_1
XANTENNA__09529__A _13135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08005_ _10944_/A _08005_/B vssd1 vssd1 vccd1 vccd1 _08044_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09956_ _09783_/A _09783_/B _09779_/X vssd1 vssd1 vccd1 vccd1 _09960_/A sky130_fd_sc_hd__a21oi_2
X_08907_ _08907_/A _08907_/B _08907_/C vssd1 vssd1 vccd1 vccd1 _08908_/C sky130_fd_sc_hd__or3_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _09887_/A vssd1 vssd1 vccd1 vccd1 _09894_/A sky130_fd_sc_hd__inv_2
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09541__A1 _13145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08838_ _08838_/A _08838_/B vssd1 vssd1 vccd1 vccd1 _08860_/B sky130_fd_sc_hd__xnor2_1
X_08769_ _08821_/B2 _09216_/B2 _08868_/B1 _08821_/A1 vssd1 vssd1 vccd1 vccd1 _08770_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10439__B1 _10981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10800_ _12668_/A _10800_/B vssd1 vssd1 vccd1 vccd1 _10801_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11780_ _11484_/X _11779_/X _12525_/A vssd1 vssd1 vccd1 vccd1 _11780_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10857__B _10981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10731_ _11562_/A _10731_/B _10731_/C vssd1 vssd1 vccd1 vccd1 _10731_/X sky130_fd_sc_hd__or3_1
XFILLER_0_67_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07855__A1 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07855__B2 _08395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11552__A_N _11550_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11034__A _12253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13450_ hold262/X _13450_/B vssd1 vssd1 vccd1 vccd1 _13450_/X sky130_fd_sc_hd__and2_1
X_10662_ _11719_/A _10662_/B vssd1 vssd1 vccd1 vccd1 _10664_/B sky130_fd_sc_hd__xnor2_1
X_12401_ _12394_/Y _12395_/X _12400_/X vssd1 vssd1 vccd1 vccd1 _12401_/X sky130_fd_sc_hd__o21ba_1
X_13381_ _13605_/A hold155/X vssd1 vssd1 vccd1 vccd1 hold156/A sky130_fd_sc_hd__and2_1
X_10593_ _10592_/A _10592_/B _10592_/Y _12047_/C1 vssd1 vssd1 vccd1 vccd1 _10593_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12332_ _12411_/A _12332_/B vssd1 vssd1 vccd1 vccd1 _12334_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__11688__B _11688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13156__A2 _13196_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12263_ _12182_/A _12182_/B _12174_/A vssd1 vssd1 vccd1 vccd1 _12278_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_105_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11214_ _11215_/B _11215_/A vssd1 vssd1 vccd1 vccd1 _11214_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_121_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12194_ _12195_/A _12195_/B vssd1 vssd1 vccd1 vccd1 _12283_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08583__A2 _10049_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11145_ _12760_/A1 _11132_/X _11144_/X _11123_/X vssd1 vssd1 vccd1 vccd1 _11145_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__07791__B1 fanout66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09174__A _10266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11076_ _11076_/A _11076_/B vssd1 vssd1 vccd1 vccd1 _11078_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08335__A2 fanout24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10027_ hold243/A _13642_/Q hold188/A vssd1 vssd1 vccd1 vccd1 _10027_/X sky130_fd_sc_hd__or3_1
XFILLER_0_98_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11978_ _07337_/Y _07431_/Y _12754_/C _11975_/Y vssd1 vssd1 vccd1 vccd1 _11978_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10929_ _10929_/A _10929_/B vssd1 vssd1 vccd1 vccd1 _10931_/B sky130_fd_sc_hd__xnor2_1
X_13717_ _13717_/CLK _13717_/D vssd1 vssd1 vccd1 vccd1 hold271/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13143__B _13207_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13648_ _13649_/CLK _13648_/D vssd1 vssd1 vccd1 vccd1 hold180/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12982__B _12982_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13395__A2 _13207_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13579_ _13579_/A _13579_/B _13579_/C vssd1 vssd1 vccd1 vccd1 _13580_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06980__B _06980_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11158__B2 _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09810_ _09642_/A _09642_/B _09640_/Y vssd1 vssd1 vccd1 vccd1 _09817_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09771__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09771__B2 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09741_ _09592_/Y _09599_/B _09597_/Y vssd1 vssd1 vccd1 vccd1 _09747_/A sky130_fd_sc_hd__o21ai_2
X_06953_ _06928_/A _06936_/B _13036_/B _06952_/X vssd1 vssd1 vccd1 vccd1 _07455_/A
+ sky130_fd_sc_hd__a31o_2
XANTENNA__08326__A2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09672_ _09670_/X _09671_/X _10005_/S vssd1 vssd1 vccd1 vccd1 _09672_/X sky130_fd_sc_hd__mux2_1
X_06884_ _06884_/A _06884_/B vssd1 vssd1 vccd1 vccd1 _11961_/A sky130_fd_sc_hd__nor2_2
XANTENNA__07534__B1 _07535_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08623_ _08653_/A _08653_/B vssd1 vssd1 vccd1 vccd1 _08982_/A sky130_fd_sc_hd__or2_1
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout267_A _06920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08554_ _08555_/B _08555_/A vssd1 vssd1 vccd1 vccd1 _08559_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_77_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09826__A2 _09426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07505_ _07505_/A _07505_/B vssd1 vssd1 vccd1 vccd1 _07506_/B sky130_fd_sc_hd__nor2_2
XANTENNA__13053__B _13054_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08485_ _08485_/A _08485_/B vssd1 vssd1 vccd1 vccd1 _08553_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07436_ reg1_val[16] _07634_/B reg1_val[17] vssd1 vssd1 vccd1 vccd1 _07436_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_64_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07367_ _07367_/A _07367_/B vssd1 vssd1 vccd1 vccd1 _10225_/A sky130_fd_sc_hd__nand2_8
XANTENNA__11397__A1 fanout44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09106_ _07347_/X _07699_/B _13151_/A fanout35/X vssd1 vssd1 vccd1 vccd1 _09107_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12594__B1 _12795_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11397__B2 _07597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07298_ _07297_/A _07192_/A _07192_/B _07521_/A vssd1 vssd1 vccd1 vccd1 _07300_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_103_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09037_ _09044_/C _09044_/D _09044_/B vssd1 vssd1 vccd1 vccd1 _09039_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12413__A _12413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout82_A _07522_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10372__A2 _07643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09939_ _10814_/A1 fanout25/X fanout23/X fanout42/X vssd1 vssd1 vccd1 vccd1 _09940_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12649__A1 _12648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08317__A2 _10538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12950_ _12935_/B _12943_/B _12956_/A vssd1 vssd1 vccd1 vccd1 _12963_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__07525__B1 _07476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11901_ _12668_/A _11901_/B vssd1 vssd1 vccd1 vccd1 _11905_/A sky130_fd_sc_hd__xnor2_1
X_12881_ reg1_val[12] curr_PC[12] _12978_/S vssd1 vssd1 vccd1 vccd1 _12883_/B sky130_fd_sc_hd__mux2_1
X_11832_ _11832_/A _11832_/B vssd1 vssd1 vccd1 vccd1 _11833_/B sky130_fd_sc_hd__nand2_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11763_ _11763_/A _11950_/A vssd1 vssd1 vccd1 vccd1 _11763_/Y sky130_fd_sc_hd__nand2_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _10715_/A _10715_/B vssd1 vssd1 vccd1 vccd1 _10714_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_82_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13502_ _13543_/A _13502_/B vssd1 vssd1 vccd1 vccd1 _13716_/D sky130_fd_sc_hd__and2_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _09860_/A _11592_/Y _11692_/Y _11693_/X vssd1 vssd1 vccd1 vccd1 _11694_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_83_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13433_ _12421_/A _13598_/C hold96/X vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__o21a_1
X_10645_ _10508_/A _10508_/B _10511_/A vssd1 vssd1 vccd1 vccd1 _10656_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_125_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13364_ _13663_/Q _13542_/B2 _13555_/A2 hold205/X vssd1 vssd1 vccd1 vccd1 hold206/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08073__A _11708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10576_ _10857_/A _10981_/A vssd1 vssd1 vccd1 vccd1 _10576_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_51_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12315_ hold282/A _12314_/X _09521_/Y vssd1 vssd1 vccd1 vccd1 _12315_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13295_ _13503_/B _13504_/A _13257_/X vssd1 vssd1 vccd1 vccd1 _13509_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12337__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12246_ _12406_/B1 _12243_/X _12245_/X vssd1 vssd1 vccd1 vccd1 dest_val[22] sky130_fd_sc_hd__o21ai_4
XFILLER_0_121_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08801__A _09371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10348__C1 _10518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12177_ _12177_/A fanout5/X vssd1 vssd1 vccd1 vccd1 _12177_/X sky130_fd_sc_hd__or2_1
XANTENNA__07764__B1 _13151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11128_ _10995_/X _10999_/X _11124_/X _11126_/Y vssd1 vssd1 vccd1 vccd1 _11129_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07136__B _13748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11059_ _11059_/A _11059_/B vssd1 vssd1 vccd1 vccd1 _11061_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11863__A2 _12163_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09269__B1 fanout4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08270_ _07283_/A _07283_/B _08328_/B2 vssd1 vssd1 vccd1 vccd1 _08272_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08492__A1 _08923_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08492__B2 _08866_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07221_ _07221_/A _07521_/A vssd1 vssd1 vccd1 vccd1 _07221_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11379__A1 _12537_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11379__B2 _12760_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12576__B1 _09429_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08244__A1 _08923_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07152_ _13748_/A _13744_/A instruction[5] _10889_/B vssd1 vssd1 vccd1 vccd1 _07152_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08244__B2 _08866_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07083_ _12642_/A _07082_/Y _07062_/Y vssd1 vssd1 vccd1 vccd1 _07083_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_112_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout104 _07276_/X vssd1 vssd1 vccd1 vccd1 _08873_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout115 _07471_/Y vssd1 vssd1 vccd1 vccd1 _11047_/A sky130_fd_sc_hd__buf_8
XANTENNA__07755__B1 _07557_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout126 _07311_/Y vssd1 vssd1 vccd1 vccd1 _08806_/B1 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10354__A2 _10787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout137 _12695_/A vssd1 vssd1 vccd1 vccd1 _12130_/A sky130_fd_sc_hd__buf_4
XANTENNA__07327__A _11126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13048__B _13048_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07985_ _07989_/A _07989_/B vssd1 vssd1 vccd1 vccd1 _07985_/X sky130_fd_sc_hd__and2_1
Xfanout159 _13196_/A2 vssd1 vssd1 vccd1 vccd1 _13194_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09724_ _09649_/A _09649_/B _09647_/X vssd1 vssd1 vccd1 vccd1 _09824_/A sky130_fd_sc_hd__a21oi_4
X_06936_ _06936_/A _06936_/B _13048_/B vssd1 vssd1 vccd1 vccd1 _06936_/X sky130_fd_sc_hd__and3_1
XANTENNA__10106__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09655_ _10298_/A _09655_/B vssd1 vssd1 vccd1 vccd1 _09656_/C sky130_fd_sc_hd__xor2_2
X_06867_ _07483_/A _07201_/A vssd1 vssd1 vccd1 vccd1 _06869_/A sky130_fd_sc_hd__and2_1
XFILLER_0_96_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08180__B1 _08486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06885__B _12981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08606_ _08606_/A _08606_/B vssd1 vssd1 vccd1 vccd1 _08609_/A sky130_fd_sc_hd__xnor2_1
X_09586_ _09779_/A _09586_/B _09586_/C vssd1 vssd1 vccd1 vccd1 _09753_/A sky130_fd_sc_hd__nand3_2
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06798_ _06796_/Y _06872_/B1 _06873_/B1 reg2_val[27] vssd1 vssd1 vccd1 vccd1 _07252_/A
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08537_ _08866_/A2 _10538_/A _08778_/B _09216_/B2 vssd1 vssd1 vccd1 vccd1 _08538_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10814__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08468_ _08413_/X _08467_/Y _08412_/X vssd1 vssd1 vccd1 vccd1 _08988_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07286__A2 _07213_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07419_ _07419_/A _07420_/B vssd1 vssd1 vccd1 vccd1 _13151_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_18_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08399_ _08408_/B _08408_/A vssd1 vssd1 vccd1 vccd1 _08399_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_80_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10430_ _10432_/A _10432_/B vssd1 vssd1 vccd1 vccd1 _10430_/X sky130_fd_sc_hd__or2_1
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10361_ _10264_/Y _10271_/B _10269_/Y vssd1 vssd1 vccd1 vccd1 _10363_/B sky130_fd_sc_hd__o21a_2
XANTENNA_clkbuf_4_1_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12100_ _12100_/A _12100_/B vssd1 vssd1 vccd1 vccd1 _12114_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11790__A1 _12760_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13080_ reg1_val[20] _13129_/B vssd1 vssd1 vccd1 vccd1 _13102_/A sky130_fd_sc_hd__xnor2_2
X_10292_ _10292_/A _10292_/B vssd1 vssd1 vccd1 vccd1 _10293_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_103_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12031_ _12032_/A _12032_/B _12032_/C vssd1 vssd1 vccd1 vccd1 _12031_/X sky130_fd_sc_hd__o21a_1
Xhold180 hold180/A vssd1 vssd1 vccd1 vccd1 hold180/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12143__A _12782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold191 hold218/X vssd1 vssd1 vccd1 vccd1 hold191/X sky130_fd_sc_hd__buf_1
XANTENNA__07210__A2 _07572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12933_ reg1_val[20] curr_PC[20] _12978_/S vssd1 vssd1 vccd1 vccd1 _12935_/B sky130_fd_sc_hd__mux2_1
XANTENNA__06795__B _12981_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12864_ _12865_/A _12865_/B _12865_/C vssd1 vssd1 vccd1 vccd1 _12872_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_96_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11815_ _11816_/A _11816_/B vssd1 vssd1 vccd1 vccd1 _11929_/A sky130_fd_sc_hd__and2_1
X_12795_ _12795_/A1 _12785_/Y _12789_/Y _12794_/X vssd1 vssd1 vccd1 vccd1 _12795_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ _11746_/A _11746_/B vssd1 vssd1 vccd1 vccd1 _11749_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07700__A _10050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11677_ _07092_/D _11674_/X _11675_/X _12047_/C1 vssd1 vssd1 vccd1 vccd1 _11677_/X
+ sky130_fd_sc_hd__o31a_1
X_10628_ _10430_/X _10573_/X _10574_/X vssd1 vssd1 vccd1 vccd1 _10628_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__07029__A2 _06928_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13416_ hold22/X _13416_/A2 _13420_/B1 _13690_/Q _13383_/A vssd1 vssd1 vccd1 vccd1
+ hold23/A sky130_fd_sc_hd__o221a_1
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11230__B1 _11600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13347_ _13359_/A hold194/X vssd1 vssd1 vccd1 vccd1 _13655_/D sky130_fd_sc_hd__and2_1
X_10559_ _10422_/A _10422_/B _10420_/X vssd1 vssd1 vccd1 vccd1 _10567_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10584__A2 _10727_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13278_ hold285/A hold7/X vssd1 vssd1 vccd1 vccd1 _13460_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_59_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08529__A2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13149__A _13149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12229_ _13663_/Q _12311_/B1 _12393_/C _12533_/B1 vssd1 vssd1 vccd1 vccd1 _12230_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__07737__B1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10336__A2 _12760_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07770_ _07770_/A _07770_/B _07770_/C vssd1 vssd1 vccd1 vccd1 _07813_/A sky130_fd_sc_hd__or3_1
XFILLER_0_75_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12089__A2 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09440_ reg1_val[3] reg1_val[28] _09463_/S vssd1 vssd1 vccd1 vccd1 _09440_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09371_ _09371_/A _09371_/B vssd1 vssd1 vccd1 vccd1 _09377_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08322_ _08322_/A _08322_/B vssd1 vssd1 vccd1 vccd1 _08401_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07610__A _10078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10272__A1 _10104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08253_ _08347_/A _08347_/B _08252_/A vssd1 vssd1 vccd1 vccd1 _08282_/A sky130_fd_sc_hd__a21o_1
XANTENNA_fanout132_A _07237_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07204_ _07212_/B _07204_/B vssd1 vssd1 vccd1 vccd1 _07204_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10328__A2_N _12235_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08184_ _13149_/A fanout28/X _08395_/B _08923_/B1 vssd1 vssd1 vccd1 vccd1 _08185_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07135_ instruction[30] instruction[23] _07135_/S vssd1 vssd1 vccd1 vccd1 reg2_idx[5]
+ sky130_fd_sc_hd__mux2_8
XFILLER_0_15_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07976__B1 _07544_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07066_ reg1_val[24] _07221_/A vssd1 vssd1 vccd1 vccd1 _07077_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08441__A _08746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07440__A2 _07435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09717__B2 _09839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07728__B1 _08704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10327__A2 _12314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ _07968_/A _08028_/A _07968_/C vssd1 vssd1 vccd1 vccd1 _07969_/B sky130_fd_sc_hd__nand3_1
XANTENNA__06896__A _06936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06919_ _11586_/A _06919_/B vssd1 vssd1 vccd1 vccd1 _07094_/A sky130_fd_sc_hd__nand2_1
X_09707_ hold262/A hold245/A _12314_/A _12796_/A1 vssd1 vssd1 vccd1 vccd1 _09707_/X
+ sky130_fd_sc_hd__a31o_1
X_07899_ _07899_/A _07899_/B vssd1 vssd1 vccd1 vccd1 _07900_/B sky130_fd_sc_hd__or2_1
X_09638_ _09390_/A _09390_/B _09388_/Y vssd1 vssd1 vccd1 vccd1 _09641_/A sky130_fd_sc_hd__o21a_1
X_09569_ fanout45/X _07307_/Y _08833_/B fanout49/X vssd1 vssd1 vccd1 vccd1 _09570_/B
+ sky130_fd_sc_hd__o22a_1
X_11600_ _11600_/A _11600_/B _11458_/B _11561_/B vssd1 vssd1 vccd1 vccd1 _12372_/B
+ sky130_fd_sc_hd__or4bb_1
XANTENNA__12788__B1 _12598_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12580_ _12738_/S _12579_/Y _12578_/X vssd1 vssd1 vccd1 vccd1 _12581_/B sky130_fd_sc_hd__a21o_1
X_11531_ _11531_/A _11531_/B vssd1 vssd1 vccd1 vccd1 _11533_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11462_ _07094_/C _11354_/B _06934_/B vssd1 vssd1 vccd1 vccd1 _11463_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13201_ hold28/X _13207_/B vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__or2_1
XFILLER_0_123_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10413_ _10414_/B _10414_/A vssd1 vssd1 vccd1 vccd1 _10413_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11393_ fanout50/X fanout20/X fanout18/X _12557_/A vssd1 vssd1 vccd1 vccd1 _11394_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13132_ _13126_/B _13128_/B _13126_/A vssd1 vssd1 vccd1 vccd1 _13133_/B sky130_fd_sc_hd__a21bo_2
X_10344_ _10344_/A _10727_/A vssd1 vssd1 vccd1 vccd1 _10344_/X sky130_fd_sc_hd__or2_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13063_ reg1_val[16] _13129_/B vssd1 vssd1 vccd1 vccd1 _13065_/A sky130_fd_sc_hd__nor2_1
X_10275_ _10275_/A _10275_/B vssd1 vssd1 vccd1 vccd1 _10277_/B sky130_fd_sc_hd__xnor2_1
X_12014_ _12014_/A _12014_/B vssd1 vssd1 vccd1 vccd1 _12024_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07195__A1 _07201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08144__B1 _07545_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12916_ _12956_/A _12910_/B _12922_/A vssd1 vssd1 vccd1 vccd1 _12917_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_69_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12847_ _13015_/B _12848_/B vssd1 vssd1 vccd1 vccd1 _12858_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_84_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _12778_/A _12778_/B vssd1 vssd1 vccd1 vccd1 _12778_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_84_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13151__B _13193_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11729_ _11802_/B _11729_/B vssd1 vssd1 vccd1 vccd1 _11735_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12990__B _12990_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09947__A1 _07175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09947__B2 _08933_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08940_ _09371_/A _08940_/B vssd1 vssd1 vccd1 vccd1 _08959_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11506__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11506__B2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08871_ _09948_/A _08871_/B vssd1 vssd1 vccd1 vccd1 _08872_/C sky130_fd_sc_hd__xnor2_1
X_07822_ _09940_/A _07822_/B vssd1 vssd1 vccd1 vccd1 _07828_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07180__B_N _07556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07605__A _10095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07753_ _09940_/A _07753_/B vssd1 vssd1 vccd1 vccd1 _07757_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07684_ _07780_/A _07684_/B vssd1 vssd1 vccd1 vccd1 _07686_/B sky130_fd_sc_hd__or2_1
XANTENNA__07489__A2 _07363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09423_ _09423_/A _09423_/B vssd1 vssd1 vccd1 vccd1 _09424_/B sky130_fd_sc_hd__xor2_4
XANTENNA__11690__B1 _12754_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09354_ fanout56/X fanout68/X fanout66/X fanout53/X vssd1 vssd1 vccd1 vccd1 _09355_/B
+ sky130_fd_sc_hd__o22a_1
X_08305_ _10236_/A _08305_/B vssd1 vssd1 vccd1 vccd1 _08377_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_35_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10245__A1 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10245__B2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09285_ _09286_/A _09286_/B vssd1 vssd1 vccd1 vccd1 _09346_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_34_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08236_ _08236_/A _08236_/B _08236_/C vssd1 vssd1 vccd1 vccd1 _08236_/X sky130_fd_sc_hd__and3_1
XFILLER_0_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08167_ _08167_/A _08235_/A _08167_/C vssd1 vssd1 vccd1 vccd1 _08167_/X sky130_fd_sc_hd__and3_1
XFILLER_0_30_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07118_ hold159/A _07118_/B vssd1 vssd1 vccd1 vccd1 busy sky130_fd_sc_hd__nor2_8
XFILLER_0_101_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08098_ _08098_/A _08098_/B vssd1 vssd1 vccd1 vccd1 _08109_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07049_ _11958_/B _11958_/C _11961_/A vssd1 vssd1 vccd1 vccd1 _07050_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__10206__A _12092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10060_ _10060_/A _10060_/B _10060_/C vssd1 vssd1 vccd1 vccd1 _10061_/B sky130_fd_sc_hd__and3_1
XANTENNA__08374__B1 _11638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13517__A _13543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12421__A _12421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10962_ _10962_/A _10962_/B vssd1 vssd1 vccd1 vccd1 _10967_/A sky130_fd_sc_hd__or2_1
XFILLER_0_15_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09730__A _11731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10298__D _10631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12701_ _12648_/A _09839_/B _12700_/X _09529_/B vssd1 vssd1 vccd1 vccd1 _12701_/X
+ sky130_fd_sc_hd__a211o_1
X_10893_ _10891_/X _10893_/B _10893_/C _10893_/D vssd1 vssd1 vccd1 vccd1 _10893_/X
+ sky130_fd_sc_hd__and4b_1
X_13681_ _13693_/CLK _13681_/D vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08429__A1 _08806_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12632_ _12728_/A _12632_/B vssd1 vssd1 vccd1 vccd1 _12733_/B sky130_fd_sc_hd__xor2_2
XANTENNA__08429__B2 _08806_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07250__A _10239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12563_ _12625_/A _12563_/B vssd1 vssd1 vccd1 vccd1 _12565_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11984__A1 _07281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11514_ _11514_/A _11514_/B vssd1 vssd1 vccd1 vccd1 _11516_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_25_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12494_ _12494_/A _12494_/B vssd1 vssd1 vccd1 vccd1 _12499_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11445_ _11445_/A _11445_/B vssd1 vssd1 vccd1 vccd1 _11447_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11376_ _11370_/Y _11371_/X _11372_/X _11375_/X vssd1 vssd1 vccd1 vccd1 _11376_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13115_ _13111_/A _13114_/B _13111_/B vssd1 vssd1 vccd1 vccd1 _13117_/A sky130_fd_sc_hd__a21bo_1
X_10327_ hold294/A _12314_/A _10325_/X _12796_/A1 vssd1 vssd1 vccd1 vccd1 _10327_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _13051_/B _13046_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[12] sky130_fd_sc_hd__and2_4
XANTENNA__09905__A _10119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10258_ _10256_/Y _10258_/B vssd1 vssd1 vccd1 vccd1 _10259_/B sky130_fd_sc_hd__and2b_1
XANTENNA__08904__A2 _09910_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10189_ _07168_/X _12235_/C _12657_/B1 reg1_val[4] vssd1 vssd1 vccd1 vccd1 _10189_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12331__A _12331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08668__A1 _08866_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08668__B2 _08950_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10786__A _11076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13413__A1 _11281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09070_ _08467_/Y _08567_/X _08469_/Y vssd1 vssd1 vccd1 vccd1 _09079_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_44_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08021_ _08021_/A _08021_/B _08021_/C vssd1 vssd1 vccd1 vccd1 _08022_/B sky130_fd_sc_hd__or3_1
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09396__A2 _07522_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout6 fanout7/A vssd1 vssd1 vccd1 vccd1 fanout6/X sky130_fd_sc_hd__buf_4
XFILLER_0_110_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09972_ _09802_/A _09802_/B _09803_/X vssd1 vssd1 vccd1 vccd1 _09974_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_110_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08923_ _08197_/A _08907_/B _08907_/C _08923_/B1 _08907_/A vssd1 vssd1 vccd1 vccd1
+ _08924_/B sky130_fd_sc_hd__o32ai_2
XFILLER_0_110_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08854_ _08197_/A _10522_/A _08868_/B1 _08907_/A vssd1 vssd1 vccd1 vccd1 _08855_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_99_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07805_ _10095_/A _07805_/B vssd1 vssd1 vccd1 vccd1 _08008_/A sky130_fd_sc_hd__xnor2_2
X_08785_ _08786_/A _08786_/B _08788_/A _08788_/B vssd1 vssd1 vccd1 vccd1 _08785_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_07736_ _10078_/A _07736_/B vssd1 vssd1 vccd1 vccd1 _07741_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_79_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07054__B _07201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07667_ _07667_/A _07667_/B vssd1 vssd1 vccd1 vccd1 _07668_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_48_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09406_ _09406_/A _09406_/B vssd1 vssd1 vccd1 vccd1 _09408_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07598_ _08907_/A fanout44/X _07597_/X _08328_/B2 vssd1 vssd1 vccd1 vccd1 _07599_/B
+ sky130_fd_sc_hd__o22a_1
X_09337_ _09337_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09338_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_35_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10769__A2 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09268_ _12717_/A _12764_/B _12718_/B vssd1 vssd1 vccd1 vccd1 fanout4/A sky130_fd_sc_hd__o21ai_2
XANTENNA__08831__A1 _08873_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08831__B2 _08891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08219_ _08256_/A _08217_/B _08291_/A vssd1 vssd1 vccd1 vccd1 _08243_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09199_ _09200_/B _09200_/A vssd1 vssd1 vccd1 vccd1 _09199_/X sky130_fd_sc_hd__and2b_1
XANTENNA__11718__A1 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10862__C _10900_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11230_ _11864_/A _12372_/A _11600_/A vssd1 vssd1 vccd1 vccd1 _11230_/X sky130_fd_sc_hd__a21o_1
XANTENNA__11718__B2 _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12391__A1 _12314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08595__B1 _09885_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11161_ _11161_/A _11161_/B _11161_/C vssd1 vssd1 vccd1 vccd1 _11162_/B sky130_fd_sc_hd__and3_1
XFILLER_0_101_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10112_ _10112_/A _10112_/B vssd1 vssd1 vccd1 vccd1 _10113_/B sky130_fd_sc_hd__xnor2_4
X_11092_ _11092_/A _11092_/B vssd1 vssd1 vccd1 vccd1 _11095_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13340__B1 _13506_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10043_ _10340_/C _10042_/X _12825_/S _10040_/Y vssd1 vssd1 vccd1 vccd1 dest_val[3]
+ sky130_fd_sc_hd__a2bb2o_4
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07570__A1 _13015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11990__A _12253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11994_ _11994_/A _11994_/B vssd1 vssd1 vccd1 vccd1 _11995_/B sky130_fd_sc_hd__and2_1
X_13733_ _13739_/CLK _13733_/D vssd1 vssd1 vccd1 vccd1 hold247/A sky130_fd_sc_hd__dfxtp_1
X_10945_ _10787_/A _07891_/X fanout10/X _07546_/X vssd1 vssd1 vccd1 vccd1 _10946_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13664_ _13719_/CLK _13664_/D vssd1 vssd1 vccd1 vccd1 hold229/A sky130_fd_sc_hd__dfxtp_1
X_10876_ _10876_/A _10876_/B vssd1 vssd1 vccd1 vccd1 _10880_/B sky130_fd_sc_hd__xor2_1
XANTENNA__10209__A1 fanout39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10209__B2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12615_ _12614_/A _12764_/B _12614_/C vssd1 vssd1 vccd1 vccd1 _12616_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13595_ hold191/X _13599_/D hold3/X vssd1 vssd1 vccd1 vccd1 _13595_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07625__A2 _07366_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12546_ curr_PC[27] _12546_/B vssd1 vssd1 vccd1 vccd1 _12546_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_41_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12477_ curr_PC[24] curr_PC[25] _12477_/C vssd1 vssd1 vccd1 vccd1 _12543_/B sky130_fd_sc_hd__and3_1
XANTENNA_4 _10464_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11428_ _11428_/A _11428_/B vssd1 vssd1 vccd1 vccd1 _11430_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11359_ reg1_val[13] curr_PC[13] vssd1 vssd1 vccd1 vccd1 _11360_/B sky130_fd_sc_hd__nand2_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08338__B1 _08395_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06978__B _07492_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ reg1_val[10] _13029_/B vssd1 vssd1 vccd1 vccd1 _13039_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09550__A2 _07643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07561__A1 _10049_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07561__B2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08570_ _08571_/A _08571_/B vssd1 vssd1 vccd1 vccd1 _08570_/X sky130_fd_sc_hd__and2_1
XFILLER_0_83_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10448__A1 _12515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07521_ _07521_/A _07521_/B vssd1 vssd1 vccd1 vccd1 _07523_/B sky130_fd_sc_hd__nor2_4
XFILLER_0_89_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07313__A1 _07300_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07313__B2 _10536_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07452_ _10889_/A _07452_/B vssd1 vssd1 vccd1 vccd1 wire122/A sky130_fd_sc_hd__xnor2_4
XANTENNA__11405__A _12417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10540__B1_N _09575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07383_ reg1_val[25] _07865_/B vssd1 vssd1 vccd1 vccd1 _07395_/A sky130_fd_sc_hd__or2_2
X_09122_ _07198_/Y _10536_/A1 _10536_/B2 _07203_/Y vssd1 vssd1 vccd1 vccd1 _09123_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09053_ _09046_/B _09046_/C _08983_/A _09046_/A _09052_/A vssd1 vssd1 vccd1 vccd1
+ _09055_/C sky130_fd_sc_hd__a2111o_1
XFILLER_0_32_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09529__B _09529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08004_ _09885_/B1 fanout84/X _08580_/B _10049_/A2 vssd1 vssd1 vccd1 vccd1 _08005_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_102_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_6_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09955_ _09955_/A _10518_/A vssd1 vssd1 vccd1 vccd1 _09961_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13322__B1 _13450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ _07367_/A _07367_/B _08197_/A vssd1 vssd1 vccd1 vccd1 _08908_/B sky130_fd_sc_hd__a21o_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ _10050_/A _09886_/B vssd1 vssd1 vccd1 vccd1 _09887_/A sky130_fd_sc_hd__xnor2_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09541__A2 _11793_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08837_ _08863_/A _08847_/B _08830_/Y vssd1 vssd1 vccd1 vccd1 _08860_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_99_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08768_ _08857_/A _08768_/B vssd1 vssd1 vccd1 vccd1 _08774_/A sky130_fd_sc_hd__xor2_1
X_07719_ _07719_/A _07719_/B vssd1 vssd1 vccd1 vccd1 _07842_/B sky130_fd_sc_hd__xnor2_2
X_08699_ _08699_/A _08699_/B vssd1 vssd1 vccd1 vccd1 _08700_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_79_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10857__C _10981_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10730_ _10729_/X _10730_/B _10730_/C vssd1 vssd1 vccd1 vccd1 _10730_/X sky130_fd_sc_hd__and3b_1
XANTENNA__07855__A2 _10915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10661_ fanout34/X fanout82/X _11423_/A fanout32/X vssd1 vssd1 vccd1 vccd1 _10662_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12400_ _09504_/Y _10596_/Y _10603_/X _12710_/B2 _12399_/X vssd1 vssd1 vccd1 vccd1
+ _12400_/X sky130_fd_sc_hd__a221o_1
XANTENNA__12061__B1 _11688_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13380_ hold224/A _13599_/D _13584_/B hold154/X vssd1 vssd1 vccd1 vccd1 hold155/A
+ sky130_fd_sc_hd__a22o_1
X_10592_ _10592_/A _10592_/B vssd1 vssd1 vccd1 vccd1 _10592_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_35_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12600__A2 _12799_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12331_ _12331_/A _12764_/B vssd1 vssd1 vccd1 vccd1 _12332_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_105_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12262_ _12336_/B _12262_/B vssd1 vssd1 vccd1 vccd1 _12280_/A sky130_fd_sc_hd__and2_1
XFILLER_0_120_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11213_ _11213_/A _11213_/B vssd1 vssd1 vccd1 vccd1 _11215_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12193_ _12283_/A _12193_/B vssd1 vssd1 vccd1 vccd1 _12195_/B sky130_fd_sc_hd__and2_1
X_11144_ _12537_/B2 _11131_/X _11143_/X _12710_/B2 _11142_/Y vssd1 vssd1 vccd1 vccd1
+ _11144_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07791__A1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07791__B2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11075_ _11076_/A _11076_/B vssd1 vssd1 vccd1 vccd1 _11075_/Y sky130_fd_sc_hd__nand2b_1
X_10026_ _10026_/A _10026_/B vssd1 vssd1 vccd1 vccd1 _10026_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__07703__A _12092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11977_ _06884_/A _09520_/X _12793_/A2 _11961_/A vssd1 vssd1 vccd1 vccd1 _11980_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11225__A _11225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13716_ _13717_/CLK _13716_/D vssd1 vssd1 vccd1 vccd1 hold291/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10928_ _10929_/A _10929_/B vssd1 vssd1 vccd1 vccd1 _10928_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13647_ _13649_/CLK _13647_/D vssd1 vssd1 vccd1 vccd1 hold237/A sky130_fd_sc_hd__dfxtp_1
X_10859_ _10302_/B _10857_/X _10858_/X _10856_/Y vssd1 vssd1 vccd1 vccd1 _10860_/B
+ sky130_fd_sc_hd__o211a_4
XFILLER_0_26_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08534__A _08951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13578_ _13605_/A hold248/X vssd1 vssd1 vccd1 vccd1 _13733_/D sky130_fd_sc_hd__and2_1
XFILLER_0_54_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10602__A1 _10457_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12529_ hold273/A _12786_/B1 _12595_/B _12528_/Y _12748_/B1 vssd1 vssd1 vccd1 vccd1
+ _12529_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_42_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11158__A2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06989__A _07110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09365__A _10507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09771__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09740_ _09740_/A _09740_/B vssd1 vssd1 vccd1 vccd1 _09808_/A sky130_fd_sc_hd__xnor2_4
X_06952_ reg2_val[10] _06980_/B vssd1 vssd1 vccd1 vccd1 _06952_/X sky130_fd_sc_hd__and2_2
XFILLER_0_94_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10118__B1 _11423_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
.ends

