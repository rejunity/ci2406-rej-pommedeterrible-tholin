// This is the unpowered netlist.
module ci2406_z80 (rst_n,
    wb_clk_i,
    io_in,
    io_oeb,
    io_out);
 input rst_n;
 input wb_clk_i;
 input [35:0] io_in;
 output [35:0] io_oeb;
 output [35:0] io_out;

 wire net185;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net186;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net187;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net217;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire clknet_0_wb_clk_i;
 wire clknet_2_0__leaf_wb_clk_i;
 wire clknet_2_1__leaf_wb_clk_i;
 wire clknet_2_2__leaf_wb_clk_i;
 wire clknet_2_3__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \z80.tv80s.di_reg[0] ;
 wire \z80.tv80s.di_reg[1] ;
 wire \z80.tv80s.di_reg[2] ;
 wire \z80.tv80s.di_reg[3] ;
 wire \z80.tv80s.di_reg[4] ;
 wire \z80.tv80s.di_reg[5] ;
 wire \z80.tv80s.di_reg[6] ;
 wire \z80.tv80s.di_reg[7] ;
 wire \z80.tv80s.i_tv80_core.ACC[0] ;
 wire \z80.tv80s.i_tv80_core.ACC[1] ;
 wire \z80.tv80s.i_tv80_core.ACC[2] ;
 wire \z80.tv80s.i_tv80_core.ACC[3] ;
 wire \z80.tv80s.i_tv80_core.ACC[4] ;
 wire \z80.tv80s.i_tv80_core.ACC[5] ;
 wire \z80.tv80s.i_tv80_core.ACC[6] ;
 wire \z80.tv80s.i_tv80_core.ACC[7] ;
 wire \z80.tv80s.i_tv80_core.ALU_Op_r[0] ;
 wire \z80.tv80s.i_tv80_core.ALU_Op_r[1] ;
 wire \z80.tv80s.i_tv80_core.ALU_Op_r[2] ;
 wire \z80.tv80s.i_tv80_core.ALU_Op_r[3] ;
 wire \z80.tv80s.i_tv80_core.Alternate ;
 wire \z80.tv80s.i_tv80_core.Ap[0] ;
 wire \z80.tv80s.i_tv80_core.Ap[1] ;
 wire \z80.tv80s.i_tv80_core.Ap[2] ;
 wire \z80.tv80s.i_tv80_core.Ap[3] ;
 wire \z80.tv80s.i_tv80_core.Ap[4] ;
 wire \z80.tv80s.i_tv80_core.Ap[5] ;
 wire \z80.tv80s.i_tv80_core.Ap[6] ;
 wire \z80.tv80s.i_tv80_core.Ap[7] ;
 wire \z80.tv80s.i_tv80_core.Arith16_r ;
 wire \z80.tv80s.i_tv80_core.Auto_Wait_t1 ;
 wire \z80.tv80s.i_tv80_core.Auto_Wait_t2 ;
 wire \z80.tv80s.i_tv80_core.BTR_r ;
 wire \z80.tv80s.i_tv80_core.BusA[0] ;
 wire \z80.tv80s.i_tv80_core.BusA[1] ;
 wire \z80.tv80s.i_tv80_core.BusA[2] ;
 wire \z80.tv80s.i_tv80_core.BusA[3] ;
 wire \z80.tv80s.i_tv80_core.BusA[4] ;
 wire \z80.tv80s.i_tv80_core.BusA[5] ;
 wire \z80.tv80s.i_tv80_core.BusA[6] ;
 wire \z80.tv80s.i_tv80_core.BusA[7] ;
 wire \z80.tv80s.i_tv80_core.BusAck ;
 wire \z80.tv80s.i_tv80_core.BusB[0] ;
 wire \z80.tv80s.i_tv80_core.BusB[1] ;
 wire \z80.tv80s.i_tv80_core.BusB[2] ;
 wire \z80.tv80s.i_tv80_core.BusB[3] ;
 wire \z80.tv80s.i_tv80_core.BusB[4] ;
 wire \z80.tv80s.i_tv80_core.BusB[5] ;
 wire \z80.tv80s.i_tv80_core.BusB[6] ;
 wire \z80.tv80s.i_tv80_core.BusB[7] ;
 wire \z80.tv80s.i_tv80_core.BusReq_s ;
 wire \z80.tv80s.i_tv80_core.F[0] ;
 wire \z80.tv80s.i_tv80_core.F[1] ;
 wire \z80.tv80s.i_tv80_core.F[2] ;
 wire \z80.tv80s.i_tv80_core.F[3] ;
 wire \z80.tv80s.i_tv80_core.F[4] ;
 wire \z80.tv80s.i_tv80_core.F[5] ;
 wire \z80.tv80s.i_tv80_core.F[6] ;
 wire \z80.tv80s.i_tv80_core.F[7] ;
 wire \z80.tv80s.i_tv80_core.Fp[0] ;
 wire \z80.tv80s.i_tv80_core.Fp[1] ;
 wire \z80.tv80s.i_tv80_core.Fp[2] ;
 wire \z80.tv80s.i_tv80_core.Fp[3] ;
 wire \z80.tv80s.i_tv80_core.Fp[4] ;
 wire \z80.tv80s.i_tv80_core.Fp[5] ;
 wire \z80.tv80s.i_tv80_core.Fp[6] ;
 wire \z80.tv80s.i_tv80_core.Fp[7] ;
 wire \z80.tv80s.i_tv80_core.Halt_FF ;
 wire \z80.tv80s.i_tv80_core.INT_s ;
 wire \z80.tv80s.i_tv80_core.IR[0] ;
 wire \z80.tv80s.i_tv80_core.IR[1] ;
 wire \z80.tv80s.i_tv80_core.IR[2] ;
 wire \z80.tv80s.i_tv80_core.IR[3] ;
 wire \z80.tv80s.i_tv80_core.IR[4] ;
 wire \z80.tv80s.i_tv80_core.IR[5] ;
 wire \z80.tv80s.i_tv80_core.IR[6] ;
 wire \z80.tv80s.i_tv80_core.IR[7] ;
 wire \z80.tv80s.i_tv80_core.ISet[0] ;
 wire \z80.tv80s.i_tv80_core.ISet[1] ;
 wire \z80.tv80s.i_tv80_core.ISet[2] ;
 wire \z80.tv80s.i_tv80_core.ISet[3] ;
 wire \z80.tv80s.i_tv80_core.IStatus[1] ;
 wire \z80.tv80s.i_tv80_core.IStatus[2] ;
 wire \z80.tv80s.i_tv80_core.I[0] ;
 wire \z80.tv80s.i_tv80_core.I[1] ;
 wire \z80.tv80s.i_tv80_core.I[2] ;
 wire \z80.tv80s.i_tv80_core.I[3] ;
 wire \z80.tv80s.i_tv80_core.I[4] ;
 wire \z80.tv80s.i_tv80_core.I[5] ;
 wire \z80.tv80s.i_tv80_core.I[6] ;
 wire \z80.tv80s.i_tv80_core.I[7] ;
 wire \z80.tv80s.i_tv80_core.IncDecZ ;
 wire \z80.tv80s.i_tv80_core.IntCycle ;
 wire \z80.tv80s.i_tv80_core.IntE ;
 wire \z80.tv80s.i_tv80_core.IntE_FF2 ;
 wire \z80.tv80s.i_tv80_core.NMICycle ;
 wire \z80.tv80s.i_tv80_core.NMI_s ;
 wire \z80.tv80s.i_tv80_core.No_BTR ;
 wire \z80.tv80s.i_tv80_core.Oldnmi_n ;
 wire \z80.tv80s.i_tv80_core.PC[0] ;
 wire \z80.tv80s.i_tv80_core.PC[10] ;
 wire \z80.tv80s.i_tv80_core.PC[11] ;
 wire \z80.tv80s.i_tv80_core.PC[12] ;
 wire \z80.tv80s.i_tv80_core.PC[13] ;
 wire \z80.tv80s.i_tv80_core.PC[14] ;
 wire \z80.tv80s.i_tv80_core.PC[15] ;
 wire \z80.tv80s.i_tv80_core.PC[1] ;
 wire \z80.tv80s.i_tv80_core.PC[2] ;
 wire \z80.tv80s.i_tv80_core.PC[3] ;
 wire \z80.tv80s.i_tv80_core.PC[4] ;
 wire \z80.tv80s.i_tv80_core.PC[5] ;
 wire \z80.tv80s.i_tv80_core.PC[6] ;
 wire \z80.tv80s.i_tv80_core.PC[7] ;
 wire \z80.tv80s.i_tv80_core.PC[8] ;
 wire \z80.tv80s.i_tv80_core.PC[9] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[1] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[2] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[3] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[4] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[5] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[6] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[7] ;
 wire \z80.tv80s.i_tv80_core.PreserveC_r ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[0] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[2] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[4] ;
 wire \z80.tv80s.i_tv80_core.RegAddrA_r[0] ;
 wire \z80.tv80s.i_tv80_core.RegAddrA_r[1] ;
 wire \z80.tv80s.i_tv80_core.RegAddrA_r[2] ;
 wire \z80.tv80s.i_tv80_core.RegAddrB_r[0] ;
 wire \z80.tv80s.i_tv80_core.RegAddrB_r[1] ;
 wire \z80.tv80s.i_tv80_core.RegAddrB_r[2] ;
 wire \z80.tv80s.i_tv80_core.RegAddrC[0] ;
 wire \z80.tv80s.i_tv80_core.RegAddrC[1] ;
 wire \z80.tv80s.i_tv80_core.RegAddrC[2] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[0] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[10] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[11] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[12] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[13] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[14] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[15] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[1] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[2] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[3] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[4] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[5] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[6] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[7] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[8] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[9] ;
 wire \z80.tv80s.i_tv80_core.SP[0] ;
 wire \z80.tv80s.i_tv80_core.SP[10] ;
 wire \z80.tv80s.i_tv80_core.SP[11] ;
 wire \z80.tv80s.i_tv80_core.SP[12] ;
 wire \z80.tv80s.i_tv80_core.SP[13] ;
 wire \z80.tv80s.i_tv80_core.SP[14] ;
 wire \z80.tv80s.i_tv80_core.SP[15] ;
 wire \z80.tv80s.i_tv80_core.SP[1] ;
 wire \z80.tv80s.i_tv80_core.SP[2] ;
 wire \z80.tv80s.i_tv80_core.SP[3] ;
 wire \z80.tv80s.i_tv80_core.SP[4] ;
 wire \z80.tv80s.i_tv80_core.SP[5] ;
 wire \z80.tv80s.i_tv80_core.SP[6] ;
 wire \z80.tv80s.i_tv80_core.SP[7] ;
 wire \z80.tv80s.i_tv80_core.SP[8] ;
 wire \z80.tv80s.i_tv80_core.SP[9] ;
 wire \z80.tv80s.i_tv80_core.Save_ALU_r ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[0] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[10] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[11] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[12] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[13] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[14] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[15] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[1] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[2] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[3] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[4] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[5] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[6] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[7] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[8] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[9] ;
 wire \z80.tv80s.i_tv80_core.XY_Ind ;
 wire \z80.tv80s.i_tv80_core.XY_State[0] ;
 wire \z80.tv80s.i_tv80_core.XY_State[1] ;
 wire \z80.tv80s.i_tv80_core.Z16_r ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[0] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][7] ;
 wire \z80.tv80s.i_tv80_core.mcycles[1] ;
 wire \z80.tv80s.i_tv80_core.mcycles[2] ;
 wire \z80.tv80s.i_tv80_core.mcycles[4] ;
 wire \z80.tv80s.i_tv80_core.mcycles[5] ;
 wire \z80.tv80s.i_tv80_core.ts[0] ;
 wire \z80.tv80s.i_tv80_core.ts[1] ;
 wire \z80.tv80s.i_tv80_core.ts[2] ;
 wire \z80.tv80s.i_tv80_core.ts[3] ;
 wire \z80.tv80s.i_tv80_core.ts[4] ;
 wire \z80.tv80s.i_tv80_core.ts[5] ;
 wire \z80.tv80s.i_tv80_core.ts[6] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0380_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_2851_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_2927_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(\z80.tv80s.i_tv80_core.INT_s ));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(\z80.tv80s.i_tv80_core.INT_s ));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\z80.tv80s.i_tv80_core.INT_s ));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(\z80.tv80s.i_tv80_core.INT_s ));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(\z80.tv80s.i_tv80_core.INT_s ));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(\z80.tv80s.i_tv80_core.INT_s ));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0562_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_0551_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_0563_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(\z80.tv80s.i_tv80_core.IncDecZ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_1765_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_1795_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(\z80.tv80s.i_tv80_core.NMICycle ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_1244_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_1455_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_2079_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_2191_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_2383_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_2706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2946__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2951__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2952__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__2955__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__2956__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__2957__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__2958__A (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2959__A (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2960__A (.DIODE(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2961__A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2968__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__2973__A (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2975__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2976__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2981__A (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2982__A (.DIODE(\z80.tv80s.i_tv80_core.Arith16_r ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2983__A (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2984__A (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2985__A (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2986__A (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2987__A (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2988__A (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2991__A (.DIODE(\z80.tv80s.i_tv80_core.PC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3002__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__3010__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3010__B (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3013__A (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3013__B (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3014__B (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3016__A (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3017__A (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3018__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3021__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3033__A (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3036__A2 (.DIODE(_2773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3041__A1 (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3042__B (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3048__A1 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3053__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3054__C_N (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3058__A (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3058__B (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3059__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__3059__B (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3062__A (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3066__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3066__C (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3068__A (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3068__B (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3069__B (.DIODE(_2812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3071__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__3071__B (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3072__A_N (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__3072__B (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3077__A1 (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3079__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3079__B1 (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3084__B1 (.DIODE(_2828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3094__A (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3102__A (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3103__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3106__D (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3108__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3109__B (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3110__B (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3111__A3 (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3117__B1 (.DIODE(_2860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3119__A3 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3121__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__3121__C (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3122__A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3122__B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3126__A2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3127__C (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3129__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3132__A (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3132__B (.DIODE(_2773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3134__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3135__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3136__A (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3143__B (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3144__A (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3147__A1 (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3147__A3 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3148__D (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3149__A (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3149__B (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3150__B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3151__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3152__A2 (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3153__A1 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3153__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__3159__A1 (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3161__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3162__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3162__B (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3163__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3163__A2 (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3163__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3164__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3164__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3165__B (.DIODE(_2828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3169__B (.DIODE(_2860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3170__A (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3171__A (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3175__A (.DIODE(_2773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3175__C (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3179__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3190__A1 (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3190__A2 (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3191__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__3191__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3192__B (.DIODE(_2860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3193__B (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__3193__C (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3199__A2 (.DIODE(_2860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3199__C1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3201__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3204__A_N (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3204__B (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3205__A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3206__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3206__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3207__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3207__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__B (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3210__C (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3212__A1 (.DIODE(_2843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3212__A2 (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3213__B (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3214__B (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3215__A (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3215__B (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3216__B1 (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3217__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3220__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__3221__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3221__A2 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3221__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3222__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3222__A2 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3222__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3223__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3225__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3225__B (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3226__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3226__B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__3227__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3229__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3229__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__3232__B (.DIODE(_2840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3233__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3236__A0 (.DIODE(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3236__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3238__A (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3240__B (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3241__C (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3242__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3243__S (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3245__D1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__3247__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3247__B (.DIODE(_0415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3250__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3250__B (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3250__C (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3251__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3251__C1 (.DIODE(_2939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3252__A (.DIODE(\z80.tv80s.i_tv80_core.IntCycle ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3252__B (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__3254__A (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3256__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__3256__A3 (.DIODE(_0415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3257__A2 (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3258__A2 (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3259__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3260__B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3263__B1 (.DIODE(_2840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3264__A (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3265__A_N (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3265__D (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3268__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3271__B1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__3274__A (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3274__B (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3276__C (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3276__D (.DIODE(_2939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3277__A (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3278__B (.DIODE(_2812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3278__C (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3280__A (.DIODE(_2773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__B (.DIODE(_0415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3284__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3286__B (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3287__A (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3288__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3291__B1 (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3292__A1 (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3292__A2 (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3293__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3295__A_N (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3296__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__3296__A2 (.DIODE(_0466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3296__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3297__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3297__A2 (.DIODE(_0466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3297__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3299__A (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3299__B (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3300__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3301__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3302__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__3304__A1 (.DIODE(_2840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__A1 (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__B1 (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3309__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__3310__A1 (.DIODE(_2860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3310__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3312__A1 (.DIODE(_0377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3312__B2 (.DIODE(\z80.tv80s.i_tv80_core.ISet[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3312__C1 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3313__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3314__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3314__B2 (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3315__A1_N (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3317__A2 (.DIODE(_0415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3318__A (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3319__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3320__A (.DIODE(\z80.tv80s.i_tv80_core.ISet[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3321__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3322__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__3323__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3326__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3327__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3329__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3335__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3336__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__3336__A3 (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3338__C1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3339__A1 (.DIODE(\z80.tv80s.i_tv80_core.ISet[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3339__D1 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3342__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__3344__A0 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__3347__A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__3348__A (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3348__B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__3349__A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__3349__B (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3350__A (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__3350__B (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__3350__C (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3352__A (.DIODE(_0446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3353__A (.DIODE(_0446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3354__A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3354__B (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3356__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__3356__B (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3356__C (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3357__A1 (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3359__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3359__B (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3360__A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3362__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__3362__B (.DIODE(\z80.tv80s.i_tv80_core.BusReq_s ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3362__C (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3362__D (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3363__A (.DIODE(_0446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3363__D_N (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3364__A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__3366__A_N (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__3368__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3370__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__3370__B (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3377__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__3377__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__3378__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__3378__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__A1 (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__A2 (.DIODE(_2828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__C1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3380__A_N (.DIODE(_2828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3381__A1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__3381__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3382__B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__3383__B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__3384__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3384__A2 (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3384__C1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3385__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3385__B (.DIODE(_2828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__C (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3387__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3387__B (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3387__C (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3389__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3389__D_N (.DIODE(_0551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3391__A1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3394__A1 (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3394__A2 (.DIODE(_0415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__A_N (.DIODE(\z80.tv80s.i_tv80_core.NMICycle ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__C (.DIODE(\z80.tv80s.i_tv80_core.IntCycle ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3397__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3398__B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3399__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3400__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3401__A1 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3403__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3403__B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3404__A2 (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3405__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3405__B (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3406__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3406__B2 (.DIODE(_0563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3407__A2 (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3407__A3 (.DIODE(_0415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3408__A2 (.DIODE(_2939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3408__B1 (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3409__A1 (.DIODE(\z80.tv80s.i_tv80_core.NMICycle ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3409__B1 (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3410__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__3412__A (.DIODE(_2773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3413__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3414__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3415__A1 (.DIODE(\z80.tv80s.i_tv80_core.ISet[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3415__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3415__A3 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3416__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3417__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3418__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3418__A2 (.DIODE(_2860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3418__A3 (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3419__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__3420__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3420__B (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3423__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3423__B2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__A1 (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__A3 (.DIODE(_0563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__B2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3425__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3426__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3426__C (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3431__A1 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3433__A (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__3433__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3433__C (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__B (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__C (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__D (.DIODE(_0563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3436__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3436__B (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3437__A2 (.DIODE(_2843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3437__B1 (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3438__B1 (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3440__C1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__A1 (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3442__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3444__C1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__B (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__A1 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3450__A2 (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__A2 (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3452__A1 (.DIODE(_2860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3452__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3453__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3453__C1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3454__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__3454__B (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__A3 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3457__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3457__B (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__A1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__A2 (.DIODE(_2840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__B1 (.DIODE(_2711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__A1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__A3 (.DIODE(_2843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__3461__B (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3462__A1 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__3462__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3463__B (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__A2 (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3465__A1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3465__A2 (.DIODE(_0613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3465__B1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3467__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3467__B (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__A2 (.DIODE(_2843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__B1 (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__D1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3469__B (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3471__A3 (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__A1_N (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__A2_N (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__B2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__A1 (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__C1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__B1 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3476__A2 (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__A2 (.DIODE(_2812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__C1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__D1 (.DIODE(_2939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3484__C (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__B (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3488__B (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3489__B2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__A2 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__B1 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__S (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3496__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3499__A1 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__A3 (.DIODE(\z80.tv80s.i_tv80_core.IncDecZ ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3503__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__3503__B (.DIODE(\z80.tv80s.i_tv80_core.BusReq_s ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3503__C (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__B (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__C_N (.DIODE(_0446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__A3 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__B (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3507__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3507__B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3507__C (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3508__B (.DIODE(\z80.tv80s.i_tv80_core.INT_s ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__A (.DIODE(_0551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__B (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3511__B (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__C (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3513__A (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3513__B (.DIODE(\z80.tv80s.i_tv80_core.IntE_FF2 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3514__A1 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__B (.DIODE(_0551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__C (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__A1 (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__A2 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__B1 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__C (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__D (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3522__A1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3524__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__B (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__3526__B (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__A (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__A1 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__B (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__C (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__B (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__C (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__B (.DIODE(\z80.tv80s.i_tv80_core.ts[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__C (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__B (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__C (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3541__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__B (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3544__A2 (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3548__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__A1 (.DIODE(_2840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__A2 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__B1 (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__A2 (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3556__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__3558__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__A1 (.DIODE(_2756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__C1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3567__B (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__A2 (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__A2 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__A1 (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3573__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__A1 (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__A1 (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3581__A1 (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3581__C1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__B1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3585__A1 (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3585__C1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__A (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__C (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__B (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3591__A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__3591__B (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3592__B (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__A2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3594__A2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__S0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__S1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3596__A2 (.DIODE(_2714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__B (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__C (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3600__A (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3600__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3601__B (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__A (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__C (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__C (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3604__A (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3604__B (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3606__A (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3606__B (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3607__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3609__A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3609__C1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__C1 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3611__A (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3611__B (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3613__A (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3613__B (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__A (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__B (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3617__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3622__B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3623__A (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__A (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3627__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3630__B (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__A3 (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3644__C (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__D (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__A (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3649__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3649__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__A (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__A (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3652__C (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3653__A2 (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3653__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__3653__C1 (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3660__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3661__B2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3663__A2 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3665__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3665__A2 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3666__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3667__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3668__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3669__S (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__B (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__B (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__C1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__C1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__A (.DIODE(_0809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__A1 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__A_N (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3680__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__B1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3690__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3690__A3 (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__B (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3694__C (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__B2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3698__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3698__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3698__B1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__B1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__A (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__B (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__S (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3706__A0 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__A2 (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__A (.DIODE(_0466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__C1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3713__A (.DIODE(_2843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__B (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__A2 (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3721__A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3721__C1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__C1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3726__C1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__C1 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3733__A (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3734__A1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3734__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3736__A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3736__B1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3737__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3738__S (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__S (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__C1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__C1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__A (.DIODE(_0809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__A1 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3748__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__B1 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__B1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3764__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__A0 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__B (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__B2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__A0 (.DIODE(_2735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__A (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__A2 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__B1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__A2 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__S (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__A2 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__B1 (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3793__C (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__C (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__B (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__C (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__A2 (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__B1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__A3 (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__B1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__A3 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__B (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__C (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__B1 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__A (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__A0 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__A (.DIODE(_0967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__A2 (.DIODE(_0967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__C1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__S0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__S1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__S (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__A (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__B (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__B1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3847__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__A0 (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__A1 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3871__B1 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__A1 (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3877__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__S0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3879__S1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__S (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__A2 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__B1 (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__A2 (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__B1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__A1 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3887__A1 (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__A3 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__A (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__A (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__S (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3919__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3923__B2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__A0 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__A2 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3928__A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__S0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__S1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3930__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3931__S (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3932__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3933__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__A3 (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__S (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__A (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__A1 (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__A1 (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__B2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3959__A (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__A2 (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3963__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__C1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3967__A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3967__C1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__A (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3971__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__S0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__S1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__S (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__S (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__C1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__C1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__A1 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3993__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__3996__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3999__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__3999__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4000__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4004__A3 (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__B (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4007__A0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4009__B (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4010__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__S (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__A (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__A (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__B (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__B2 (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__A0 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4032__A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__S0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__S1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__S (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__B (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__C (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4039__B (.DIODE(_2812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__A2 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__B (.DIODE(_2773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__C (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__A1 (.DIODE(_2939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4051__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__A1 (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__A1 (.DIODE(_2840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__A2 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__B1 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4059__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4059__C1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__C1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__A1 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__B1 (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__A4 (.DIODE(_2939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__B1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4068__A1 (.DIODE(_2773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4068__A3 (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4070__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__4070__B (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__A1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__B2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__4074__A (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4074__B (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4074__C (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4074__D_N (.DIODE(_1204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4078__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__4079__A1 (.DIODE(_2939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4080__A2 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__B1 (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__A3 (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__C1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__4086__A2 (.DIODE(_2860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4086__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__B2 (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4089__A2 (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4089__B2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__B2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__B2 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4092__A2 (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__A2 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__A1 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__B1 (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4100__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__4102__B2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__4103__B2 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__A (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__B (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__C (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__D_N (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__S (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4109__S (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4110__S (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4111__S (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4112__S (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4113__S (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4114__S (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4115__S (.DIODE(_1236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4116__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4116__B (.DIODE(_2814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__4120__B1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__A (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__4123__A0 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4124__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__4124__D (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4126__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__B1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__4128__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__4128__A2 (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__A1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4133__S0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4133__S1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4136__B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__4148__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4149__B1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4153__A2 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4153__B1 (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__A2 (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4155__B1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4162__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4163__C1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__S0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__S1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__A2 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__B1 (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__A2 (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4170__B1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4177__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4178__A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4178__C1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4179__S0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4182__A2 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4182__B1 (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4184__A2 (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4185__B1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4190__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4192__S0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__A2 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__B1 (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4200__A2 (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4201__B1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4208__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4209__A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4210__S0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4210__S1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4213__A2 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4213__B1 (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4215__A2 (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4216__B1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4223__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__S0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__S1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4229__A2 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4229__B1 (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4230__A2 (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4231__B1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__4239__A (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4240__A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4241__S0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__A2 (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__B1 (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__A2 (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4248__B1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__A1 (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__B1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__S (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4257__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4257__C1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__C1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__A (.DIODE(_0809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4260__A1 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4264__S (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__S (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4266__S (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__S (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__S (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__S (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4270__S (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__S (.DIODE(_1374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4272__B (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4273__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__S (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__S (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__S (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4287__S (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4288__S (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4289__S (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__S (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4291__S (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__S (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4294__S (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4295__S (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__S (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__S (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__S (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4299__S (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__S (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__S (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4303__S (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__S (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__S (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__S (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4307__S (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4308__S (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__S (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__S (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4312__S (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__S (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4314__S (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4315__S (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__S (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__S (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4318__S (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4320__S (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__S (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4322__S (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__S (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__S (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4325__S (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__S (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__S (.DIODE(_1381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__S (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__S (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4331__S (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__S (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__S (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__S (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4335__S (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__S (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4338__S (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__S (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4340__S (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4341__S (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__S (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__S (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__S (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__S (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4347__S (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4348__S (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4349__S (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4350__S (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__S (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__S (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__S (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__S (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4356__S (.DIODE(_1385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4357__S (.DIODE(_1385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4358__S (.DIODE(_1385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4359__S (.DIODE(_1385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__S (.DIODE(_1385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__S (.DIODE(_1385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__S (.DIODE(_1385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4363__S (.DIODE(_1385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4365__S (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__S (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4367__S (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__S (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__S (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4370__S (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__S (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4372__S (.DIODE(_1386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__B (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__4378__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4380__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__4382__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4382__A2 (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4382__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__4383__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4383__A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__4383__A3 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__A1 (.DIODE(_2773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__4387__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__C1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__4391__A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4391__B (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4393__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__4393__C1 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4394__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__A (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4396__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__4396__B1 (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__A2 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__B1 (.DIODE(_0377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__A2 (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__B1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__A1 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__A2 (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__B1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4403__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__A1 (.DIODE(_1204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__A2 (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__B1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4405__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__B (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__A1 (.DIODE(_2773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__A2 (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__A3 (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__A1 (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__A1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__B2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__B (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__A1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__A2 (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__4414__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4417__C (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__B1 (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__B2 (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__A1 (.DIODE(_1411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__B1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4424__A (.DIODE(_2773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__A2 (.DIODE(_2812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__A1 (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__A2 (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__B1 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__B2 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__B (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__C (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__A2 (.DIODE(_2843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__B2 (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__B2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__A1 (.DIODE(_0377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__A2 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__B2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__B (.DIODE(_2939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__A1 (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__A1 (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__A2 (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__B (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__C1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__A2 (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__A_N (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__C (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__D (.DIODE(\z80.tv80s.i_tv80_core.ISet[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__B1 (.DIODE(_0563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__B2 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__A1 (.DIODE(\z80.tv80s.i_tv80_core.NMICycle ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__A2 (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__B1 (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__A1 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__A2 (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__A1 (.DIODE(_2703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__A1 (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__D (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__B2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__S0 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__S1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__S0 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__S1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__A2 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__A3 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__A (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__B (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4474__A (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__4474__B (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__B (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__A1 (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__C1 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__4478__A (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__4479__A (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__B2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__A0 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__S (.DIODE(_1465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__B (.DIODE(_2828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__C (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__A (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__A2 (.DIODE(_1465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__A3 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__C1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__S0 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__S1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__S0 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__S1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__A0 (.DIODE(\z80.tv80s.i_tv80_core.SP[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__S (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__A (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__A2 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__B2 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__A0 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__S (.DIODE(_1465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4507__B (.DIODE(_2735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__S0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__S1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__S0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__S1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__A (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__A2 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__B2 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4519__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__A0 (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__S (.DIODE(_1465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__S0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__S1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__S0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__S1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__A (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4532__A0 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__A0 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__S (.DIODE(_1465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__B (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__S0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__S1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__S0 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__S1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__A1 (.DIODE(_1536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__A (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__A0 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__A0 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__S (.DIODE(_1465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__A_N (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__S0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__S1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__S0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__S1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__A1 (.DIODE(_1551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__A (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__A0 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__A0 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__S (.DIODE(_1465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__S0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__S1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__S0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__S1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__A1 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__A (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__A1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__A2 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__B2 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__A0 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__S (.DIODE(_1465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__A1 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__S0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__S1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__S0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__S1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__A1 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__A2 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__B2 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__S (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__A0 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__S (.DIODE(_1465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__S0 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__S1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__S0 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__S1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4603__A1 (.DIODE(_1593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__B (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__A (.DIODE(_2773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__B (.DIODE(_2812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__C (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4619__A1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4619__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__A1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__B1 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__A2 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__B1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__4623__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__S0 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__S1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__S0 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__S1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__A1 (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__A2 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__B2 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__B1 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__A2 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__S0 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__S1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__S0 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__S1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4640__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__A2 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__B2 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__B1 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__A1 (.DIODE(_2735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__A2 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__S0 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__S1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__S0 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__S1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__A1 (.DIODE(_1644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__A2 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__B2 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__B1 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__A1 (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__A2 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__S0 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__S1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__S0 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__S1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__A1 (.DIODE(_1657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__A2 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4678__B2 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__B1 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__A1 (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__A2 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4682__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__S0 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__S1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__S0 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__S1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__A1 (.DIODE(_1671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__C1 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__A1 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__A2 (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__S0 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__S1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__S0 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__S1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__A1 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__A2 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__B2 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__B1 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__A1 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__A2 (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__S0 (.DIODE(\z80.tv80s.i_tv80_core.RegAddrC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__S1 (.DIODE(\z80.tv80s.i_tv80_core.RegAddrC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__S0 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__S1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__S (.DIODE(\z80.tv80s.i_tv80_core.RegAddrC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__A2 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__B2 (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__B1 (.DIODE(_1610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__A1 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__A2 (.DIODE(_1611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__D (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__A2 (.DIODE(_2860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__A2 (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__A3 (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__A (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__B (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__B (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__A1 (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__A2 (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__A1 (.DIODE(_0377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__A1_N (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__B1 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__B2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__4748__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__A2_N (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__A1 (.DIODE(_0466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__B (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__A1 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__A2 (.DIODE(_2812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__C1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__A (.DIODE(_0384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__B (.DIODE(_0466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__A (.DIODE(\z80.tv80s.i_tv80_core.NMICycle ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__B (.DIODE(\z80.tv80s.i_tv80_core.IntCycle ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__B (.DIODE(\z80.tv80s.i_tv80_core.IntCycle ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4772__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__A1 (.DIODE(_2702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__A2 (.DIODE(_2812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__A (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4777__B (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__A0 (.DIODE(\z80.tv80s.i_tv80_core.PC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__S (.DIODE(_0446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__B (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__A1 (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__C1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__B2 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__C1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__A1 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__A2 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4782__B1 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4787__S (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__A1 (.DIODE(_1765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__A2 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__B1 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4791__B2 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__A0 (.DIODE(\z80.tv80s.i_tv80_core.PC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__S (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__C (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__A2 (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__B2 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__A1 (.DIODE(\z80.tv80s.i_tv80_core.SP[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4799__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4799__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4802__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__S (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__A1 (.DIODE(_1780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__C (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__S (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__C1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__A1 (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__A2 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__B (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__S (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__A1 (.DIODE(_1795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__B (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__S (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__C1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__A1 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__A2 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4834__S (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__A1 (.DIODE(_1809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__B (.DIODE(_1536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__S (.DIODE(_0446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__A0 (.DIODE(_1536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__B1 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__B2 (.DIODE(_1536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__C1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__A1 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__A2 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__S (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__A1 (.DIODE(_1822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__B (.DIODE(_1551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__S (.DIODE(_0446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__A0 (.DIODE(_1551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__4855__B1 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__B2 (.DIODE(_1551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__C1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__A1 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__A2 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__S (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__A1 (.DIODE(_1836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__B (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__S (.DIODE(_0446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__A0 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__S (.DIODE(_0444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__B1 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__B2 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__C1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__A1 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__A2 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__S (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__A1 (.DIODE(_1849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__B (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__S (.DIODE(_0446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__A0 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__B2 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__C1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__C1 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__A1 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__A2 (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__S (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4894__A1 (.DIODE(_1864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4894__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__B (.DIODE(_1593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__A (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__B (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__B2 (.DIODE(_1593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__A0 (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__S (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__A0 (.DIODE(_1593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__A0 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__S (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__B2 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__A2 (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__A1 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__S (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__A1 (.DIODE(_1879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__B (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__A (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__B (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4913__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4913__B2 (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__A0 (.DIODE(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__S (.DIODE(_0446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__B (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4916__A1 (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4916__C1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__A (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__B (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__B1 (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__A1 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4922__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4922__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__4925__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__A1 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__S (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__4928__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__A (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4929__B (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4930__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__S (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__A0 (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__S (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__B2 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__A (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__A1 (.DIODE(_1909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__S (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4943__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4943__B (.DIODE(_1644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__A (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__B (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4945__B2 (.DIODE(_1644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__A0 (.DIODE(\z80.tv80s.i_tv80_core.PC[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__S (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__A0 (.DIODE(_1644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__A0 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__S (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__B2 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__4957__A1 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__S (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__B (.DIODE(_1657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__A (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__B (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4961__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4961__B2 (.DIODE(_1657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__S (.DIODE(_0446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__B (.DIODE(_1657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__A1 (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__C1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4967__A (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4967__B (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4968__B1 (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__A1 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__A1 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__S (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__B (.DIODE(_1671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__A (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__B (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__B2 (.DIODE(_1671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__S (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__A0 (.DIODE(_1671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__S (.DIODE(_0444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__A0 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__S (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__B2 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__A1 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__S (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__B (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__A (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__B (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__B2 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__S (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__A0 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__S (.DIODE(_0444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__A0 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__S (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__B2 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__A2 (.DIODE(_1744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__A1 (.DIODE(_1238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__A (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__S (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5007__A (.DIODE(_1238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__A (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__B (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__B1 (.DIODE(_1747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5010__S (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__S (.DIODE(_0444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__A0 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__S (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__A1 (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__B2 (.DIODE(_1749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__A2 (.DIODE(_1744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__A1 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__S (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__A2 (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__B1_N (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__A1 (.DIODE(_2711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__A1 (.DIODE(_2711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__A2 (.DIODE(\z80.tv80s.i_tv80_core.Arith16_r ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__C1 (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__A2 (.DIODE(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__B2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__A2 (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__B2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__B2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__D (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__B2 (.DIODE(_2711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__A_N (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__B (.DIODE(_2011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__D (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A1 (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5071__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__S (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__A0 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__A2 (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__B1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__B2 (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__A3 (.DIODE(_2891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__B2 (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__C1 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__A (.DIODE(_2027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__A (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__B (.DIODE(_2027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A1 (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A2 (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A3 (.DIODE(_2027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__A (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__A1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__B2 (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__B (.DIODE(_0415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__B1 (.DIODE(_0396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__A2 (.DIODE(_2805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__C1 (.DIODE(_2936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__B2 (.DIODE(_2920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__B1 (.DIODE(_2834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__A1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A (.DIODE(_2045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__B (.DIODE(_2046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__A (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__B (.DIODE(_2046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__A (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__A1 (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__A2 (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__B1 (.DIODE(_2027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5110__C1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__C1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__C1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__C1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__A (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__A2 (.DIODE(_0809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__B1 (.DIODE(_2045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5116__A (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__A1 (.DIODE(_0809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__B1 (.DIODE(_2046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__A (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__B (.DIODE(_2045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__A (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__B (.DIODE(_2045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__A2 (.DIODE(_2059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5125__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5125__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__A1 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__B2 (.DIODE(\z80.tv80s.i_tv80_core.PC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__A1 (.DIODE(\z80.tv80s.i_tv80_core.SP[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__B2 (.DIODE(\z80.tv80s.i_tv80_core.PC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__C1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__C1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__A (.DIODE(_0809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__A1 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__B1 (.DIODE(_2045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__A2 (.DIODE(_2046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5137__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__B2 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__C1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5143__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5143__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5143__C1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__A (.DIODE(_0809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__A1 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__B1 (.DIODE(_2045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__A1 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__A2 (.DIODE(_2046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__B2 (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__A1 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__B2 (.DIODE(\z80.tv80s.i_tv80_core.PC[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__C1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__C1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__C1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__C1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__S0 (.DIODE(_2045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__S1 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__A1 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__C1 (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__C1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__C1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__C1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__S0 (.DIODE(_2045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__S1 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5175__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__S (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__B2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__S (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__S (.DIODE(_2045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__S (.DIODE(_2045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5186__S (.DIODE(_0809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__B1 (.DIODE(_2125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__A1 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__B2 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__C1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__C1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__C1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__C1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__S0 (.DIODE(_2045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__S1 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__C1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__C1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__A (.DIODE(_0809_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A1 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__B1 (.DIODE(_2046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__A2 (.DIODE(_2045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__A1 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__A (.DIODE(_0446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5231__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__B2 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__A1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__B2 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__A2 (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__B1 (.DIODE(_1221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__A0 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__A1 (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__A2 (.DIODE(_2169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__B1_N (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__A1 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__A2 (.DIODE(_1204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__B1 (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__B (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__A (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__B (.DIODE(_1204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__A1 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__A2 (.DIODE(_1204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__B1 (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__A (.DIODE(_0760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__A (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__B (.DIODE(_1204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__C_N (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5252__A (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__A (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__A1 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__B2 (.DIODE(_2183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__A1 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__A1 (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__A1 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5274__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__A1 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__A1 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__A1 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__A1 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__B2 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__A2 (.DIODE(_1204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__B1 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__A1 (.DIODE(_1204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__S (.DIODE(_2213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__S (.DIODE(_2213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__S (.DIODE(_2213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__S (.DIODE(_2213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__S (.DIODE(_2213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5303__S (.DIODE(_2213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__S (.DIODE(_2213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__S (.DIODE(_2213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__A0 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__S (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__A0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__S (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__S (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__S (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__S (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__S (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__A0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__S (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__A0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__A1 (.DIODE(net853));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__S (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__A (.DIODE(net749));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__B (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__C1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__A (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A1 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__B2 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__B2 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__A2 (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__A2 (.DIODE(_0642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__A (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__A2 (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__B (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__B (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__A2 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__A3 (.DIODE(_2812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__B1 (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__A2 (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__B2 (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__A0 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__B (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__5352__A (.DIODE(_2243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__A2 (.DIODE(_2789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__A3 (.DIODE(_2812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__B1 (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__A1_N (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__B2 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__B (.DIODE(\z80.tv80s.i_tv80_core.ts[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__D (.DIODE(_0377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__A (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__A (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__C (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__A (.DIODE(_2252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__C (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__D (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__B (.DIODE(_2252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__C (.DIODE(_2254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__B2 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A1 (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A1 (.DIODE(\z80.tv80s.i_tv80_core.IntE_FF2 ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__S (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A2 (.DIODE(\z80.tv80s.i_tv80_core.Arith16_r ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__B1 (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__A1 (.DIODE(\z80.tv80s.i_tv80_core.Arith16_r ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5383__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__A (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__B1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__A2 (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__A (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__B (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__A (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__B (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__A (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__B (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__A (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__B (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__A (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__B (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__A (.DIODE(_2840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__C (.DIODE(_0587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__B1 (.DIODE(_2315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5426__B (.DIODE(_2315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__A1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__A1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__A2 (.DIODE(_2243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__A2 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__C1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__A2 (.DIODE(_2860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__B1 (.DIODE(_2254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__A2 (.DIODE(_2254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__A1 (.DIODE(_0967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__B1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__B1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__A1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__A2 (.DIODE(_2236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__C1 (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__B (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__B2 (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5452__B2 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5453__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__A2 (.DIODE(_2243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5455__A2 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__C1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__A2 (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5461__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5461__A2 (.DIODE(_2860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5462__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__B1 (.DIODE(_2254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__A2_N (.DIODE(_2254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__A0 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5466__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__B1 (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__A1 (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__A1 (.DIODE(_2011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__A (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__B (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__C (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__D (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__A (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__B (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__A0 (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__A0 (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__A0 (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__S (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__B1 (.DIODE(_2252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5486__A1 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5487__A0 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__A (.DIODE(\z80.tv80s.i_tv80_core.ts[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__S (.DIODE(_2374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__S (.DIODE(_2374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__S (.DIODE(_2374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__S (.DIODE(_2374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__S (.DIODE(_2374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__S (.DIODE(_2374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__S (.DIODE(_2374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__S (.DIODE(_2374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__A2 (.DIODE(_0546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__C1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__A3 (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__B1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__B (.DIODE(_2773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__B1 (.DIODE(_0385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__A1 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__B (.DIODE(_0613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__A2 (.DIODE(_0613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__A2 (.DIODE(_0374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__B1 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__A1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__B1 (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__B (.DIODE(_2387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__A (.DIODE(\z80.tv80s.i_tv80_core.PC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__S (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__S (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__S (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__S (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5522__A1 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__S (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__S (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__S (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5534__S (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__A1 (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5541__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5543__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__S (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__A2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__S (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__A1 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__S (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__5560__S (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__S (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5563__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5564__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__S (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__S (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__A1 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__S (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__S (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__S (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__A1 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__S (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__S (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__A1 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__S (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__S (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__S (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__A1 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5602__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5607__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__5609__S (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__S (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__S (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__A1 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__S (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__S (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__A1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__A1 (.DIODE(_0518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__B (.DIODE(_2387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__A1 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__B2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__A2 (.DIODE(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__A1_N (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__A1 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__5655__S (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__S (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__A2 (.DIODE(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__A4 (.DIODE(\z80.tv80s.i_tv80_core.PC[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__A1 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__5670__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__S (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5674__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5675__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__A1 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5677__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__B2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5685__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__B (.DIODE(_2471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5693__A2 (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__A1_N (.DIODE(_2377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__B (.DIODE(_2471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__5703__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__A1 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__S (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__5707__S (.DIODE(_2377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5710__A2 (.DIODE(\z80.tv80s.i_tv80_core.ts[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5710__B1 (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__A1 (.DIODE(_1237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__A2 (.DIODE(_2572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__A1 (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__B1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__B (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__A2 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__A1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__A2 (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5718__B2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__A1 (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__A2 (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__B2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__A1 (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__A2 (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__B2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__A1 (.DIODE(_0968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__A2 (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__B2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__A2 (.DIODE(_1536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__A1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__A2 (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__B2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__A2 (.DIODE(_1551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__A1 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__A2 (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5733__B2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__A1 (.DIODE(_1237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__A2 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__A1 (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__A2 (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__B2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5737__A1 (.DIODE(_1237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5737__A2 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5737__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__A1 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__A2 (.DIODE(_2570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5739__B2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__A2 (.DIODE(_2593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__B1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__B (.DIODE(_2593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__A2 (.DIODE(_1593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__A1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__A2 (.DIODE(_2593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5745__B2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__A2 (.DIODE(_1616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__A1 (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__A2 (.DIODE(_2593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__B2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__A1 (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__A2 (.DIODE(_2593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__B2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__A2 (.DIODE(_1644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__A1 (.DIODE(_0968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__A2 (.DIODE(_2593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__B2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__A2 (.DIODE(_1657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__A1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__A2 (.DIODE(_2593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__B2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__A2 (.DIODE(_1671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__A1 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__A2 (.DIODE(_2593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__B2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__B (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__C (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__B1_N (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__B (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__A2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__A3 (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__B1 (.DIODE(_2593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__B1 (.DIODE(_2593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__B2 (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5769__A3 (.DIODE(_2572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5769__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__A0 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__S (.DIODE(_2593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__S (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5774__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5778__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__A0 (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__A0 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__A0 (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__A0 (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__A0 (.DIODE(\z80.tv80s.i_tv80_core.F[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__A0 (.DIODE(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__A0 (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__A2 (.DIODE(_2243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__A1_N (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__A2_N (.DIODE(_2243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5796__A1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5798__A1_N (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5798__A2_N (.DIODE(_2243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5801__A1 (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__A1_N (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__A2_N (.DIODE(_2243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5806__A1 (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5811__A1 (.DIODE(_0968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__A1_N (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__A2_N (.DIODE(_2243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5814__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__A1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__A1 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__A1_N (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__A2_N (.DIODE(_2243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__A1 (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5828__A1_N (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5828__A2_N (.DIODE(_2243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__A1 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__A1 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5832__A0 (.DIODE(net808));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__A1 (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__B1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__A (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__A (.DIODE(_0671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5838__A (.DIODE(_0377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5838__B (.DIODE(_0379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__S (.DIODE(_2659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5841__A1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5842__A2 (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5842__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__S (.DIODE(_2659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5846__A1_N (.DIODE(_0845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__A1_N (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__S (.DIODE(_2659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5850__A1 (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__A2 (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5852__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5852__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5852__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__S (.DIODE(_2659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__A1 (.DIODE(_0968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__A2 (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__S (.DIODE(_2659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__A1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__A2 (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__B2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__S (.DIODE(_2659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5862__A1 (.DIODE(_1060_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5863__A2 (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5863__B2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5865__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5865__S (.DIODE(_2659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__A1 (.DIODE(_1092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5867__A2 (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5867__B2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__S (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__S (.DIODE(_2659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5870__A1 (.DIODE(_1162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5871__A2 (.DIODE(_2656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5871__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5873__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__A1 (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__B (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5876__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__5900__RESET_B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__RESET_B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__RESET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__RESET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__CLK (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__RESET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__RESET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6042__RESET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__RESET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__RESET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__RESET_B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__RESET_B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6051__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6052__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__RESET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6054__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6056__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__RESET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6058__RESET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6059__RESET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6060__RESET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__RESET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__RESET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6095__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__RESET_B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6125__RESET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__RESET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__RESET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6128__RESET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__RESET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6169__RESET_B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__6175__SET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__SET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6189__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6191__RESET_B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6192__RESET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__RESET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__RESET_B (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6195__RESET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__RESET_B (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__RESET_B (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6202__RESET_B (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__RESET_B (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__SET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__SET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6206__SET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6207__SET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6208__SET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6209__SET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6210__SET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6211__SET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__SET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6244__RESET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__RESET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6250__RESET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__RESET_B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__6293__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__6294__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__6295__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__6296__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__6297__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__6298__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout102_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout103_A (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_A (.DIODE(_0444_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(_0377_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(\z80.tv80s.i_tv80_core.ts[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(\z80.tv80s.i_tv80_core.ts[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net869));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(\z80.tv80s.i_tv80_core.RegAddrC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_A (.DIODE(\z80.tv80s.i_tv80_core.RegAddrC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_A (.DIODE(net805));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout53_A (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout54_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout57_A (.DIODE(_1744_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout58_A (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout59_A (.DIODE(_2377_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_A (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout61_A (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_A (.DIODE(_1739_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_A (.DIODE(_2572_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout67_A (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_A (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout71_A (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_A (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout74_A (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout76_A (.DIODE(_2471_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_A (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout78_A (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_A (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_A (.DIODE(_1237_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_A (.DIODE(_1238_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_A (.DIODE(_1743_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_A (.DIODE(_1743_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold181_A (.DIODE(\z80.tv80s.i_tv80_core.ts[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold268_A (.DIODE(\z80.tv80s.i_tv80_core.IncDecZ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold302_A (.DIODE(\z80.tv80s.i_tv80_core.NMICycle ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold338_A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold343_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold363_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold365_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold369_A (.DIODE(\z80.tv80s.i_tv80_core.ISet[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold373_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold384_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold388_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold396_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold400_A (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold408_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold410_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold419_A (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold435_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold482_A (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold484_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold494_A (.DIODE(\z80.tv80s.i_tv80_core.Arith16_r ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold506_A (.DIODE(\z80.tv80s.i_tv80_core.SP[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold508_A (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold512_A (.DIODE(\z80.tv80s.i_tv80_core.PC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold522_A (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold525_A (.DIODE(\z80.tv80s.i_tv80_core.PC[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold529_A (.DIODE(\z80.tv80s.i_tv80_core.IntCycle ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold531_A (.DIODE(\z80.tv80s.i_tv80_core.PC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold532_A (.DIODE(\z80.tv80s.i_tv80_core.BusReq_s ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold544_A (.DIODE(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold556_A (.DIODE(\z80.tv80s.i_tv80_core.ts[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold561_A (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold567_A (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold573_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold576_A (.DIODE(\z80.tv80s.i_tv80_core.F[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold588_A (.DIODE(\z80.tv80s.i_tv80_core.ISet[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold590_A (.DIODE(\z80.tv80s.i_tv80_core.RegAddrC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold591_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold593_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold594_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold595_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold596_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold598_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold599_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold601_A (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold603_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold604_A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold606_A (.DIODE(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold611_A (.DIODE(\z80.tv80s.i_tv80_core.IntE_FF2 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold614_A (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold616_A (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold619_A (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold623_A (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold629_A (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold630_A (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold631_A (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold632_A (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold635_A (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold636_A (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold637_A (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold647_A (.DIODE(\z80.tv80s.i_tv80_core.RegAddrC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold648_A (.DIODE(\z80.tv80s.i_tv80_core.RegAddrC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold649_A (.DIODE(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold651_A (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold652_A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold656_A (.DIODE(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_output21_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_output31_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_output32_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_output33_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_output34_A (.DIODE(net34));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _2946_ (.A(net142),
    .Y(_2697_));
 sky130_fd_sc_hd__inv_2 _2947_ (.A(net134),
    .Y(_2698_));
 sky130_fd_sc_hd__inv_2 _2948_ (.A(net135),
    .Y(_2699_));
 sky130_fd_sc_hd__inv_2 _2949_ (.A(net132),
    .Y(_2700_));
 sky130_fd_sc_hd__inv_2 _2950_ (.A(net130),
    .Y(_2701_));
 sky130_fd_sc_hd__inv_4 _2951_ (.A(net125),
    .Y(_2702_));
 sky130_fd_sc_hd__inv_6 _2952_ (.A(net122),
    .Y(_2703_));
 sky130_fd_sc_hd__inv_2 _2953_ (.A(\z80.tv80s.i_tv80_core.IR[7] ),
    .Y(_2704_));
 sky130_fd_sc_hd__inv_2 _2954_ (.A(net145),
    .Y(_2705_));
 sky130_fd_sc_hd__inv_2 _2955_ (.A(net149),
    .Y(_2706_));
 sky130_fd_sc_hd__inv_2 _2956_ (.A(net168),
    .Y(_2707_));
 sky130_fd_sc_hd__inv_2 _2957_ (.A(net163),
    .Y(_2708_));
 sky130_fd_sc_hd__inv_2 _2958_ (.A(\z80.tv80s.i_tv80_core.F[2] ),
    .Y(_2709_));
 sky130_fd_sc_hd__inv_2 _2959_ (.A(\z80.tv80s.i_tv80_core.F[0] ),
    .Y(_2710_));
 sky130_fd_sc_hd__inv_2 _2960_ (.A(\z80.tv80s.i_tv80_core.F[6] ),
    .Y(_2711_));
 sky130_fd_sc_hd__inv_2 _2961_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .Y(_2712_));
 sky130_fd_sc_hd__inv_2 _2962_ (.A(net656),
    .Y(_2713_));
 sky130_fd_sc_hd__inv_4 _2963_ (.A(net859),
    .Y(_2714_));
 sky130_fd_sc_hd__inv_2 _2964_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ),
    .Y(_2715_));
 sky130_fd_sc_hd__inv_2 _2965_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ),
    .Y(_2716_));
 sky130_fd_sc_hd__inv_2 _2966_ (.A(net509),
    .Y(_2717_));
 sky130_fd_sc_hd__inv_2 _2967_ (.A(net741),
    .Y(_2718_));
 sky130_fd_sc_hd__inv_2 _2968_ (.A(net155),
    .Y(net33));
 sky130_fd_sc_hd__inv_2 _2969_ (.A(\z80.tv80s.i_tv80_core.Halt_FF ),
    .Y(net22));
 sky130_fd_sc_hd__inv_2 _2970_ (.A(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .Y(_2719_));
 sky130_fd_sc_hd__inv_2 _2971_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ),
    .Y(_2720_));
 sky130_fd_sc_hd__inv_2 _2972_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ),
    .Y(_2721_));
 sky130_fd_sc_hd__inv_2 _2973_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .Y(_2722_));
 sky130_fd_sc_hd__inv_2 _2974_ (.A(net154),
    .Y(_2723_));
 sky130_fd_sc_hd__inv_2 _2975_ (.A(\z80.tv80s.i_tv80_core.BusA[1] ),
    .Y(_2724_));
 sky130_fd_sc_hd__inv_2 _2976_ (.A(\z80.tv80s.i_tv80_core.BusA[2] ),
    .Y(_2725_));
 sky130_fd_sc_hd__inv_2 _2977_ (.A(net652),
    .Y(_2726_));
 sky130_fd_sc_hd__inv_2 _2978_ (.A(net627),
    .Y(_2727_));
 sky130_fd_sc_hd__inv_2 _2979_ (.A(net590),
    .Y(_2728_));
 sky130_fd_sc_hd__inv_2 _2980_ (.A(net601),
    .Y(_2729_));
 sky130_fd_sc_hd__inv_2 _2981_ (.A(\z80.tv80s.i_tv80_core.F[4] ),
    .Y(_2730_));
 sky130_fd_sc_hd__inv_2 _2982_ (.A(\z80.tv80s.i_tv80_core.Arith16_r ),
    .Y(_2731_));
 sky130_fd_sc_hd__inv_2 _2983_ (.A(\z80.tv80s.di_reg[1] ),
    .Y(_2732_));
 sky130_fd_sc_hd__inv_2 _2984_ (.A(\z80.tv80s.di_reg[0] ),
    .Y(_2733_));
 sky130_fd_sc_hd__inv_2 _2985_ (.A(\z80.tv80s.di_reg[3] ),
    .Y(_2734_));
 sky130_fd_sc_hd__inv_2 _2986_ (.A(\z80.tv80s.di_reg[2] ),
    .Y(_2735_));
 sky130_fd_sc_hd__inv_2 _2987_ (.A(\z80.tv80s.di_reg[4] ),
    .Y(_2736_));
 sky130_fd_sc_hd__inv_2 _2988_ (.A(\z80.tv80s.di_reg[6] ),
    .Y(_2737_));
 sky130_fd_sc_hd__inv_2 _2989_ (.A(net816),
    .Y(_2738_));
 sky130_fd_sc_hd__inv_2 _2990_ (.A(net813),
    .Y(_2739_));
 sky130_fd_sc_hd__inv_2 _2991_ (.A(\z80.tv80s.i_tv80_core.PC[1] ),
    .Y(_2740_));
 sky130_fd_sc_hd__inv_2 _2992_ (.A(net609),
    .Y(_2741_));
 sky130_fd_sc_hd__inv_2 _2993_ (.A(net642),
    .Y(_2742_));
 sky130_fd_sc_hd__inv_2 _2994_ (.A(\z80.tv80s.i_tv80_core.PC[4] ),
    .Y(_2743_));
 sky130_fd_sc_hd__inv_2 _2995_ (.A(\z80.tv80s.i_tv80_core.PC[5] ),
    .Y(_2744_));
 sky130_fd_sc_hd__inv_2 _2996_ (.A(net631),
    .Y(_2745_));
 sky130_fd_sc_hd__inv_2 _2997_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .Y(_2746_));
 sky130_fd_sc_hd__inv_2 _2998_ (.A(\z80.tv80s.i_tv80_core.SP[8] ),
    .Y(_2747_));
 sky130_fd_sc_hd__inv_2 _2999_ (.A(net521),
    .Y(_2748_));
 sky130_fd_sc_hd__inv_2 _3000_ (.A(net9),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _3001_ (.A(net12),
    .Y(_0023_));
 sky130_fd_sc_hd__o31a_1 _3002_ (.A1(net167),
    .A2(net586),
    .A3(net309),
    .B1(net142),
    .X(_2749_));
 sky130_fd_sc_hd__nor2_1 _3003_ (.A(net123),
    .B(net120),
    .Y(_2750_));
 sky130_fd_sc_hd__or2_4 _3004_ (.A(net123),
    .B(net120),
    .X(_2751_));
 sky130_fd_sc_hd__and2_1 _3005_ (.A(\z80.tv80s.i_tv80_core.IR[7] ),
    .B(\z80.tv80s.i_tv80_core.IR[6] ),
    .X(_2752_));
 sky130_fd_sc_hd__nand2_8 _3006_ (.A(\z80.tv80s.i_tv80_core.IR[7] ),
    .B(\z80.tv80s.i_tv80_core.IR[6] ),
    .Y(_2753_));
 sky130_fd_sc_hd__or4bb_4 _3007_ (.A(net124),
    .B(net121),
    .C_N(\z80.tv80s.i_tv80_core.IR[7] ),
    .D_N(\z80.tv80s.i_tv80_core.IR[6] ),
    .X(_2754_));
 sky130_fd_sc_hd__and3_1 _3008_ (.A(net133),
    .B(net135),
    .C(_2700_),
    .X(_2755_));
 sky130_fd_sc_hd__nand3b_4 _3009_ (.A_N(net131),
    .B(net135),
    .C(net133),
    .Y(_2756_));
 sky130_fd_sc_hd__nor2_2 _3010_ (.A(net128),
    .B(_2756_),
    .Y(_2757_));
 sky130_fd_sc_hd__inv_2 _3011_ (.A(_2757_),
    .Y(_2758_));
 sky130_fd_sc_hd__nor2_1 _3012_ (.A(_2754_),
    .B(_2758_),
    .Y(_2759_));
 sky130_fd_sc_hd__nor2_1 _3013_ (.A(_2702_),
    .B(net122),
    .Y(_2760_));
 sky130_fd_sc_hd__nand2_1 _3014_ (.A(net123),
    .B(_2703_),
    .Y(_2761_));
 sky130_fd_sc_hd__nand2_2 _3015_ (.A(_2752_),
    .B(_2760_),
    .Y(_2762_));
 sky130_fd_sc_hd__nor2_1 _3016_ (.A(_2756_),
    .B(_2762_),
    .Y(_2763_));
 sky130_fd_sc_hd__or2_1 _3017_ (.A(_2756_),
    .B(_2762_),
    .X(_2764_));
 sky130_fd_sc_hd__nor2_1 _3018_ (.A(net118),
    .B(_2764_),
    .Y(_2765_));
 sky130_fd_sc_hd__or2_4 _3019_ (.A(\z80.tv80s.i_tv80_core.IR[7] ),
    .B(\z80.tv80s.i_tv80_core.IR[6] ),
    .X(_2766_));
 sky130_fd_sc_hd__or3_4 _3020_ (.A(net133),
    .B(net135),
    .C(net131),
    .X(_2767_));
 sky130_fd_sc_hd__nor4_4 _3021_ (.A(net128),
    .B(_2751_),
    .C(_2766_),
    .D(_2767_),
    .Y(_2768_));
 sky130_fd_sc_hd__nor2_2 _3022_ (.A(net126),
    .B(_2764_),
    .Y(_2769_));
 sky130_fd_sc_hd__or3_1 _3023_ (.A(_2759_),
    .B(_2763_),
    .C(_2768_),
    .X(_2770_));
 sky130_fd_sc_hd__or3b_4 _3024_ (.A(net134),
    .B(net132),
    .C_N(net135),
    .X(_2771_));
 sky130_fd_sc_hd__or2_2 _3025_ (.A(net127),
    .B(_2771_),
    .X(_2772_));
 sky130_fd_sc_hd__nor2_4 _3026_ (.A(_2766_),
    .B(_2772_),
    .Y(_2773_));
 sky130_fd_sc_hd__nor2_4 _3027_ (.A(_2698_),
    .B(net135),
    .Y(_2774_));
 sky130_fd_sc_hd__or3b_4 _3028_ (.A(net135),
    .B(net131),
    .C_N(net133),
    .X(_2775_));
 sky130_fd_sc_hd__or2_2 _3029_ (.A(net121),
    .B(_2766_),
    .X(_2776_));
 sky130_fd_sc_hd__nor2_2 _3030_ (.A(_2775_),
    .B(_2776_),
    .Y(_2777_));
 sky130_fd_sc_hd__or2_1 _3031_ (.A(_2775_),
    .B(_2776_),
    .X(_2778_));
 sky130_fd_sc_hd__or3b_4 _3032_ (.A(\z80.tv80s.i_tv80_core.IR[7] ),
    .B(\z80.tv80s.i_tv80_core.IR[6] ),
    .C_N(net121),
    .X(_2779_));
 sky130_fd_sc_hd__or2_1 _3033_ (.A(_2702_),
    .B(_2779_),
    .X(_2780_));
 sky130_fd_sc_hd__nor2_2 _3034_ (.A(_2775_),
    .B(_2780_),
    .Y(_2781_));
 sky130_fd_sc_hd__or2_1 _3035_ (.A(_2775_),
    .B(_2780_),
    .X(_2782_));
 sky130_fd_sc_hd__a211o_1 _3036_ (.A1(net121),
    .A2(_2773_),
    .B1(_2777_),
    .C1(_2781_),
    .X(_2783_));
 sky130_fd_sc_hd__or4b_2 _3037_ (.A(net121),
    .B(\z80.tv80s.i_tv80_core.IR[7] ),
    .C(\z80.tv80s.i_tv80_core.IR[6] ),
    .D_N(net124),
    .X(_2784_));
 sky130_fd_sc_hd__nor2_2 _3038_ (.A(_2767_),
    .B(_2784_),
    .Y(_2785_));
 sky130_fd_sc_hd__nor2_1 _3039_ (.A(net127),
    .B(net123),
    .Y(_2786_));
 sky130_fd_sc_hd__or2_2 _3040_ (.A(net127),
    .B(net123),
    .X(_2787_));
 sky130_fd_sc_hd__a211oi_1 _3041_ (.A1(_2756_),
    .A2(_2767_),
    .B1(_2779_),
    .C1(_2787_),
    .Y(_2788_));
 sky130_fd_sc_hd__nor2_4 _3042_ (.A(net127),
    .B(_2702_),
    .Y(_2789_));
 sky130_fd_sc_hd__nand2_4 _3043_ (.A(net119),
    .B(net124),
    .Y(_2790_));
 sky130_fd_sc_hd__nor2_1 _3044_ (.A(_2767_),
    .B(_2779_),
    .Y(_2791_));
 sky130_fd_sc_hd__or2_1 _3045_ (.A(_2767_),
    .B(_2779_),
    .X(_2792_));
 sky130_fd_sc_hd__nor2_1 _3046_ (.A(_2753_),
    .B(_2767_),
    .Y(_2793_));
 sky130_fd_sc_hd__and2_1 _3047_ (.A(_2751_),
    .B(_2793_),
    .X(_2794_));
 sky130_fd_sc_hd__a2111o_1 _3048_ (.A1(_2789_),
    .A2(_2791_),
    .B1(_2794_),
    .C1(_2788_),
    .D1(_2785_),
    .X(_2795_));
 sky130_fd_sc_hd__nand2_1 _3049_ (.A(_2698_),
    .B(net131),
    .Y(_2796_));
 sky130_fd_sc_hd__and3b_1 _3050_ (.A_N(net133),
    .B(net131),
    .C(net130),
    .X(_2797_));
 sky130_fd_sc_hd__and3_1 _3051_ (.A(\z80.tv80s.i_tv80_core.IR[0] ),
    .B(\z80.tv80s.i_tv80_core.IR[7] ),
    .C(\z80.tv80s.i_tv80_core.IR[6] ),
    .X(_2798_));
 sky130_fd_sc_hd__and3_2 _3052_ (.A(_2750_),
    .B(_2797_),
    .C(_2798_),
    .X(_2799_));
 sky130_fd_sc_hd__nor2_1 _3053_ (.A(net118),
    .B(_2771_),
    .Y(_2800_));
 sky130_fd_sc_hd__or4bb_4 _3054_ (.A(net133),
    .B(net131),
    .C_N(net128),
    .D_N(net135),
    .X(_2801_));
 sky130_fd_sc_hd__a21oi_1 _3055_ (.A1(_2767_),
    .A2(_2801_),
    .B1(_2754_),
    .Y(_2802_));
 sky130_fd_sc_hd__or2_1 _3056_ (.A(_2799_),
    .B(_2802_),
    .X(_2803_));
 sky130_fd_sc_hd__or4_1 _3057_ (.A(_2770_),
    .B(_2783_),
    .C(_2795_),
    .D(_2803_),
    .X(_2804_));
 sky130_fd_sc_hd__nor2_4 _3058_ (.A(_2702_),
    .B(_2703_),
    .Y(_2805_));
 sky130_fd_sc_hd__nand2_2 _3059_ (.A(net125),
    .B(net122),
    .Y(_2806_));
 sky130_fd_sc_hd__nor2_1 _3060_ (.A(_2753_),
    .B(_2806_),
    .Y(_2807_));
 sky130_fd_sc_hd__or2_2 _3061_ (.A(_2753_),
    .B(_2806_),
    .X(_2808_));
 sky130_fd_sc_hd__nor2_1 _3062_ (.A(_2756_),
    .B(_2808_),
    .Y(_2809_));
 sky130_fd_sc_hd__and3_1 _3063_ (.A(net133),
    .B(net135),
    .C(net131),
    .X(_2810_));
 sky130_fd_sc_hd__or3_4 _3064_ (.A(_2698_),
    .B(_2699_),
    .C(_2700_),
    .X(_2811_));
 sky130_fd_sc_hd__nor2_4 _3065_ (.A(_2779_),
    .B(_2811_),
    .Y(_2812_));
 sky130_fd_sc_hd__nor3_2 _3066_ (.A(net118),
    .B(_2754_),
    .C(_2756_),
    .Y(_2813_));
 sky130_fd_sc_hd__nor2_2 _3067_ (.A(_2801_),
    .B(_2808_),
    .Y(_2814_));
 sky130_fd_sc_hd__or2_2 _3068_ (.A(_2813_),
    .B(_2814_),
    .X(_2815_));
 sky130_fd_sc_hd__or3_1 _3069_ (.A(_2809_),
    .B(_2812_),
    .C(_2815_),
    .X(_2816_));
 sky130_fd_sc_hd__nor2_1 _3070_ (.A(_2776_),
    .B(_2811_),
    .Y(_2817_));
 sky130_fd_sc_hd__nor2_2 _3071_ (.A(net125),
    .B(_2703_),
    .Y(_2818_));
 sky130_fd_sc_hd__nand2b_2 _3072_ (.A_N(net125),
    .B(net122),
    .Y(_2819_));
 sky130_fd_sc_hd__nor2_2 _3073_ (.A(_2753_),
    .B(_2819_),
    .Y(_2820_));
 sky130_fd_sc_hd__nor2_1 _3074_ (.A(net119),
    .B(_2811_),
    .Y(_2821_));
 sky130_fd_sc_hd__and2_1 _3075_ (.A(_2800_),
    .B(_2820_),
    .X(_2822_));
 sky130_fd_sc_hd__a221o_1 _3076_ (.A1(_2807_),
    .A2(_2810_),
    .B1(_2820_),
    .B2(_2821_),
    .C1(_2822_),
    .X(_2823_));
 sky130_fd_sc_hd__a31o_1 _3077_ (.A1(_2756_),
    .A2(_2796_),
    .A3(_2801_),
    .B1(_2776_),
    .X(_2824_));
 sky130_fd_sc_hd__or2_1 _3078_ (.A(net124),
    .B(_2779_),
    .X(_2825_));
 sky130_fd_sc_hd__a22o_1 _3079_ (.A1(_2700_),
    .A2(net118),
    .B1(_2756_),
    .B2(net133),
    .X(_2826_));
 sky130_fd_sc_hd__o21ai_1 _3080_ (.A1(_2825_),
    .A2(_2826_),
    .B1(_2824_),
    .Y(_2827_));
 sky130_fd_sc_hd__and3_2 _3081_ (.A(_2751_),
    .B(_2797_),
    .C(_2798_),
    .X(_2828_));
 sky130_fd_sc_hd__nor2_1 _3082_ (.A(_2753_),
    .B(_2811_),
    .Y(_2829_));
 sky130_fd_sc_hd__nand2_1 _3083_ (.A(net121),
    .B(_2787_),
    .Y(_2830_));
 sky130_fd_sc_hd__a31o_1 _3084_ (.A1(_2752_),
    .A2(_2810_),
    .A3(_2830_),
    .B1(_2828_),
    .X(_2831_));
 sky130_fd_sc_hd__or4_1 _3085_ (.A(_2817_),
    .B(_2823_),
    .C(_2827_),
    .D(_2831_),
    .X(_2832_));
 sky130_fd_sc_hd__or3_2 _3086_ (.A(_2804_),
    .B(_2816_),
    .C(_2832_),
    .X(_2833_));
 sky130_fd_sc_hd__nor2_4 _3087_ (.A(_2704_),
    .B(\z80.tv80s.i_tv80_core.IR[6] ),
    .Y(_2834_));
 sky130_fd_sc_hd__or2_4 _3088_ (.A(_2704_),
    .B(\z80.tv80s.i_tv80_core.IR[6] ),
    .X(_2835_));
 sky130_fd_sc_hd__nand3b_4 _3089_ (.A_N(\z80.tv80s.i_tv80_core.IR[6] ),
    .B(\z80.tv80s.i_tv80_core.IR[7] ),
    .C(net120),
    .Y(_2836_));
 sky130_fd_sc_hd__nor2_1 _3090_ (.A(_2767_),
    .B(_2836_),
    .Y(_2837_));
 sky130_fd_sc_hd__or2_2 _3091_ (.A(_2767_),
    .B(_2836_),
    .X(_2838_));
 sky130_fd_sc_hd__or2_2 _3092_ (.A(_2771_),
    .B(_2836_),
    .X(_2839_));
 sky130_fd_sc_hd__or3_4 _3093_ (.A(net134),
    .B(net132),
    .C(_2836_),
    .X(_2840_));
 sky130_fd_sc_hd__or2_2 _3094_ (.A(_2756_),
    .B(_2836_),
    .X(_2841_));
 sky130_fd_sc_hd__or2_2 _3095_ (.A(_2775_),
    .B(_2836_),
    .X(_2842_));
 sky130_fd_sc_hd__or3_4 _3096_ (.A(_2698_),
    .B(net132),
    .C(_2836_),
    .X(_2843_));
 sky130_fd_sc_hd__nand2_2 _3097_ (.A(_2841_),
    .B(_2842_),
    .Y(_2844_));
 sky130_fd_sc_hd__nor2_2 _3098_ (.A(net131),
    .B(_2836_),
    .Y(_2845_));
 sky130_fd_sc_hd__nand2_2 _3099_ (.A(net132),
    .B(net119),
    .Y(_2846_));
 sky130_fd_sc_hd__inv_2 _3100_ (.A(_2846_),
    .Y(_2847_));
 sky130_fd_sc_hd__nor2_1 _3101_ (.A(_2774_),
    .B(_2846_),
    .Y(_2848_));
 sky130_fd_sc_hd__or4_1 _3102_ (.A(_2702_),
    .B(_2774_),
    .C(_2836_),
    .D(_2846_),
    .X(_2849_));
 sky130_fd_sc_hd__or4_1 _3103_ (.A(net118),
    .B(net124),
    .C(_2811_),
    .D(_2836_),
    .X(_2850_));
 sky130_fd_sc_hd__and2_1 _3104_ (.A(_2704_),
    .B(\z80.tv80s.i_tv80_core.IR[6] ),
    .X(_2851_));
 sky130_fd_sc_hd__nand2_4 _3105_ (.A(_2704_),
    .B(\z80.tv80s.i_tv80_core.IR[6] ),
    .Y(_2852_));
 sky130_fd_sc_hd__or4_4 _3106_ (.A(_2698_),
    .B(_2699_),
    .C(_2700_),
    .D(net95),
    .X(_2853_));
 sky130_fd_sc_hd__nor2_1 _3107_ (.A(net120),
    .B(_2853_),
    .Y(_2854_));
 sky130_fd_sc_hd__or2_1 _3108_ (.A(net122),
    .B(_2853_),
    .X(_2855_));
 sky130_fd_sc_hd__nor2_2 _3109_ (.A(_2775_),
    .B(net95),
    .Y(_2856_));
 sky130_fd_sc_hd__or2_4 _3110_ (.A(_2775_),
    .B(net95),
    .X(_2857_));
 sky130_fd_sc_hd__a32o_1 _3111_ (.A1(net127),
    .A2(net120),
    .A3(_2856_),
    .B1(_2854_),
    .B2(net123),
    .X(_2858_));
 sky130_fd_sc_hd__and3_2 _3112_ (.A(net134),
    .B(_2699_),
    .C(net132),
    .X(_2859_));
 sky130_fd_sc_hd__nand2_8 _3113_ (.A(net131),
    .B(_2774_),
    .Y(_2860_));
 sky130_fd_sc_hd__and3_2 _3114_ (.A(net127),
    .B(net123),
    .C(net121),
    .X(_2861_));
 sky130_fd_sc_hd__nand3_1 _3115_ (.A(net127),
    .B(net123),
    .C(net120),
    .Y(_2862_));
 sky130_fd_sc_hd__nor2_1 _3116_ (.A(_2811_),
    .B(_2862_),
    .Y(_2863_));
 sky130_fd_sc_hd__a221o_1 _3117_ (.A1(net120),
    .A2(_2797_),
    .B1(_2860_),
    .B2(_2750_),
    .C1(_2863_),
    .X(_2864_));
 sky130_fd_sc_hd__or3_4 _3118_ (.A(net133),
    .B(net135),
    .C(_2700_),
    .X(_2865_));
 sky130_fd_sc_hd__o311a_1 _3119_ (.A1(net133),
    .A2(_2699_),
    .A3(net128),
    .B1(_2775_),
    .C1(_2865_),
    .X(_2866_));
 sky130_fd_sc_hd__nor2_1 _3120_ (.A(_2753_),
    .B(_2866_),
    .Y(_2867_));
 sky130_fd_sc_hd__and3_1 _3121_ (.A(net146),
    .B(_2852_),
    .C(net94),
    .X(_2868_));
 sky130_fd_sc_hd__nor2_1 _3122_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ),
    .B(net151),
    .Y(_2869_));
 sky130_fd_sc_hd__o211a_1 _3123_ (.A1(net133),
    .A2(_2846_),
    .B1(_2865_),
    .C1(_2775_),
    .X(_2870_));
 sky130_fd_sc_hd__a21oi_1 _3124_ (.A1(_2754_),
    .A2(_2808_),
    .B1(_2866_),
    .Y(_2871_));
 sky130_fd_sc_hd__or4_1 _3125_ (.A(net128),
    .B(net124),
    .C(_2836_),
    .D(_2865_),
    .X(_2872_));
 sky130_fd_sc_hd__a211o_1 _3126_ (.A1(_2700_),
    .A2(net128),
    .B1(_2757_),
    .C1(_2848_),
    .X(_2873_));
 sky130_fd_sc_hd__and4_1 _3127_ (.A(\z80.tv80s.i_tv80_core.IR[0] ),
    .B(_2818_),
    .C(_2834_),
    .D(_2847_),
    .X(_2874_));
 sky130_fd_sc_hd__a211o_1 _3128_ (.A1(net133),
    .A2(net135),
    .B1(net131),
    .C1(net127),
    .X(_2875_));
 sky130_fd_sc_hd__o31a_1 _3129_ (.A1(_2700_),
    .A2(net118),
    .A3(_2774_),
    .B1(_2875_),
    .X(_2876_));
 sky130_fd_sc_hd__a21oi_1 _3130_ (.A1(_2758_),
    .A2(_2826_),
    .B1(_2780_),
    .Y(_2877_));
 sky130_fd_sc_hd__nor2_2 _3131_ (.A(_2775_),
    .B(_2825_),
    .Y(_2878_));
 sky130_fd_sc_hd__and2_1 _3132_ (.A(_2703_),
    .B(_2773_),
    .X(_2879_));
 sky130_fd_sc_hd__or2_1 _3133_ (.A(_2878_),
    .B(_2879_),
    .X(_2880_));
 sky130_fd_sc_hd__and3_4 _3134_ (.A(net128),
    .B(_2755_),
    .C(_2820_),
    .X(_2881_));
 sky130_fd_sc_hd__nor4_1 _3135_ (.A(net118),
    .B(_2751_),
    .C(_2766_),
    .D(_2767_),
    .Y(_2882_));
 sky130_fd_sc_hd__or2_1 _3136_ (.A(_2881_),
    .B(_2882_),
    .X(_2883_));
 sky130_fd_sc_hd__nor2_1 _3137_ (.A(_2762_),
    .B(_2801_),
    .Y(_2884_));
 sky130_fd_sc_hd__and2_4 _3138_ (.A(_2757_),
    .B(_2820_),
    .X(_2885_));
 sky130_fd_sc_hd__or2_1 _3139_ (.A(_2884_),
    .B(_2885_),
    .X(_2886_));
 sky130_fd_sc_hd__or4_1 _3140_ (.A(_2877_),
    .B(_2880_),
    .C(_2883_),
    .D(_2886_),
    .X(_2887_));
 sky130_fd_sc_hd__a31o_1 _3141_ (.A1(_2699_),
    .A2(net127),
    .A3(net120),
    .B1(net131),
    .X(_2888_));
 sky130_fd_sc_hd__o211ai_1 _3142_ (.A1(_2699_),
    .A2(net123),
    .B1(_2888_),
    .C1(net134),
    .Y(_2889_));
 sky130_fd_sc_hd__nor2_2 _3143_ (.A(_2771_),
    .B(net95),
    .Y(_2890_));
 sky130_fd_sc_hd__nor2_8 _3144_ (.A(_2703_),
    .B(_2790_),
    .Y(_2891_));
 sky130_fd_sc_hd__nand3b_4 _3145_ (.A_N(net127),
    .B(net123),
    .C(net120),
    .Y(_2892_));
 sky130_fd_sc_hd__nor2_1 _3146_ (.A(_2853_),
    .B(_2892_),
    .Y(_2893_));
 sky130_fd_sc_hd__a32o_1 _3147_ (.A1(_2805_),
    .A2(_2821_),
    .A3(net96),
    .B1(_2890_),
    .B2(_2750_),
    .X(_2894_));
 sky130_fd_sc_hd__or4_4 _3148_ (.A(net133),
    .B(_2699_),
    .C(_2700_),
    .D(net95),
    .X(_2895_));
 sky130_fd_sc_hd__nor2_1 _3149_ (.A(_2756_),
    .B(net95),
    .Y(_2896_));
 sky130_fd_sc_hd__nand2_2 _3150_ (.A(_2755_),
    .B(net96),
    .Y(_2897_));
 sky130_fd_sc_hd__o211a_1 _3151_ (.A1(_2751_),
    .A2(_2771_),
    .B1(net96),
    .C1(_2889_),
    .X(_2898_));
 sky130_fd_sc_hd__a31o_1 _3152_ (.A1(_2760_),
    .A2(_2834_),
    .A3(_2873_),
    .B1(_2871_),
    .X(_2899_));
 sky130_fd_sc_hd__o32a_1 _3153_ (.A1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ),
    .A2(net151),
    .A3(_2868_),
    .B1(_2870_),
    .B2(_2762_),
    .X(_2900_));
 sky130_fd_sc_hd__or4b_1 _3154_ (.A(_2874_),
    .B(_2893_),
    .C(_2898_),
    .D_N(_2900_),
    .X(_2901_));
 sky130_fd_sc_hd__o32a_1 _3155_ (.A1(_2761_),
    .A2(_2835_),
    .A3(_2876_),
    .B1(_2762_),
    .B2(_2772_),
    .X(_2902_));
 sky130_fd_sc_hd__o311a_1 _3156_ (.A1(_2751_),
    .A2(_2801_),
    .A3(_2835_),
    .B1(_2872_),
    .C1(_2902_),
    .X(_2903_));
 sky130_fd_sc_hd__and4b_1 _3157_ (.A_N(_2845_),
    .B(_2849_),
    .C(_2850_),
    .D(_2903_),
    .X(_2904_));
 sky130_fd_sc_hd__or4b_1 _3158_ (.A(_2894_),
    .B(_2899_),
    .C(_2901_),
    .D_N(_2904_),
    .X(_2905_));
 sky130_fd_sc_hd__a21o_1 _3159_ (.A1(_2834_),
    .A2(_2864_),
    .B1(_2858_),
    .X(_2906_));
 sky130_fd_sc_hd__a2111o_1 _3160_ (.A1(_2818_),
    .A2(_2867_),
    .B1(_2887_),
    .C1(_2905_),
    .D1(_2906_),
    .X(_2907_));
 sky130_fd_sc_hd__o21ai_4 _3161_ (.A1(_2833_),
    .A2(_2907_),
    .B1(net163),
    .Y(_2908_));
 sky130_fd_sc_hd__nor2_1 _3162_ (.A(net94),
    .B(_2891_),
    .Y(_2909_));
 sky130_fd_sc_hd__a21o_1 _3163_ (.A1(net94),
    .A2(_2891_),
    .B1(net116),
    .X(_2910_));
 sky130_fd_sc_hd__o31ai_1 _3164_ (.A1(net95),
    .A2(_2909_),
    .A3(_2910_),
    .B1(net165),
    .Y(_2911_));
 sky130_fd_sc_hd__or2_1 _3165_ (.A(_2822_),
    .B(_2828_),
    .X(_2912_));
 sky130_fd_sc_hd__nor2_1 _3166_ (.A(_2753_),
    .B(_2775_),
    .Y(_2913_));
 sky130_fd_sc_hd__or2_2 _3167_ (.A(_2759_),
    .B(_2913_),
    .X(_2914_));
 sky130_fd_sc_hd__or4_1 _3168_ (.A(_2883_),
    .B(_2884_),
    .C(_2912_),
    .D(_2914_),
    .X(_2915_));
 sky130_fd_sc_hd__nor2_1 _3169_ (.A(_2753_),
    .B(_2860_),
    .Y(_2916_));
 sky130_fd_sc_hd__nor2_2 _3170_ (.A(_2756_),
    .B(_2766_),
    .Y(_2917_));
 sky130_fd_sc_hd__or2_1 _3171_ (.A(_2756_),
    .B(_2766_),
    .X(_2918_));
 sky130_fd_sc_hd__or2_1 _3172_ (.A(_2785_),
    .B(_2791_),
    .X(_2919_));
 sky130_fd_sc_hd__nor2_4 _3173_ (.A(_2766_),
    .B(_2801_),
    .Y(_2920_));
 sky130_fd_sc_hd__or2_1 _3174_ (.A(_2766_),
    .B(_2801_),
    .X(_2921_));
 sky130_fd_sc_hd__or3_1 _3175_ (.A(_2773_),
    .B(_2919_),
    .C(_2920_),
    .X(_2922_));
 sky130_fd_sc_hd__or4_1 _3176_ (.A(_2817_),
    .B(_2916_),
    .C(_2917_),
    .D(_2922_),
    .X(_2923_));
 sky130_fd_sc_hd__nor3_1 _3177_ (.A(_2816_),
    .B(_2915_),
    .C(_2923_),
    .Y(_2924_));
 sky130_fd_sc_hd__and3_2 _3178_ (.A(_2698_),
    .B(_2798_),
    .C(_2847_),
    .X(_2925_));
 sky130_fd_sc_hd__o2111a_2 _3179_ (.A1(net133),
    .A2(net118),
    .B1(_2752_),
    .C1(net135),
    .D1(net131),
    .X(_2926_));
 sky130_fd_sc_hd__nor2_2 _3180_ (.A(_2753_),
    .B(_2772_),
    .Y(_2927_));
 sky130_fd_sc_hd__or3_2 _3181_ (.A(net126),
    .B(_2753_),
    .C(_2771_),
    .X(_2928_));
 sky130_fd_sc_hd__nor2_1 _3182_ (.A(_2754_),
    .B(_2801_),
    .Y(_2929_));
 sky130_fd_sc_hd__o22a_1 _3183_ (.A1(_2753_),
    .A2(_2767_),
    .B1(_2801_),
    .B2(_2754_),
    .X(_2930_));
 sky130_fd_sc_hd__or2_1 _3184_ (.A(_2793_),
    .B(_2929_),
    .X(_2931_));
 sky130_fd_sc_hd__and3b_1 _3185_ (.A_N(_2926_),
    .B(_2928_),
    .C(_2930_),
    .X(_2932_));
 sky130_fd_sc_hd__nor2_2 _3186_ (.A(_2766_),
    .B(_2796_),
    .Y(_2933_));
 sky130_fd_sc_hd__or2_2 _3187_ (.A(_2766_),
    .B(_2796_),
    .X(_2934_));
 sky130_fd_sc_hd__nor2_2 _3188_ (.A(net145),
    .B(net147),
    .Y(_2935_));
 sky130_fd_sc_hd__or2_4 _3189_ (.A(net145),
    .B(net147),
    .X(_2936_));
 sky130_fd_sc_hd__a21oi_1 _3190_ (.A1(_2891_),
    .A2(_2936_),
    .B1(_2934_),
    .Y(_2937_));
 sky130_fd_sc_hd__a21oi_1 _3191_ (.A1(net149),
    .A2(net94),
    .B1(_2835_),
    .Y(_2938_));
 sky130_fd_sc_hd__nor2_4 _3192_ (.A(_2766_),
    .B(_2860_),
    .Y(_2939_));
 sky130_fd_sc_hd__and3_2 _3193_ (.A(net121),
    .B(net146),
    .C(_2789_),
    .X(_2940_));
 sky130_fd_sc_hd__nor2_2 _3194_ (.A(_2753_),
    .B(_2865_),
    .Y(_2941_));
 sky130_fd_sc_hd__or2_2 _3195_ (.A(_2753_),
    .B(_2865_),
    .X(_2942_));
 sky130_fd_sc_hd__or2_2 _3196_ (.A(_2799_),
    .B(_2941_),
    .X(_2943_));
 sky130_fd_sc_hd__nor3_1 _3197_ (.A(net97),
    .B(_2937_),
    .C(_2943_),
    .Y(_2944_));
 sky130_fd_sc_hd__nor2_1 _3198_ (.A(_2885_),
    .B(_2938_),
    .Y(_2945_));
 sky130_fd_sc_hd__o311a_1 _3199_ (.A1(_2766_),
    .A2(_2860_),
    .A3(_2940_),
    .B1(_2945_),
    .C1(net95),
    .X(_0370_));
 sky130_fd_sc_hd__and3_1 _3200_ (.A(_2932_),
    .B(_2944_),
    .C(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__o221a_1 _3201_ (.A1(net150),
    .A2(_2778_),
    .B1(_2779_),
    .B2(_2775_),
    .C1(_2764_),
    .X(_0372_));
 sky130_fd_sc_hd__a31o_1 _3202_ (.A1(_2924_),
    .A2(_0371_),
    .A3(_0372_),
    .B1(_2911_),
    .X(_0373_));
 sky130_fd_sc_hd__or4_4 _3203_ (.A(_2698_),
    .B(net135),
    .C(_2780_),
    .D(_2846_),
    .X(_0374_));
 sky130_fd_sc_hd__nand2b_1 _3204_ (.A_N(_2813_),
    .B(_0374_),
    .Y(_0375_));
 sky130_fd_sc_hd__nand2_1 _3205_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ),
    .B(_0375_),
    .Y(_0376_));
 sky130_fd_sc_hd__nor2_4 _3206_ (.A(net164),
    .B(net163),
    .Y(_0377_));
 sky130_fd_sc_hd__or2_1 _3207_ (.A(net164),
    .B(net163),
    .X(_0378_));
 sky130_fd_sc_hd__nor2_4 _3208_ (.A(_2819_),
    .B(_2853_),
    .Y(_0379_));
 sky130_fd_sc_hd__nor2_1 _3209_ (.A(_2845_),
    .B(_0379_),
    .Y(_0380_));
 sky130_fd_sc_hd__or3_2 _3210_ (.A(net133),
    .B(net131),
    .C(net95),
    .X(_0381_));
 sky130_fd_sc_hd__nand4_2 _3211_ (.A(_2895_),
    .B(_2897_),
    .C(_0380_),
    .D(_0381_),
    .Y(_0382_));
 sky130_fd_sc_hd__o221a_1 _3212_ (.A1(_2843_),
    .A2(_2936_),
    .B1(_0381_),
    .B2(net147),
    .C1(_2895_),
    .X(_0383_));
 sky130_fd_sc_hd__nor2_4 _3213_ (.A(net145),
    .B(net143),
    .Y(_0384_));
 sky130_fd_sc_hd__or2_4 _3214_ (.A(net145),
    .B(net143),
    .X(_0385_));
 sky130_fd_sc_hd__nand2_1 _3215_ (.A(_0379_),
    .B(_0384_),
    .Y(_0386_));
 sky130_fd_sc_hd__o221a_1 _3216_ (.A1(net147),
    .A2(_2839_),
    .B1(_2936_),
    .B2(_2838_),
    .C1(_2897_),
    .X(_0387_));
 sky130_fd_sc_hd__a41o_1 _3217_ (.A1(_0382_),
    .A2(_0383_),
    .A3(_0386_),
    .A4(_0387_),
    .B1(net105),
    .X(_0388_));
 sky130_fd_sc_hd__nand4_4 _3218_ (.A(_2908_),
    .B(_0373_),
    .C(_0376_),
    .D(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__and2b_1 _3219_ (.A_N(_2749_),
    .B(_0389_),
    .X(_0390_));
 sky130_fd_sc_hd__o21a_1 _3220_ (.A1(net146),
    .A2(_2764_),
    .B1(_2924_),
    .X(_0391_));
 sky130_fd_sc_hd__o21a_2 _3221_ (.A1(net143),
    .A2(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .B1(net117),
    .X(_0392_));
 sky130_fd_sc_hd__o21ai_4 _3222_ (.A1(net143),
    .A2(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .B1(net117),
    .Y(_0393_));
 sky130_fd_sc_hd__o32a_1 _3223_ (.A1(net150),
    .A2(_2751_),
    .A3(_2766_),
    .B1(_2825_),
    .B2(_0392_),
    .X(_0394_));
 sky130_fd_sc_hd__a21o_1 _3224_ (.A1(_2784_),
    .A2(_0394_),
    .B1(_2775_),
    .X(_0395_));
 sky130_fd_sc_hd__and2_4 _3225_ (.A(net117),
    .B(net143),
    .X(_0396_));
 sky130_fd_sc_hd__nand2_1 _3226_ (.A(net117),
    .B(net144),
    .Y(_0397_));
 sky130_fd_sc_hd__nor2_1 _3227_ (.A(net128),
    .B(_2782_),
    .Y(_0398_));
 sky130_fd_sc_hd__nand2_1 _3228_ (.A(_0397_),
    .B(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__o311a_1 _3229_ (.A1(net118),
    .A2(net144),
    .A3(_2782_),
    .B1(_0395_),
    .C1(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__a31o_1 _3230_ (.A1(_0371_),
    .A2(_0391_),
    .A3(_0400_),
    .B1(_2911_),
    .X(_0401_));
 sky130_fd_sc_hd__o21a_1 _3231_ (.A1(_2897_),
    .A2(_0392_),
    .B1(_0386_),
    .X(_0402_));
 sky130_fd_sc_hd__or2_1 _3232_ (.A(net147),
    .B(_2840_),
    .X(_0403_));
 sky130_fd_sc_hd__a41o_1 _3233_ (.A1(_0382_),
    .A2(_0383_),
    .A3(_0402_),
    .A4(_0403_),
    .B1(net105),
    .X(_0404_));
 sky130_fd_sc_hd__and4_2 _3234_ (.A(_2908_),
    .B(_0376_),
    .C(_0401_),
    .D(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__or2_2 _3235_ (.A(_2749_),
    .B(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__mux2_2 _3236_ (.A0(\z80.tv80s.i_tv80_core.F[6] ),
    .A1(\z80.tv80s.i_tv80_core.F[0] ),
    .S(net124),
    .X(_0407_));
 sky130_fd_sc_hd__xnor2_4 _3237_ (.A(net119),
    .B(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__nor2_1 _3238_ (.A(_2703_),
    .B(_2787_),
    .Y(_0409_));
 sky130_fd_sc_hd__or3b_1 _3239_ (.A(net127),
    .B(net123),
    .C_N(net120),
    .X(_0410_));
 sky130_fd_sc_hd__and3_2 _3240_ (.A(net127),
    .B(_2702_),
    .C(net120),
    .X(_0411_));
 sky130_fd_sc_hd__and4b_1 _3241_ (.A_N(net123),
    .B(net120),
    .C(\z80.tv80s.i_tv80_core.F[2] ),
    .D(net127),
    .X(_0412_));
 sky130_fd_sc_hd__o21ba_1 _3242_ (.A1(\z80.tv80s.i_tv80_core.F[2] ),
    .A2(_0410_),
    .B1_N(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _3243_ (.A0(_2892_),
    .A1(_2862_),
    .S(\z80.tv80s.i_tv80_core.F[7] ),
    .X(_0414_));
 sky130_fd_sc_hd__o211a_2 _3244_ (.A1(net120),
    .A2(_0408_),
    .B1(_0413_),
    .C1(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__o2111a_2 _3245_ (.A1(net120),
    .A2(_0408_),
    .B1(_0413_),
    .C1(_0414_),
    .D1(net144),
    .X(_0416_));
 sky130_fd_sc_hd__or2_1 _3246_ (.A(_0393_),
    .B(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__nand2_1 _3247_ (.A(net150),
    .B(_0415_),
    .Y(_0418_));
 sky130_fd_sc_hd__and3_2 _3248_ (.A(_2706_),
    .B(_2757_),
    .C(_2820_),
    .X(_0419_));
 sky130_fd_sc_hd__nor2_1 _3249_ (.A(_2775_),
    .B(_2779_),
    .Y(_0420_));
 sky130_fd_sc_hd__or4_1 _3250_ (.A(net115),
    .B(_2834_),
    .C(net96),
    .D(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__a2111o_1 _3251_ (.A1(net116),
    .A2(_2777_),
    .B1(_2933_),
    .C1(_2939_),
    .D1(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__or2_4 _3252_ (.A(\z80.tv80s.i_tv80_core.IntCycle ),
    .B(net519),
    .X(_0423_));
 sky130_fd_sc_hd__inv_2 _3253_ (.A(_0423_),
    .Y(_0424_));
 sky130_fd_sc_hd__nand2_1 _3254_ (.A(_2936_),
    .B(_0423_),
    .Y(_0425_));
 sky130_fd_sc_hd__a221o_1 _3255_ (.A1(_2799_),
    .A2(_0393_),
    .B1(_0425_),
    .B2(net97),
    .C1(_0422_),
    .X(_0426_));
 sky130_fd_sc_hd__a32o_1 _3256_ (.A1(net149),
    .A2(_2793_),
    .A3(_0415_),
    .B1(_0417_),
    .B2(_2941_),
    .X(_0427_));
 sky130_fd_sc_hd__a311o_1 _3257_ (.A1(_2712_),
    .A2(_0384_),
    .A3(_0419_),
    .B1(_0426_),
    .C1(_0427_),
    .X(_0428_));
 sky130_fd_sc_hd__o21ba_1 _3258_ (.A1(_2932_),
    .A2(_2936_),
    .B1_N(_0428_),
    .X(_0429_));
 sky130_fd_sc_hd__nor2_4 _3259_ (.A(net117),
    .B(net147),
    .Y(_0430_));
 sky130_fd_sc_hd__nand2_4 _3260_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ),
    .B(net116),
    .Y(_0431_));
 sky130_fd_sc_hd__a21o_1 _3261_ (.A1(_2841_),
    .A2(_2895_),
    .B1(_0430_),
    .X(_0432_));
 sky130_fd_sc_hd__a22o_1 _3262_ (.A1(net147),
    .A2(_2841_),
    .B1(_2842_),
    .B2(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__a21oi_1 _3263_ (.A1(_2839_),
    .A2(_0430_),
    .B1(_2840_),
    .Y(_0434_));
 sky130_fd_sc_hd__or2_2 _3264_ (.A(_0379_),
    .B(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__and4b_1 _3265_ (.A_N(_0435_),
    .B(_0433_),
    .C(_2897_),
    .D(net115),
    .X(_0436_));
 sky130_fd_sc_hd__o21a_1 _3266_ (.A1(net147),
    .A2(_0381_),
    .B1(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__a22oi_2 _3267_ (.A1(_0391_),
    .A2(_0429_),
    .B1(_0437_),
    .B2(_0382_),
    .Y(_0438_));
 sky130_fd_sc_hd__nor3_2 _3268_ (.A(net163),
    .B(_2749_),
    .C(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__inv_2 _3269_ (.A(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__and3b_2 _3270_ (.A_N(_0390_),
    .B(_0406_),
    .C(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__a21o_1 _3271_ (.A1(net148),
    .A2(_0375_),
    .B1(net58),
    .X(_0442_));
 sky130_fd_sc_hd__nor2_2 _3272_ (.A(net576),
    .B(net507),
    .Y(_0443_));
 sky130_fd_sc_hd__or2_4 _3273_ (.A(\z80.tv80s.i_tv80_core.XY_State[1] ),
    .B(\z80.tv80s.i_tv80_core.XY_State[0] ),
    .X(_0444_));
 sky130_fd_sc_hd__nor2_2 _3274_ (.A(\z80.tv80s.i_tv80_core.XY_Ind ),
    .B(_0443_),
    .Y(_0445_));
 sky130_fd_sc_hd__nand2_8 _3275_ (.A(_0442_),
    .B(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__or4_1 _3276_ (.A(_2777_),
    .B(_2781_),
    .C(net96),
    .D(_2939_),
    .X(_0447_));
 sky130_fd_sc_hd__or2_1 _3277_ (.A(_2834_),
    .B(_2916_),
    .X(_0448_));
 sky130_fd_sc_hd__or4_1 _3278_ (.A(_2809_),
    .B(_2812_),
    .C(_2813_),
    .D(_2817_),
    .X(_0449_));
 sky130_fd_sc_hd__or3_1 _3279_ (.A(_2763_),
    .B(_2878_),
    .C(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__or4_1 _3280_ (.A(_2773_),
    .B(_2927_),
    .C(_0447_),
    .D(_0448_),
    .X(_0451_));
 sky130_fd_sc_hd__or3_1 _3281_ (.A(_2915_),
    .B(_0450_),
    .C(_0451_),
    .X(_0452_));
 sky130_fd_sc_hd__or2_1 _3282_ (.A(_2926_),
    .B(_2931_),
    .X(_0453_));
 sky130_fd_sc_hd__nor2_1 _3283_ (.A(_0397_),
    .B(_0415_),
    .Y(_0454_));
 sky130_fd_sc_hd__o21a_1 _3284_ (.A1(net150),
    .A2(_0454_),
    .B1(_2941_),
    .X(_0455_));
 sky130_fd_sc_hd__nor2_1 _3285_ (.A(_2799_),
    .B(_2919_),
    .Y(_0456_));
 sky130_fd_sc_hd__nor2_1 _3286_ (.A(net147),
    .B(_0396_),
    .Y(_0457_));
 sky130_fd_sc_hd__nand2_1 _3287_ (.A(_0385_),
    .B(_0423_),
    .Y(_0458_));
 sky130_fd_sc_hd__and2_1 _3288_ (.A(net116),
    .B(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__inv_2 _3289_ (.A(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__or3_1 _3290_ (.A(_2933_),
    .B(_0452_),
    .C(_0453_),
    .X(_0461_));
 sky130_fd_sc_hd__a2111o_1 _3291_ (.A1(_2933_),
    .A2(_2940_),
    .B1(_2814_),
    .C1(_2885_),
    .D1(_2917_),
    .X(_0462_));
 sky130_fd_sc_hd__a221o_1 _3292_ (.A1(_2920_),
    .A2(_2936_),
    .B1(_0460_),
    .B2(net97),
    .C1(_0462_),
    .X(_0463_));
 sky130_fd_sc_hd__a2bb2o_1 _3293_ (.A1_N(_0456_),
    .A2_N(_0457_),
    .B1(_0461_),
    .B2(net150),
    .X(_0464_));
 sky130_fd_sc_hd__or3_1 _3294_ (.A(_0455_),
    .B(_0463_),
    .C(_0464_),
    .X(_0465_));
 sky130_fd_sc_hd__and2b_2 _3295_ (.A_N(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .B(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ),
    .X(_0466_));
 sky130_fd_sc_hd__o21a_1 _3296_ (.A1(net144),
    .A2(_0466_),
    .B1(net117),
    .X(_0467_));
 sky130_fd_sc_hd__o21ai_1 _3297_ (.A1(net143),
    .A2(_0466_),
    .B1(net117),
    .Y(_0468_));
 sky130_fd_sc_hd__nand2_1 _3298_ (.A(_0419_),
    .B(_0468_),
    .Y(_0469_));
 sky130_fd_sc_hd__nand2_2 _3299_ (.A(_0379_),
    .B(_0396_),
    .Y(_0470_));
 sky130_fd_sc_hd__nor2_1 _3300_ (.A(net143),
    .B(_2712_),
    .Y(_0471_));
 sky130_fd_sc_hd__and2_2 _3301_ (.A(net117),
    .B(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__or2_1 _3302_ (.A(net149),
    .B(_0472_),
    .X(_0473_));
 sky130_fd_sc_hd__or2_1 _3303_ (.A(_2841_),
    .B(_0473_),
    .X(_0474_));
 sky130_fd_sc_hd__a21o_1 _3304_ (.A1(_2840_),
    .A2(_2842_),
    .B1(_0392_),
    .X(_0475_));
 sky130_fd_sc_hd__a22o_1 _3305_ (.A1(_2856_),
    .A2(_2935_),
    .B1(_0379_),
    .B2(_0457_),
    .X(_0476_));
 sky130_fd_sc_hd__and3_1 _3306_ (.A(_2855_),
    .B(_2857_),
    .C(_0380_),
    .X(_0477_));
 sky130_fd_sc_hd__nor2_1 _3307_ (.A(_0476_),
    .B(_0477_),
    .Y(_0478_));
 sky130_fd_sc_hd__a31o_1 _3308_ (.A1(_0474_),
    .A2(_0475_),
    .A3(_0478_),
    .B1(net147),
    .X(_0479_));
 sky130_fd_sc_hd__nand2_2 _3309_ (.A(net146),
    .B(_2869_),
    .Y(_0480_));
 sky130_fd_sc_hd__o21a_2 _3310_ (.A1(_2860_),
    .A2(_0480_),
    .B1(net116),
    .X(_0481_));
 sky130_fd_sc_hd__inv_2 _3311_ (.A(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__a221o_1 _3312_ (.A1(_0377_),
    .A2(_0479_),
    .B1(_0482_),
    .B2(\z80.tv80s.i_tv80_core.ISet[2] ),
    .C1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ),
    .X(_0483_));
 sky130_fd_sc_hd__a31o_1 _3313_ (.A1(net165),
    .A2(_0465_),
    .A3(_0469_),
    .B1(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__a2bb2o_1 _3314_ (.A1_N(_2934_),
    .A2_N(_2940_),
    .B1(net117),
    .B2(_2920_),
    .X(_0485_));
 sky130_fd_sc_hd__a2bb2o_1 _3315_ (.A1_N(_0396_),
    .A2_N(_0456_),
    .B1(_0458_),
    .B2(net97),
    .X(_0486_));
 sky130_fd_sc_hd__o41a_1 _3316_ (.A1(_0452_),
    .A2(_0453_),
    .A3(_0485_),
    .A4(_0486_),
    .B1(_2706_),
    .X(_0487_));
 sky130_fd_sc_hd__o211a_1 _3317_ (.A1(_0397_),
    .A2(_0415_),
    .B1(_2706_),
    .C1(_2941_),
    .X(_0488_));
 sky130_fd_sc_hd__or3b_1 _3318_ (.A(_2814_),
    .B(_2917_),
    .C_N(_0469_),
    .X(_0489_));
 sky130_fd_sc_hd__o31ai_1 _3319_ (.A1(_0487_),
    .A2(_0488_),
    .A3(_0489_),
    .B1(net165),
    .Y(_0490_));
 sky130_fd_sc_hd__nand2_1 _3320_ (.A(\z80.tv80s.i_tv80_core.ISet[2] ),
    .B(_0481_),
    .Y(_0491_));
 sky130_fd_sc_hd__or2_1 _3321_ (.A(net106),
    .B(_0479_),
    .X(_0492_));
 sky130_fd_sc_hd__a31o_1 _3322_ (.A1(_0490_),
    .A2(_0491_),
    .A3(_0492_),
    .B1(net142),
    .X(_0493_));
 sky130_fd_sc_hd__or3_1 _3323_ (.A(net118),
    .B(_2767_),
    .C(_2784_),
    .X(_0494_));
 sky130_fd_sc_hd__nand2_1 _3324_ (.A(_2792_),
    .B(_0494_),
    .Y(_0495_));
 sky130_fd_sc_hd__o31a_1 _3325_ (.A1(_0452_),
    .A2(_0485_),
    .A3(_0495_),
    .B1(_2706_),
    .X(_0496_));
 sky130_fd_sc_hd__and2_2 _3326_ (.A(net118),
    .B(_2785_),
    .X(_0497_));
 sky130_fd_sc_hd__nand2_2 _3327_ (.A(net118),
    .B(_2785_),
    .Y(_0498_));
 sky130_fd_sc_hd__nor2_1 _3328_ (.A(_2706_),
    .B(_0424_),
    .Y(_0499_));
 sky130_fd_sc_hd__nand2_1 _3329_ (.A(net150),
    .B(_0423_),
    .Y(_0500_));
 sky130_fd_sc_hd__o21a_1 _3330_ (.A1(_0459_),
    .A2(_0499_),
    .B1(net97),
    .X(_0501_));
 sky130_fd_sc_hd__o21ai_1 _3331_ (.A1(_2799_),
    .A2(_2885_),
    .B1(_0457_),
    .Y(_0502_));
 sky130_fd_sc_hd__a21o_1 _3332_ (.A1(_2792_),
    .A2(_0494_),
    .B1(_0397_),
    .X(_0503_));
 sky130_fd_sc_hd__nand2_1 _3333_ (.A(_0502_),
    .B(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__or4_1 _3334_ (.A(_0453_),
    .B(_0497_),
    .C(_0501_),
    .D(_0504_),
    .X(_0505_));
 sky130_fd_sc_hd__o31a_1 _3335_ (.A1(_0488_),
    .A2(_0496_),
    .A3(_0505_),
    .B1(net165),
    .X(_0506_));
 sky130_fd_sc_hd__o311a_1 _3336_ (.A1(net149),
    .A2(_2842_),
    .A3(_0396_),
    .B1(_2855_),
    .C1(_2841_),
    .X(_0507_));
 sky130_fd_sc_hd__and4bb_1 _3337_ (.A_N(_0476_),
    .B_N(_0477_),
    .C(_0507_),
    .D(_0403_),
    .X(_0508_));
 sky130_fd_sc_hd__a211oi_1 _3338_ (.A1(net147),
    .A2(_0477_),
    .B1(_0508_),
    .C1(net105),
    .Y(_0509_));
 sky130_fd_sc_hd__a2111o_1 _3339_ (.A1(\z80.tv80s.i_tv80_core.ISet[2] ),
    .A2(_0481_),
    .B1(_0506_),
    .C1(_0509_),
    .D1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ),
    .X(_0510_));
 sky130_fd_sc_hd__and2b_1 _3340_ (.A_N(_0493_),
    .B(_0510_),
    .X(_0511_));
 sky130_fd_sc_hd__nor2_1 _3341_ (.A(_0493_),
    .B(_0510_),
    .Y(_0512_));
 sky130_fd_sc_hd__mux2_1 _3342_ (.A0(\z80.tv80s.i_tv80_core.ts[2] ),
    .A1(net136),
    .S(_0510_),
    .X(_0513_));
 sky130_fd_sc_hd__nor3b_1 _3343_ (.A(_0484_),
    .B(_0493_),
    .C_N(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__mux2_1 _3344_ (.A0(net398),
    .A1(net255),
    .S(_0510_),
    .X(_0515_));
 sky130_fd_sc_hd__a221o_1 _3345_ (.A1(net497),
    .A2(_0512_),
    .B1(_0515_),
    .B2(_0493_),
    .C1(_0514_),
    .X(_0516_));
 sky130_fd_sc_hd__a31oi_1 _3346_ (.A1(\z80.tv80s.i_tv80_core.ts[0] ),
    .A2(_0484_),
    .A3(_0511_),
    .B1(_0516_),
    .Y(_0517_));
 sky130_fd_sc_hd__inv_6 _3347_ (.A(net54),
    .Y(_0518_));
 sky130_fd_sc_hd__nor2_4 _3348_ (.A(_2714_),
    .B(net11),
    .Y(_0519_));
 sky130_fd_sc_hd__nor2_1 _3349_ (.A(net54),
    .B(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__or3_4 _3350_ (.A(net749),
    .B(net54),
    .C(_0519_),
    .X(_0521_));
 sky130_fd_sc_hd__inv_2 _3351_ (.A(_0521_),
    .Y(_0522_));
 sky130_fd_sc_hd__nor2_1 _3352_ (.A(_0446_),
    .B(_0521_),
    .Y(_0523_));
 sky130_fd_sc_hd__or2_4 _3353_ (.A(_0446_),
    .B(_0521_),
    .X(_0524_));
 sky130_fd_sc_hd__or3_1 _3354_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ),
    .B(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .C(net267),
    .X(_0525_));
 sky130_fd_sc_hd__inv_2 _3355_ (.A(_0525_),
    .Y(_0526_));
 sky130_fd_sc_hd__or4_1 _3356_ (.A(net142),
    .B(net117),
    .C(net143),
    .D(_0525_),
    .X(_0527_));
 sky130_fd_sc_hd__a21oi_1 _3357_ (.A1(_0374_),
    .A2(_0527_),
    .B1(_0524_),
    .Y(_0528_));
 sky130_fd_sc_hd__a21o_1 _3358_ (.A1(net259),
    .A2(_0524_),
    .B1(_0528_),
    .X(_0007_));
 sky130_fd_sc_hd__and3_1 _3359_ (.A(_2697_),
    .B(_0374_),
    .C(_0523_),
    .X(_0529_));
 sky130_fd_sc_hd__and2_1 _3360_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ),
    .B(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__a21o_1 _3361_ (.A1(net273),
    .A2(_0524_),
    .B1(_0530_),
    .X(_0008_));
 sky130_fd_sc_hd__or4_1 _3362_ (.A(net142),
    .B(\z80.tv80s.i_tv80_core.BusReq_s ),
    .C(_0385_),
    .D(_0519_),
    .X(_0531_));
 sky130_fd_sc_hd__or4b_1 _3363_ (.A(_0446_),
    .B(_0525_),
    .C(_0531_),
    .D_N(_0374_),
    .X(_0532_));
 sky130_fd_sc_hd__nor2_1 _3364_ (.A(net54),
    .B(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__a21o_1 _3365_ (.A1(net261),
    .A2(_0524_),
    .B1(_0533_),
    .X(_0009_));
 sky130_fd_sc_hd__and2b_1 _3366_ (.A_N(net555),
    .B(_0529_),
    .X(_0534_));
 sky130_fd_sc_hd__a22o_1 _3367_ (.A1(net461),
    .A2(_0524_),
    .B1(_0534_),
    .B2(net267),
    .X(_0010_));
 sky130_fd_sc_hd__and3_1 _3368_ (.A(net143),
    .B(_0526_),
    .C(_0529_),
    .X(_0535_));
 sky130_fd_sc_hd__a21o_1 _3369_ (.A1(net250),
    .A2(_0524_),
    .B1(_0535_),
    .X(_0011_));
 sky130_fd_sc_hd__and3_1 _3370_ (.A(net142),
    .B(_0374_),
    .C(_0523_),
    .X(_0536_));
 sky130_fd_sc_hd__a21o_1 _3371_ (.A1(net490),
    .A2(_0524_),
    .B1(_0536_),
    .X(_0012_));
 sky130_fd_sc_hd__or2_1 _3372_ (.A(_0535_),
    .B(_0536_),
    .X(_0537_));
 sky130_fd_sc_hd__o41a_1 _3373_ (.A1(net261),
    .A2(\z80.tv80s.i_tv80_core.Pre_XY_F_M[5] ),
    .A3(net250),
    .A4(\z80.tv80s.i_tv80_core.Pre_XY_F_M[7] ),
    .B1(_0524_),
    .X(_0538_));
 sky130_fd_sc_hd__a2111o_1 _3374_ (.A1(net267),
    .A2(_0534_),
    .B1(_0537_),
    .C1(_0538_),
    .D1(_0533_),
    .X(_0029_));
 sky130_fd_sc_hd__o41a_1 _3375_ (.A1(\z80.tv80s.i_tv80_core.Pre_XY_F_M[2] ),
    .A2(\z80.tv80s.i_tv80_core.Pre_XY_F_M[3] ),
    .A3(net250),
    .A4(\z80.tv80s.i_tv80_core.Pre_XY_F_M[7] ),
    .B1(_0524_),
    .X(_0539_));
 sky130_fd_sc_hd__or4_1 _3376_ (.A(_0528_),
    .B(_0530_),
    .C(_0537_),
    .D(net251),
    .X(_0030_));
 sky130_fd_sc_hd__o31a_2 _3377_ (.A1(net136),
    .A2(\z80.tv80s.i_tv80_core.ts[1] ),
    .A3(\z80.tv80s.i_tv80_core.ts[2] ),
    .B1(net151),
    .X(_0540_));
 sky130_fd_sc_hd__o31ai_2 _3378_ (.A1(net136),
    .A2(net656),
    .A3(net870),
    .B1(net151),
    .Y(_0541_));
 sky130_fd_sc_hd__o211a_1 _3379_ (.A1(_2813_),
    .A2(_2828_),
    .B1(_2819_),
    .C1(net164),
    .X(_0542_));
 sky130_fd_sc_hd__and2b_1 _3380_ (.A_N(_2828_),
    .B(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__a21oi_1 _3381_ (.A1(net555),
    .A2(_0543_),
    .B1(net103),
    .Y(_0544_));
 sky130_fd_sc_hd__and2_4 _3382_ (.A(net859),
    .B(net11),
    .X(_0545_));
 sky130_fd_sc_hd__nand2_8 _3383_ (.A(net844),
    .B(net11),
    .Y(_0546_));
 sky130_fd_sc_hd__a211o_1 _3384_ (.A1(net103),
    .A2(_0546_),
    .B1(_0544_),
    .C1(net155),
    .X(_0547_));
 sky130_fd_sc_hd__and2_1 _3385_ (.A(net164),
    .B(_2828_),
    .X(_0548_));
 sky130_fd_sc_hd__and3_1 _3386_ (.A(net148),
    .B(net109),
    .C(_0545_),
    .X(_0549_));
 sky130_fd_sc_hd__or3_2 _3387_ (.A(net116),
    .B(net155),
    .C(_0546_),
    .X(_0550_));
 sky130_fd_sc_hd__or2_2 _3388_ (.A(_0542_),
    .B(_0548_),
    .X(_0551_));
 sky130_fd_sc_hd__or4b_1 _3389_ (.A(net163),
    .B(net586),
    .C(net309),
    .D_N(_0551_),
    .X(_0552_));
 sky130_fd_sc_hd__a22o_1 _3390_ (.A1(_2819_),
    .A2(_0548_),
    .B1(_0549_),
    .B2(_0552_),
    .X(_0553_));
 sky130_fd_sc_hd__a21o_1 _3391_ (.A1(net164),
    .A2(_0547_),
    .B1(net798),
    .X(_0000_));
 sky130_fd_sc_hd__nor2_1 _3392_ (.A(_0542_),
    .B(_0550_),
    .Y(_0554_));
 sky130_fd_sc_hd__a22o_1 _3393_ (.A1(net586),
    .A2(_0550_),
    .B1(_0554_),
    .B2(_0548_),
    .X(_0001_));
 sky130_fd_sc_hd__a21oi_1 _3394_ (.A1(_0396_),
    .A2(_0415_),
    .B1(_2942_),
    .Y(_0555_));
 sky130_fd_sc_hd__and3b_1 _3395_ (.A_N(\z80.tv80s.i_tv80_core.NMICycle ),
    .B(net97),
    .C(\z80.tv80s.i_tv80_core.IntCycle ),
    .X(_0556_));
 sky130_fd_sc_hd__or4_1 _3396_ (.A(_2799_),
    .B(_2878_),
    .C(_2885_),
    .D(_0556_),
    .X(_0557_));
 sky130_fd_sc_hd__o21a_1 _3397_ (.A1(_0555_),
    .A2(_0557_),
    .B1(net165),
    .X(_0558_));
 sky130_fd_sc_hd__nor2_1 _3398_ (.A(_2897_),
    .B(net105),
    .Y(_0559_));
 sky130_fd_sc_hd__or2_1 _3399_ (.A(net155),
    .B(_0559_),
    .X(_0560_));
 sky130_fd_sc_hd__o22a_1 _3400_ (.A1(net110),
    .A2(net420),
    .B1(_0558_),
    .B2(_0560_),
    .X(_0015_));
 sky130_fd_sc_hd__a32o_1 _3401_ (.A1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .A2(_2715_),
    .A3(_0534_),
    .B1(_0524_),
    .B2(net257),
    .X(_0006_));
 sky130_fd_sc_hd__or4_1 _3402_ (.A(net274),
    .B(_0010_),
    .C(net491),
    .D(net258),
    .X(_0031_));
 sky130_fd_sc_hd__nor2_2 _3403_ (.A(net155),
    .B(net106),
    .Y(_0561_));
 sky130_fd_sc_hd__o21a_2 _3404_ (.A1(_2845_),
    .A2(_0379_),
    .B1(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__nor2_2 _3405_ (.A(net115),
    .B(net155),
    .Y(_0563_));
 sky130_fd_sc_hd__a221o_1 _3406_ (.A1(net155),
    .A2(net452),
    .B1(_2781_),
    .B2(_0563_),
    .C1(_0562_),
    .X(_0013_));
 sky130_fd_sc_hd__a32o_1 _3407_ (.A1(_2941_),
    .A2(_0396_),
    .A3(_0415_),
    .B1(_0418_),
    .B2(_2793_),
    .X(_0564_));
 sky130_fd_sc_hd__o21a_1 _3408_ (.A1(_2933_),
    .A2(_2939_),
    .B1(_2891_),
    .X(_0565_));
 sky130_fd_sc_hd__a2111o_1 _3409_ (.A1(\z80.tv80s.i_tv80_core.NMICycle ),
    .A2(net97),
    .B1(_2920_),
    .C1(_0565_),
    .D1(_2765_),
    .X(_0566_));
 sky130_fd_sc_hd__a21oi_1 _3410_ (.A1(net146),
    .A2(_0408_),
    .B1(_2792_),
    .Y(_0567_));
 sky130_fd_sc_hd__or4_1 _3411_ (.A(_2769_),
    .B(_2785_),
    .C(_2926_),
    .D(_2929_),
    .X(_0568_));
 sky130_fd_sc_hd__or4_1 _3412_ (.A(_2773_),
    .B(_2914_),
    .C(_2927_),
    .D(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__o41a_1 _3413_ (.A1(_0564_),
    .A2(_0566_),
    .A3(_0567_),
    .A4(_0569_),
    .B1(net165),
    .X(_0570_));
 sky130_fd_sc_hd__a21oi_1 _3414_ (.A1(_2857_),
    .A2(_2895_),
    .B1(net106),
    .Y(_0571_));
 sky130_fd_sc_hd__a311o_1 _3415_ (.A1(\z80.tv80s.i_tv80_core.ISet[2] ),
    .A2(net95),
    .A3(net94),
    .B1(_0570_),
    .C1(_0571_),
    .X(_0572_));
 sky130_fd_sc_hd__mux2_1 _3416_ (.A0(net343),
    .A1(_0572_),
    .S(net110),
    .X(_0016_));
 sky130_fd_sc_hd__a311o_1 _3417_ (.A1(_2704_),
    .A2(net94),
    .A3(_2892_),
    .B1(_2916_),
    .C1(_2777_),
    .X(_0573_));
 sky130_fd_sc_hd__a31o_1 _3418_ (.A1(net96),
    .A2(_2860_),
    .A3(_2891_),
    .B1(_0573_),
    .X(_0574_));
 sky130_fd_sc_hd__a31o_1 _3419_ (.A1(net146),
    .A2(_2791_),
    .A3(_0408_),
    .B1(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__nand2_1 _3420_ (.A(net96),
    .B(net94),
    .Y(_0576_));
 sky130_fd_sc_hd__inv_2 _3421_ (.A(_0576_),
    .Y(_0577_));
 sky130_fd_sc_hd__nor2_1 _3422_ (.A(net105),
    .B(_0381_),
    .Y(_0578_));
 sky130_fd_sc_hd__a221o_1 _3423_ (.A1(net165),
    .A2(_0575_),
    .B1(_0577_),
    .B2(net163),
    .C1(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__a32o_1 _3424_ (.A1(_2834_),
    .A2(net94),
    .A3(_0563_),
    .B1(net594),
    .B2(net155),
    .X(_0580_));
 sky130_fd_sc_hd__a21o_1 _3425_ (.A1(net110),
    .A2(_0579_),
    .B1(net595),
    .X(_0014_));
 sky130_fd_sc_hd__and3_1 _3426_ (.A(net128),
    .B(net123),
    .C(_2703_),
    .X(_0581_));
 sky130_fd_sc_hd__a31o_1 _3427_ (.A1(net96),
    .A2(net94),
    .A3(_0581_),
    .B1(_2893_),
    .X(_0582_));
 sky130_fd_sc_hd__nor2_1 _3428_ (.A(_2861_),
    .B(_0576_),
    .Y(_0583_));
 sky130_fd_sc_hd__o21ai_1 _3429_ (.A1(_2893_),
    .A2(_0583_),
    .B1(_0561_),
    .Y(_0584_));
 sky130_fd_sc_hd__a22o_1 _3430_ (.A1(_0561_),
    .A2(_0582_),
    .B1(_0584_),
    .B2(net517),
    .X(_0004_));
 sky130_fd_sc_hd__a32o_1 _3431_ (.A1(_2789_),
    .A2(_0561_),
    .A3(_0577_),
    .B1(_0584_),
    .B2(net263),
    .X(_0005_));
 sky130_fd_sc_hd__and2_1 _3432_ (.A(net309),
    .B(_0550_),
    .X(_0003_));
 sky130_fd_sc_hd__and3_1 _3433_ (.A(net555),
    .B(net110),
    .C(net101),
    .X(_0585_));
 sky130_fd_sc_hd__and4_1 _3434_ (.A(net148),
    .B(_2813_),
    .C(_0545_),
    .D(_0563_),
    .X(_0586_));
 sky130_fd_sc_hd__a221o_1 _3435_ (.A1(net163),
    .A2(_0550_),
    .B1(_0585_),
    .B2(_0543_),
    .C1(_0586_),
    .X(_0002_));
 sky130_fd_sc_hd__nand2_8 _3436_ (.A(net116),
    .B(_0396_),
    .Y(_0587_));
 sky130_fd_sc_hd__a21oi_1 _3437_ (.A1(_2838_),
    .A2(_2843_),
    .B1(_0587_),
    .Y(_0588_));
 sky130_fd_sc_hd__a21oi_2 _3438_ (.A1(_2712_),
    .A2(_2715_),
    .B1(_0385_),
    .Y(_0589_));
 sky130_fd_sc_hd__nor2_1 _3439_ (.A(net126),
    .B(_2897_),
    .Y(_0590_));
 sky130_fd_sc_hd__a221o_1 _3440_ (.A1(_2890_),
    .A2(_0430_),
    .B1(_0589_),
    .B2(_0590_),
    .C1(net105),
    .X(_0591_));
 sky130_fd_sc_hd__a211o_1 _3441_ (.A1(_0379_),
    .A2(_0472_),
    .B1(_0588_),
    .C1(_0591_),
    .X(_0592_));
 sky130_fd_sc_hd__a21o_1 _3442_ (.A1(net118),
    .A2(_2878_),
    .B1(_2799_),
    .X(_0593_));
 sky130_fd_sc_hd__o21a_1 _3443_ (.A1(_2941_),
    .A2(_0593_),
    .B1(_0589_),
    .X(_0594_));
 sky130_fd_sc_hd__o211a_1 _3444_ (.A1(_2934_),
    .A2(_2935_),
    .B1(_0565_),
    .C1(net144),
    .X(_0595_));
 sky130_fd_sc_hd__a221o_1 _3445_ (.A1(_0419_),
    .A2(_0467_),
    .B1(_0472_),
    .B2(_0398_),
    .C1(_0595_),
    .X(_0596_));
 sky130_fd_sc_hd__nand2_1 _3446_ (.A(net116),
    .B(_0385_),
    .Y(_0597_));
 sky130_fd_sc_hd__a21o_1 _3447_ (.A1(net97),
    .A2(_0423_),
    .B1(_2926_),
    .X(_0598_));
 sky130_fd_sc_hd__nor2_1 _3448_ (.A(net126),
    .B(_2778_),
    .Y(_0599_));
 sky130_fd_sc_hd__o211a_1 _3449_ (.A1(_2702_),
    .A2(net116),
    .B1(_0599_),
    .C1(net145),
    .X(_0600_));
 sky130_fd_sc_hd__a211o_1 _3450_ (.A1(_2769_),
    .A2(_0396_),
    .B1(_0594_),
    .C1(_0600_),
    .X(_0601_));
 sky130_fd_sc_hd__a31o_1 _3451_ (.A1(net116),
    .A2(_0385_),
    .A3(_0598_),
    .B1(_0596_),
    .X(_0602_));
 sky130_fd_sc_hd__a21o_1 _3452_ (.A1(_2860_),
    .A2(_2940_),
    .B1(net95),
    .X(_0603_));
 sky130_fd_sc_hd__o311a_1 _3453_ (.A1(net96),
    .A2(_0601_),
    .A3(_0602_),
    .B1(_0603_),
    .C1(net165),
    .X(_0604_));
 sky130_fd_sc_hd__nor2_1 _3454_ (.A(net142),
    .B(_0587_),
    .Y(_0605_));
 sky130_fd_sc_hd__a41o_1 _3455_ (.A1(net163),
    .A2(net95),
    .A3(net94),
    .A4(_0605_),
    .B1(net107),
    .X(_0606_));
 sky130_fd_sc_hd__o21ai_4 _3456_ (.A1(_0604_),
    .A2(_0606_),
    .B1(_0592_),
    .Y(net21));
 sky130_fd_sc_hd__or3b_1 _3457_ (.A(net105),
    .B(_0587_),
    .C_N(_2845_),
    .X(_0607_));
 sky130_fd_sc_hd__o21a_1 _3458_ (.A1(net784),
    .A2(_2840_),
    .B1(_2711_),
    .X(_0608_));
 sky130_fd_sc_hd__a31o_1 _3459_ (.A1(net784),
    .A2(_2839_),
    .A3(_2843_),
    .B1(_0608_),
    .X(_0609_));
 sky130_fd_sc_hd__a21oi_1 _3460_ (.A1(net125),
    .A2(_0609_),
    .B1(_0607_),
    .Y(_0028_));
 sky130_fd_sc_hd__nor2_1 _3461_ (.A(net656),
    .B(_0519_),
    .Y(_0610_));
 sky130_fd_sc_hd__o21ai_1 _3462_ (.A1(net746),
    .A2(_0610_),
    .B1(net150),
    .Y(_0611_));
 sky130_fd_sc_hd__nor2_2 _3463_ (.A(_2921_),
    .B(_0384_),
    .Y(_0612_));
 sky130_fd_sc_hd__o21ai_4 _3464_ (.A1(_0498_),
    .A2(_0587_),
    .B1(_0503_),
    .Y(_0613_));
 sky130_fd_sc_hd__o21a_1 _3465_ (.A1(_0612_),
    .A2(_0613_),
    .B1(net165),
    .X(_0614_));
 sky130_fd_sc_hd__nor2_1 _3466_ (.A(_0610_),
    .B(_0614_),
    .Y(_0615_));
 sky130_fd_sc_hd__nor2_2 _3467_ (.A(net143),
    .B(_2936_),
    .Y(_0616_));
 sky130_fd_sc_hd__a2111o_1 _3468_ (.A1(_2838_),
    .A2(_2843_),
    .B1(_2936_),
    .C1(_2712_),
    .D1(net143),
    .X(_0617_));
 sky130_fd_sc_hd__nor2_2 _3469_ (.A(_2857_),
    .B(_0384_),
    .Y(_0618_));
 sky130_fd_sc_hd__o31ai_1 _3470_ (.A1(net147),
    .A2(_2839_),
    .A3(_0393_),
    .B1(_0617_),
    .Y(_0619_));
 sky130_fd_sc_hd__a311oi_1 _3471_ (.A1(net126),
    .A2(net145),
    .A3(_0379_),
    .B1(_0618_),
    .C1(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hd__o2bb2a_1 _3472_ (.A1_N(net142),
    .A2_N(_0374_),
    .B1(_0620_),
    .B2(net164),
    .X(_0621_));
 sky130_fd_sc_hd__o211a_1 _3473_ (.A1(net805),
    .A2(_0621_),
    .B1(_0615_),
    .C1(net21),
    .X(_0622_));
 sky130_fd_sc_hd__o21ai_1 _3474_ (.A1(net150),
    .A2(_0622_),
    .B1(_0611_),
    .Y(_0019_));
 sky130_fd_sc_hd__a21o_1 _3475_ (.A1(_2842_),
    .A2(_0381_),
    .B1(_0431_),
    .X(_0623_));
 sky130_fd_sc_hd__o21a_1 _3476_ (.A1(_2841_),
    .A2(_0587_),
    .B1(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__or3_1 _3477_ (.A(_2883_),
    .B(_2925_),
    .C(_2927_),
    .X(_0625_));
 sky130_fd_sc_hd__nor2_1 _3478_ (.A(_2880_),
    .B(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__or3_1 _3479_ (.A(_2914_),
    .B(_2919_),
    .C(_2931_),
    .X(_0627_));
 sky130_fd_sc_hd__or2_1 _3480_ (.A(_2809_),
    .B(_2917_),
    .X(_0628_));
 sky130_fd_sc_hd__or2_1 _3481_ (.A(_2817_),
    .B(_0628_),
    .X(_0629_));
 sky130_fd_sc_hd__a2111o_1 _3482_ (.A1(net124),
    .A2(_2812_),
    .B1(_2831_),
    .C1(net96),
    .D1(_2939_),
    .X(_0630_));
 sky130_fd_sc_hd__or4_1 _3483_ (.A(_2783_),
    .B(_2823_),
    .C(_0629_),
    .D(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__or3_1 _3484_ (.A(_2763_),
    .B(_2768_),
    .C(_2920_),
    .X(_0632_));
 sky130_fd_sc_hd__inv_2 _3485_ (.A(_0632_),
    .Y(_0633_));
 sky130_fd_sc_hd__or3_1 _3486_ (.A(_2886_),
    .B(_2933_),
    .C(_0448_),
    .X(_0634_));
 sky130_fd_sc_hd__nand2_1 _3487_ (.A(net165),
    .B(_0396_),
    .Y(_0635_));
 sky130_fd_sc_hd__or3_1 _3488_ (.A(_2768_),
    .B(_2920_),
    .C(_0635_),
    .X(_0636_));
 sky130_fd_sc_hd__o32a_1 _3489_ (.A1(_0633_),
    .A2(_0634_),
    .A3(_0636_),
    .B1(_0624_),
    .B2(net106),
    .X(_0637_));
 sky130_fd_sc_hd__o21ba_1 _3490_ (.A1(net21),
    .A2(_0610_),
    .B1_N(_0622_),
    .X(_0638_));
 sky130_fd_sc_hd__or2_1 _3491_ (.A(_0637_),
    .B(_0638_),
    .X(_0639_));
 sky130_fd_sc_hd__o21ai_1 _3492_ (.A1(net656),
    .A2(_0519_),
    .B1(net746),
    .Y(_0640_));
 sky130_fd_sc_hd__mux2_1 _3493_ (.A0(_0639_),
    .A1(_0640_),
    .S(net150),
    .X(_0017_));
 sky130_fd_sc_hd__and2b_1 _3494_ (.A_N(_0638_),
    .B(_0637_),
    .X(_0641_));
 sky130_fd_sc_hd__o21ai_1 _3495_ (.A1(net150),
    .A2(_0641_),
    .B1(_0611_),
    .Y(_0018_));
 sky130_fd_sc_hd__or3_4 _3496_ (.A(net115),
    .B(_2935_),
    .C(_0498_),
    .X(_0642_));
 sky130_fd_sc_hd__or4_1 _3497_ (.A(\z80.tv80s.i_tv80_core.mcycles[1] ),
    .B(\z80.tv80s.i_tv80_core.mcycles[4] ),
    .C(\z80.tv80s.i_tv80_core.mcycles[2] ),
    .D(\z80.tv80s.i_tv80_core.mcycles[5] ),
    .X(_0643_));
 sky130_fd_sc_hd__nor2_1 _3498_ (.A(_2706_),
    .B(_0643_),
    .Y(_0644_));
 sky130_fd_sc_hd__a221o_1 _3499_ (.A1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .A2(\z80.tv80s.i_tv80_core.mcycles[1] ),
    .B1(\z80.tv80s.i_tv80_core.mcycles[2] ),
    .B2(net145),
    .C1(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__a221o_2 _3500_ (.A1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ),
    .A2(\z80.tv80s.i_tv80_core.mcycles[4] ),
    .B1(\z80.tv80s.i_tv80_core.mcycles[5] ),
    .B2(net143),
    .C1(_0645_),
    .X(_0646_));
 sky130_fd_sc_hd__a41o_1 _3501_ (.A1(net146),
    .A2(net166),
    .A3(\z80.tv80s.i_tv80_core.IncDecZ ),
    .A4(_0497_),
    .B1(_0646_),
    .X(_0647_));
 sky130_fd_sc_hd__nor2_1 _3502_ (.A(net862),
    .B(_0647_),
    .Y(_0648_));
 sky130_fd_sc_hd__or4_1 _3503_ (.A(net142),
    .B(\z80.tv80s.i_tv80_core.BusReq_s ),
    .C(_0519_),
    .D(_0648_),
    .X(_0649_));
 sky130_fd_sc_hd__or3b_4 _3504_ (.A(_0649_),
    .B(net54),
    .C_N(_0446_),
    .X(_0650_));
 sky130_fd_sc_hd__a31o_1 _3505_ (.A1(net150),
    .A2(\z80.tv80s.i_tv80_core.ts[2] ),
    .A3(net11),
    .B1(net720),
    .X(_0651_));
 sky130_fd_sc_hd__and3b_1 _3506_ (.A_N(net716),
    .B(_0650_),
    .C(net721),
    .X(_0032_));
 sky130_fd_sc_hd__or4_2 _3507_ (.A(net118),
    .B(net115),
    .C(_2756_),
    .D(_2808_),
    .X(_0652_));
 sky130_fd_sc_hd__and3_1 _3508_ (.A(net662),
    .B(\z80.tv80s.i_tv80_core.INT_s ),
    .C(_0652_),
    .X(_0653_));
 sky130_fd_sc_hd__nor2_1 _3509_ (.A(_0551_),
    .B(_0650_),
    .Y(_0654_));
 sky130_fd_sc_hd__o21a_1 _3510_ (.A1(net504),
    .A2(_0653_),
    .B1(_0654_),
    .X(_0655_));
 sky130_fd_sc_hd__and4_1 _3511_ (.A(net166),
    .B(net136),
    .C(_2757_),
    .D(_2807_),
    .X(_0656_));
 sky130_fd_sc_hd__or3_2 _3512_ (.A(_2895_),
    .B(net106),
    .C(_0587_),
    .X(_0657_));
 sky130_fd_sc_hd__or3_1 _3513_ (.A(_2714_),
    .B(\z80.tv80s.i_tv80_core.IntE_FF2 ),
    .C(_0657_),
    .X(_0658_));
 sky130_fd_sc_hd__o21ai_1 _3514_ (.A1(net519),
    .A2(_0652_),
    .B1(_0657_),
    .Y(_0659_));
 sky130_fd_sc_hd__a21o_1 _3515_ (.A1(\z80.tv80s.i_tv80_core.ts[2] ),
    .A2(_0659_),
    .B1(net662),
    .X(_0660_));
 sky130_fd_sc_hd__and4bb_1 _3516_ (.A_N(_0655_),
    .B_N(_0656_),
    .C(_0658_),
    .D(net663),
    .X(_0026_));
 sky130_fd_sc_hd__or4b_1 _3517_ (.A(net504),
    .B(_0551_),
    .C(_0650_),
    .D_N(_0653_),
    .X(_0661_));
 sky130_fd_sc_hd__o21bai_1 _3518_ (.A1(_2714_),
    .A2(_0652_),
    .B1_N(net828),
    .Y(_0662_));
 sky130_fd_sc_hd__and3b_1 _3519_ (.A_N(_0656_),
    .B(_0661_),
    .C(net829),
    .X(_0027_));
 sky130_fd_sc_hd__a21oi_2 _3520_ (.A1(net155),
    .A2(net749),
    .B1(_0519_),
    .Y(_0663_));
 sky130_fd_sc_hd__and4_1 _3521_ (.A(net165),
    .B(net96),
    .C(net94),
    .D(_2891_),
    .X(_0664_));
 sky130_fd_sc_hd__a32o_1 _3522_ (.A1(_0518_),
    .A2(_0663_),
    .A3(_0664_),
    .B1(_0424_),
    .B2(net619),
    .X(_0024_));
 sky130_fd_sc_hd__nor2_1 _3523_ (.A(net515),
    .B(_0637_),
    .Y(_0665_));
 sky130_fd_sc_hd__o21a_1 _3524_ (.A1(_0499_),
    .A2(_0665_),
    .B1(net54),
    .X(_0021_));
 sky130_fd_sc_hd__or3_1 _3525_ (.A(net150),
    .B(net21),
    .C(_0610_),
    .X(_0020_));
 sky130_fd_sc_hd__and2_1 _3526_ (.A(net450),
    .B(net54),
    .X(_0022_));
 sky130_fd_sc_hd__nand2_1 _3527_ (.A(net382),
    .B(net413),
    .Y(_0666_));
 sky130_fd_sc_hd__nand2_1 _3528_ (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ),
    .B(net542),
    .Y(_0667_));
 sky130_fd_sc_hd__nand2_1 _3529_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .B(net154),
    .Y(_0668_));
 sky130_fd_sc_hd__nand3_4 _3530_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .C(net154),
    .Y(_0669_));
 sky130_fd_sc_hd__nor2_1 _3531_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .B(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__or2_2 _3532_ (.A(_2713_),
    .B(net450),
    .X(_0671_));
 sky130_fd_sc_hd__mux2_2 _3533_ (.A0(_0670_),
    .A1(_0671_),
    .S(_2719_),
    .X(_0672_));
 sky130_fd_sc_hd__nor2_1 _3534_ (.A(_0666_),
    .B(_0672_),
    .Y(_0673_));
 sky130_fd_sc_hd__or4b_2 _3535_ (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ),
    .B(_0672_),
    .C(_0666_),
    .D_N(_0667_),
    .X(_0674_));
 sky130_fd_sc_hd__and3_1 _3536_ (.A(net164),
    .B(net136),
    .C(_2881_),
    .X(_0675_));
 sky130_fd_sc_hd__nand3_4 _3537_ (.A(net164),
    .B(net136),
    .C(_2881_),
    .Y(_0676_));
 sky130_fd_sc_hd__and3_2 _3538_ (.A(net167),
    .B(\z80.tv80s.i_tv80_core.ts[4] ),
    .C(_2881_),
    .X(_0677_));
 sky130_fd_sc_hd__nand3_4 _3539_ (.A(net167),
    .B(net398),
    .C(_2881_),
    .Y(_0678_));
 sky130_fd_sc_hd__or2_1 _3540_ (.A(net147),
    .B(_0468_),
    .X(_0679_));
 sky130_fd_sc_hd__a21o_1 _3541_ (.A1(_2885_),
    .A2(_0679_),
    .B1(net115),
    .X(_0680_));
 sky130_fd_sc_hd__nor2_1 _3542_ (.A(_2942_),
    .B(_0417_),
    .Y(_0681_));
 sky130_fd_sc_hd__nand2_1 _3543_ (.A(_2926_),
    .B(_2936_),
    .Y(_0682_));
 sky130_fd_sc_hd__a32o_1 _3544_ (.A1(_2768_),
    .A2(_2936_),
    .A3(_0423_),
    .B1(_0392_),
    .B2(_2799_),
    .X(_0683_));
 sky130_fd_sc_hd__nor2_2 _3545_ (.A(_2885_),
    .B(_0683_),
    .Y(_0684_));
 sky130_fd_sc_hd__a21o_1 _3546_ (.A1(_2928_),
    .A2(_2930_),
    .B1(_0597_),
    .X(_0685_));
 sky130_fd_sc_hd__o311a_1 _3547_ (.A1(_2942_),
    .A2(_0393_),
    .A3(_0416_),
    .B1(_0682_),
    .C1(_0685_),
    .X(_0686_));
 sky130_fd_sc_hd__nand2_1 _3548_ (.A(net122),
    .B(_2917_),
    .Y(_0687_));
 sky130_fd_sc_hd__a31o_1 _3549_ (.A1(_0684_),
    .A2(_0686_),
    .A3(_0687_),
    .B1(_0680_),
    .X(_0688_));
 sky130_fd_sc_hd__a21o_1 _3550_ (.A1(_2841_),
    .A2(_2895_),
    .B1(_0597_),
    .X(_0689_));
 sky130_fd_sc_hd__o221a_1 _3551_ (.A1(_2840_),
    .A2(_0431_),
    .B1(_0587_),
    .B2(_2842_),
    .C1(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__o21a_1 _3552_ (.A1(net105),
    .A2(_0690_),
    .B1(_0688_),
    .X(_0691_));
 sky130_fd_sc_hd__o21ai_2 _3553_ (.A1(net105),
    .A2(_0690_),
    .B1(_0688_),
    .Y(_0692_));
 sky130_fd_sc_hd__or2_1 _3554_ (.A(_2895_),
    .B(_0597_),
    .X(_0693_));
 sky130_fd_sc_hd__o21a_1 _3555_ (.A1(_2838_),
    .A2(_0587_),
    .B1(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__nand2_1 _3556_ (.A(net125),
    .B(_2917_),
    .Y(_0695_));
 sky130_fd_sc_hd__a31o_1 _3557_ (.A1(_0684_),
    .A2(_0686_),
    .A3(_0695_),
    .B1(_0680_),
    .X(_0696_));
 sky130_fd_sc_hd__o21ai_4 _3558_ (.A1(net105),
    .A2(_0694_),
    .B1(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__nand2_1 _3559_ (.A(_0692_),
    .B(_0697_),
    .Y(_0698_));
 sky130_fd_sc_hd__a31o_1 _3560_ (.A1(_2918_),
    .A2(_0684_),
    .A3(_0686_),
    .B1(_0680_),
    .X(_0699_));
 sky130_fd_sc_hd__o21a_1 _3561_ (.A1(_2756_),
    .A2(_2836_),
    .B1(net145),
    .X(_0700_));
 sky130_fd_sc_hd__o21ai_1 _3562_ (.A1(net147),
    .A2(_0700_),
    .B1(_2839_),
    .Y(_0701_));
 sky130_fd_sc_hd__nand2_1 _3563_ (.A(_2842_),
    .B(_2935_),
    .Y(_0702_));
 sky130_fd_sc_hd__a21oi_1 _3564_ (.A1(_0701_),
    .A2(_0702_),
    .B1(_2837_),
    .Y(_0703_));
 sky130_fd_sc_hd__o211a_1 _3565_ (.A1(_0616_),
    .A2(_0703_),
    .B1(_0693_),
    .C1(net107),
    .X(_0704_));
 sky130_fd_sc_hd__a21oi_2 _3566_ (.A1(net105),
    .A2(_0699_),
    .B1(_0704_),
    .Y(_0705_));
 sky130_fd_sc_hd__nand2_1 _3567_ (.A(net148),
    .B(net136),
    .Y(_0706_));
 sky130_fd_sc_hd__o21ai_1 _3568_ (.A1(net148),
    .A2(_0546_),
    .B1(_0706_),
    .Y(_0707_));
 sky130_fd_sc_hd__nand3_2 _3569_ (.A(_0698_),
    .B(_0705_),
    .C(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__a41o_4 _3570_ (.A1(_0674_),
    .A2(_0676_),
    .A3(_0678_),
    .A4(_0708_),
    .B1(net157),
    .X(_0709_));
 sky130_fd_sc_hd__a211o_2 _3571_ (.A1(net105),
    .A2(_0699_),
    .B1(_0704_),
    .C1(_0706_),
    .X(_0710_));
 sky130_fd_sc_hd__a21oi_4 _3572_ (.A1(_2714_),
    .A2(_0710_),
    .B1(net104),
    .Y(_0711_));
 sky130_fd_sc_hd__or3_2 _3573_ (.A(net90),
    .B(_0677_),
    .C(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__o31ai_2 _3574_ (.A1(net90),
    .A2(_0677_),
    .A3(_0711_),
    .B1(_2718_),
    .Y(_0713_));
 sky130_fd_sc_hd__a21oi_1 _3575_ (.A1(_2714_),
    .A2(_0710_),
    .B1(_0697_),
    .Y(_0714_));
 sky130_fd_sc_hd__a211oi_4 _3576_ (.A1(_2714_),
    .A2(_0710_),
    .B1(_0697_),
    .C1(_0691_),
    .Y(_0715_));
 sky130_fd_sc_hd__mux2_1 _3577_ (.A0(\z80.tv80s.i_tv80_core.RegAddrA_r[2] ),
    .A1(\z80.tv80s.i_tv80_core.XY_State[1] ),
    .S(_0715_),
    .X(_0716_));
 sky130_fd_sc_hd__o21a_4 _3578_ (.A1(_0712_),
    .A2(_0716_),
    .B1(_0713_),
    .X(_0717_));
 sky130_fd_sc_hd__o21ai_2 _3579_ (.A1(_0712_),
    .A2(_0716_),
    .B1(_0713_),
    .Y(_0718_));
 sky130_fd_sc_hd__a21o_1 _3580_ (.A1(\z80.tv80s.i_tv80_core.RegAddrA_r[1] ),
    .A2(net89),
    .B1(net90),
    .X(_0719_));
 sky130_fd_sc_hd__a211o_1 _3581_ (.A1(_2714_),
    .A2(_0710_),
    .B1(_0692_),
    .C1(net104),
    .X(_0720_));
 sky130_fd_sc_hd__o31ai_4 _3582_ (.A1(_0711_),
    .A2(_0715_),
    .A3(_0719_),
    .B1(_0720_),
    .Y(_0721_));
 sky130_fd_sc_hd__o31a_2 _3583_ (.A1(_0711_),
    .A2(_0715_),
    .A3(_0719_),
    .B1(_0720_),
    .X(_0722_));
 sky130_fd_sc_hd__o21a_4 _3584_ (.A1(\z80.tv80s.i_tv80_core.RegAddrA_r[0] ),
    .A2(_0677_),
    .B1(_0676_),
    .X(_0723_));
 sky130_fd_sc_hd__a211o_4 _3585_ (.A1(_2714_),
    .A2(_0710_),
    .B1(_0697_),
    .C1(net104),
    .X(_0724_));
 sky130_fd_sc_hd__o31ai_4 _3586_ (.A1(_0711_),
    .A2(net75),
    .A3(_0723_),
    .B1(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__o31a_4 _3587_ (.A1(_0711_),
    .A2(net75),
    .A3(_0723_),
    .B1(_0724_),
    .X(_0726_));
 sky130_fd_sc_hd__and3_4 _3588_ (.A(_0717_),
    .B(net71),
    .C(net70),
    .X(_0727_));
 sky130_fd_sc_hd__or3_4 _3589_ (.A(net65),
    .B(net72),
    .C(net69),
    .X(_0728_));
 sky130_fd_sc_hd__nor2_4 _3590_ (.A(_0709_),
    .B(_0728_),
    .Y(_0729_));
 sky130_fd_sc_hd__nor2_1 _3591_ (.A(net140),
    .B(net90),
    .Y(_0730_));
 sky130_fd_sc_hd__nand2_1 _3592_ (.A(_2718_),
    .B(net90),
    .Y(_0731_));
 sky130_fd_sc_hd__o21a_1 _3593_ (.A1(\z80.tv80s.i_tv80_core.RegAddrB_r[2] ),
    .A2(net90),
    .B1(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__o21ai_2 _3594_ (.A1(\z80.tv80s.i_tv80_core.RegAddrB_r[2] ),
    .A2(net90),
    .B1(_0731_),
    .Y(_0733_));
 sky130_fd_sc_hd__mux4_1 _3595_ (.A0(net406),
    .A1(net434),
    .A2(net303),
    .A3(net301),
    .S0(net82),
    .S1(net81),
    .X(_0734_));
 sky130_fd_sc_hd__o21ai_1 _3596_ (.A1(net148),
    .A2(_2714_),
    .B1(_0706_),
    .Y(_0735_));
 sky130_fd_sc_hd__and2_2 _3597_ (.A(_0705_),
    .B(_0735_),
    .X(_0736_));
 sky130_fd_sc_hd__nand2_2 _3598_ (.A(_0705_),
    .B(_0735_),
    .Y(_0737_));
 sky130_fd_sc_hd__and3_4 _3599_ (.A(net65),
    .B(net72),
    .C(net70),
    .X(_0738_));
 sky130_fd_sc_hd__or3_1 _3600_ (.A(_0717_),
    .B(net71),
    .C(net69),
    .X(_0739_));
 sky130_fd_sc_hd__and3_4 _3601_ (.A(net65),
    .B(net72),
    .C(net69),
    .X(_0740_));
 sky130_fd_sc_hd__or3_1 _3602_ (.A(_0717_),
    .B(net71),
    .C(net70),
    .X(_0741_));
 sky130_fd_sc_hd__and3_4 _3603_ (.A(net65),
    .B(net71),
    .C(net70),
    .X(_0742_));
 sky130_fd_sc_hd__or3_1 _3604_ (.A(_0717_),
    .B(net72),
    .C(net69),
    .X(_0743_));
 sky130_fd_sc_hd__and3_4 _3605_ (.A(net65),
    .B(net71),
    .C(net69),
    .X(_0744_));
 sky130_fd_sc_hd__or3_1 _3606_ (.A(_0717_),
    .B(net72),
    .C(_0725_),
    .X(_0745_));
 sky130_fd_sc_hd__mux2_1 _3607_ (.A0(net406),
    .A1(net434),
    .S(net70),
    .X(_0746_));
 sky130_fd_sc_hd__o311a_1 _3608_ (.A1(_0711_),
    .A2(net75),
    .A3(_0723_),
    .B1(_0724_),
    .C1(_2716_),
    .X(_0747_));
 sky130_fd_sc_hd__a211oi_1 _3609_ (.A1(_2717_),
    .A2(net70),
    .B1(_0747_),
    .C1(net72),
    .Y(_0748_));
 sky130_fd_sc_hd__a211o_1 _3610_ (.A1(net72),
    .A2(_0746_),
    .B1(_0748_),
    .C1(_0717_),
    .X(_0749_));
 sky130_fd_sc_hd__and3_4 _3611_ (.A(_0717_),
    .B(net72),
    .C(_0725_),
    .X(_0750_));
 sky130_fd_sc_hd__or3_4 _3612_ (.A(net65),
    .B(net71),
    .C(net69),
    .X(_0751_));
 sky130_fd_sc_hd__and3_4 _3613_ (.A(_0717_),
    .B(net72),
    .C(net69),
    .X(_0752_));
 sky130_fd_sc_hd__or3_4 _3614_ (.A(net65),
    .B(net71),
    .C(_0725_),
    .X(_0753_));
 sky130_fd_sc_hd__and3_4 _3615_ (.A(_0717_),
    .B(net71),
    .C(net69),
    .X(_0754_));
 sky130_fd_sc_hd__or3_4 _3616_ (.A(net65),
    .B(net72),
    .C(_0725_),
    .X(_0755_));
 sky130_fd_sc_hd__mux2_1 _3617_ (.A0(net303),
    .A1(net301),
    .S(net70),
    .X(_0756_));
 sky130_fd_sc_hd__mux2_1 _3618_ (.A0(net347),
    .A1(net333),
    .S(net70),
    .X(_0757_));
 sky130_fd_sc_hd__mux2_1 _3619_ (.A0(_0756_),
    .A1(_0757_),
    .S(net71),
    .X(_0758_));
 sky130_fd_sc_hd__o21a_1 _3620_ (.A1(net65),
    .A2(_0758_),
    .B1(_0749_),
    .X(_0759_));
 sky130_fd_sc_hd__o21ai_4 _3621_ (.A1(net65),
    .A2(_0758_),
    .B1(_0749_),
    .Y(_0760_));
 sky130_fd_sc_hd__and3_4 _3622_ (.A(net166),
    .B(net96),
    .C(_2909_),
    .X(_0761_));
 sky130_fd_sc_hd__and2_1 _3623_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .B(_0669_),
    .X(_0762_));
 sky130_fd_sc_hd__nand2_4 _3624_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .B(_0669_),
    .Y(_0763_));
 sky130_fd_sc_hd__and2b_2 _3625_ (.A_N(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .B(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .X(_0764_));
 sky130_fd_sc_hd__xor2_2 _3626_ (.A(net154),
    .B(\z80.tv80s.i_tv80_core.BusB[0] ),
    .X(_0765_));
 sky130_fd_sc_hd__and2_1 _3627_ (.A(\z80.tv80s.i_tv80_core.BusA[0] ),
    .B(_0765_),
    .X(_0766_));
 sky130_fd_sc_hd__or2_1 _3628_ (.A(net154),
    .B(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__xor2_2 _3629_ (.A(\z80.tv80s.i_tv80_core.BusA[0] ),
    .B(_0765_),
    .X(_0768_));
 sky130_fd_sc_hd__and2b_1 _3630_ (.A_N(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(\z80.tv80s.i_tv80_core.F[0] ),
    .X(_0769_));
 sky130_fd_sc_hd__nor2_1 _3631_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .B(net154),
    .Y(_0770_));
 sky130_fd_sc_hd__or2_1 _3632_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .B(net154),
    .X(_0771_));
 sky130_fd_sc_hd__xor2_1 _3633_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .B(net154),
    .X(_0772_));
 sky130_fd_sc_hd__mux2_1 _3634_ (.A0(net154),
    .A1(_0772_),
    .S(_0769_),
    .X(_0773_));
 sky130_fd_sc_hd__or2_1 _3635_ (.A(_0768_),
    .B(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__nand2_1 _3636_ (.A(_0768_),
    .B(_0773_),
    .Y(_0775_));
 sky130_fd_sc_hd__and2_2 _3637_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(_0668_),
    .X(_0776_));
 sky130_fd_sc_hd__nand2_4 _3638_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(_0668_),
    .Y(_0777_));
 sky130_fd_sc_hd__and3_2 _3639_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .C(net108),
    .X(_0778_));
 sky130_fd_sc_hd__a22o_1 _3640_ (.A1(_0764_),
    .A2(_0767_),
    .B1(_0768_),
    .B2(_0778_),
    .X(_0779_));
 sky130_fd_sc_hd__a31o_1 _3641_ (.A1(_0774_),
    .A2(_0775_),
    .A3(_0777_),
    .B1(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__o41a_2 _3642_ (.A1(net108),
    .A2(\z80.tv80s.i_tv80_core.BusA[0] ),
    .A3(\z80.tv80s.i_tv80_core.BusB[0] ),
    .A4(_0777_),
    .B1(_0780_),
    .X(_0781_));
 sky130_fd_sc_hd__nor2_1 _3643_ (.A(net120),
    .B(_2787_),
    .Y(_0782_));
 sky130_fd_sc_hd__and3b_1 _3644_ (.A_N(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(\z80.tv80s.i_tv80_core.ALU_Op_r[1] ),
    .C(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .X(_0783_));
 sky130_fd_sc_hd__and2b_4 _3645_ (.A_N(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .B(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__and4b_4 _3646_ (.A_N(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .C(net108),
    .D(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .X(_0785_));
 sky130_fd_sc_hd__and3_2 _3647_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .B(_0771_),
    .C(_0776_),
    .X(_0786_));
 sky130_fd_sc_hd__inv_2 _3648_ (.A(_0786_),
    .Y(_0787_));
 sky130_fd_sc_hd__mux2_1 _3649_ (.A0(\z80.tv80s.i_tv80_core.BusB[0] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[4] ),
    .S(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .X(_0788_));
 sky130_fd_sc_hd__and3_2 _3650_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .B(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .C(_0770_),
    .X(_0789_));
 sky130_fd_sc_hd__nand3_2 _3651_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .B(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .C(_0770_),
    .Y(_0790_));
 sky130_fd_sc_hd__and3b_4 _3652_ (.A_N(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(_0770_),
    .C(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .X(_0791_));
 sky130_fd_sc_hd__a221o_1 _3653_ (.A1(net123),
    .A2(\z80.tv80s.i_tv80_core.F[0] ),
    .B1(net139),
    .B2(_2750_),
    .C1(_2805_),
    .X(_0792_));
 sky130_fd_sc_hd__mux2_1 _3654_ (.A0(\z80.tv80s.i_tv80_core.BusA[1] ),
    .A1(_0792_),
    .S(net119),
    .X(_0793_));
 sky130_fd_sc_hd__nand2_2 _3655_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .B(_0783_),
    .Y(_0794_));
 sky130_fd_sc_hd__inv_2 _3656_ (.A(_0794_),
    .Y(_0795_));
 sky130_fd_sc_hd__nor2_1 _3657_ (.A(_0782_),
    .B(_0794_),
    .Y(_0796_));
 sky130_fd_sc_hd__a211o_1 _3658_ (.A1(_0782_),
    .A2(_0785_),
    .B1(_0796_),
    .C1(_0784_),
    .X(_0797_));
 sky130_fd_sc_hd__a22o_1 _3659_ (.A1(_0782_),
    .A2(_0784_),
    .B1(_0786_),
    .B2(_0788_),
    .X(_0798_));
 sky130_fd_sc_hd__a211o_1 _3660_ (.A1(\z80.tv80s.i_tv80_core.BusA[0] ),
    .A2(_0789_),
    .B1(_0798_),
    .C1(_0763_),
    .X(_0799_));
 sky130_fd_sc_hd__a22o_1 _3661_ (.A1(_0791_),
    .A2(_0793_),
    .B1(_0797_),
    .B2(\z80.tv80s.i_tv80_core.BusB[0] ),
    .X(_0800_));
 sky130_fd_sc_hd__o221a_1 _3662_ (.A1(_0762_),
    .A2(_0781_),
    .B1(_0799_),
    .B2(_0800_),
    .C1(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(_0801_));
 sky130_fd_sc_hd__a21o_1 _3663_ (.A1(_2719_),
    .A2(\z80.tv80s.di_reg[0] ),
    .B1(_0801_),
    .X(_0802_));
 sky130_fd_sc_hd__mux2_4 _3664_ (.A0(_0802_),
    .A1(net580),
    .S(_0761_),
    .X(_0803_));
 sky130_fd_sc_hd__a21oi_1 _3665_ (.A1(net74),
    .A2(_0803_),
    .B1(_0677_),
    .Y(_0804_));
 sky130_fd_sc_hd__o21ai_1 _3666_ (.A1(net74),
    .A2(_0759_),
    .B1(_0804_),
    .Y(_0805_));
 sky130_fd_sc_hd__a21oi_1 _3667_ (.A1(_2748_),
    .A2(_0677_),
    .B1(net90),
    .Y(_0806_));
 sky130_fd_sc_hd__a22o_2 _3668_ (.A1(net90),
    .A2(_0734_),
    .B1(_0805_),
    .B2(_0806_),
    .X(_0807_));
 sky130_fd_sc_hd__mux2_1 _3669_ (.A0(net333),
    .A1(_0807_),
    .S(_0729_),
    .X(_0036_));
 sky130_fd_sc_hd__and2_4 _3670_ (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ),
    .B(_0676_),
    .X(_0808_));
 sky130_fd_sc_hd__nand2_4 _3671_ (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ),
    .B(_0676_),
    .Y(_0809_));
 sky130_fd_sc_hd__mux2_1 _3672_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ),
    .S(net82),
    .X(_0810_));
 sky130_fd_sc_hd__mux2_1 _3673_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][1] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][1] ),
    .S(net82),
    .X(_0811_));
 sky130_fd_sc_hd__mux2_1 _3674_ (.A0(_0810_),
    .A1(_0811_),
    .S(net79),
    .X(_0812_));
 sky130_fd_sc_hd__o221a_1 _3675_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][1] ),
    .A2(net140),
    .B1(net82),
    .B2(net875),
    .C1(net81),
    .X(_0813_));
 sky130_fd_sc_hd__o221a_1 _3676_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ),
    .A2(net140),
    .B1(net82),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ),
    .C1(net79),
    .X(_0814_));
 sky130_fd_sc_hd__or3_1 _3677_ (.A(_0809_),
    .B(_0813_),
    .C(_0814_),
    .X(_0815_));
 sky130_fd_sc_hd__o21a_1 _3678_ (.A1(_0808_),
    .A2(_0812_),
    .B1(_0815_),
    .X(_0816_));
 sky130_fd_sc_hd__and2b_1 _3679_ (.A_N(\z80.tv80s.i_tv80_core.BusB[1] ),
    .B(net154),
    .X(_0817_));
 sky130_fd_sc_hd__and2b_1 _3680_ (.A_N(net154),
    .B(\z80.tv80s.i_tv80_core.BusB[1] ),
    .X(_0818_));
 sky130_fd_sc_hd__o21ai_1 _3681_ (.A1(_0817_),
    .A2(_0818_),
    .B1(\z80.tv80s.i_tv80_core.BusA[1] ),
    .Y(_0819_));
 sky130_fd_sc_hd__nand2_1 _3682_ (.A(net108),
    .B(_0819_),
    .Y(_0820_));
 sky130_fd_sc_hd__or3_1 _3683_ (.A(\z80.tv80s.i_tv80_core.BusA[1] ),
    .B(_0817_),
    .C(_0818_),
    .X(_0821_));
 sky130_fd_sc_hd__and2_1 _3684_ (.A(_0819_),
    .B(_0821_),
    .X(_0822_));
 sky130_fd_sc_hd__a21o_1 _3685_ (.A1(_0768_),
    .A2(_0773_),
    .B1(_0766_),
    .X(_0823_));
 sky130_fd_sc_hd__or2_1 _3686_ (.A(_0822_),
    .B(_0823_),
    .X(_0824_));
 sky130_fd_sc_hd__nand2_1 _3687_ (.A(_0822_),
    .B(_0823_),
    .Y(_0825_));
 sky130_fd_sc_hd__a22o_1 _3688_ (.A1(_0764_),
    .A2(_0820_),
    .B1(_0822_),
    .B2(_0778_),
    .X(_0826_));
 sky130_fd_sc_hd__a31o_1 _3689_ (.A1(_0777_),
    .A2(_0824_),
    .A3(_0825_),
    .B1(_0826_),
    .X(_0827_));
 sky130_fd_sc_hd__o41a_2 _3690_ (.A1(net108),
    .A2(\z80.tv80s.i_tv80_core.BusA[1] ),
    .A3(\z80.tv80s.i_tv80_core.BusB[1] ),
    .A4(_0777_),
    .B1(_0827_),
    .X(_0828_));
 sky130_fd_sc_hd__mux2_1 _3691_ (.A0(\z80.tv80s.i_tv80_core.BusB[1] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[5] ),
    .S(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .X(_0829_));
 sky130_fd_sc_hd__mux2_1 _3692_ (.A0(\z80.tv80s.i_tv80_core.BusA[0] ),
    .A1(\z80.tv80s.i_tv80_core.BusA[2] ),
    .S(net129),
    .X(_0830_));
 sky130_fd_sc_hd__a22o_1 _3693_ (.A1(_0786_),
    .A2(_0829_),
    .B1(_0830_),
    .B2(_0791_),
    .X(_0831_));
 sky130_fd_sc_hd__and3_1 _3694_ (.A(net127),
    .B(_2702_),
    .C(_2703_),
    .X(_0832_));
 sky130_fd_sc_hd__nor2_1 _3695_ (.A(_0794_),
    .B(_0832_),
    .Y(_0833_));
 sky130_fd_sc_hd__a211o_1 _3696_ (.A1(_0785_),
    .A2(_0832_),
    .B1(_0833_),
    .C1(_0784_),
    .X(_0834_));
 sky130_fd_sc_hd__a221o_1 _3697_ (.A1(_0784_),
    .A2(_0832_),
    .B1(_0834_),
    .B2(\z80.tv80s.i_tv80_core.BusB[1] ),
    .C1(_0831_),
    .X(_0835_));
 sky130_fd_sc_hd__o21a_1 _3698_ (.A1(\z80.tv80s.i_tv80_core.BusA[1] ),
    .A2(\z80.tv80s.i_tv80_core.BusA[2] ),
    .B1(\z80.tv80s.i_tv80_core.BusA[3] ),
    .X(_0836_));
 sky130_fd_sc_hd__o21ai_1 _3699_ (.A1(\z80.tv80s.i_tv80_core.BusA[1] ),
    .A2(\z80.tv80s.i_tv80_core.BusA[2] ),
    .B1(\z80.tv80s.i_tv80_core.BusA[3] ),
    .Y(_0837_));
 sky130_fd_sc_hd__nor2_1 _3700_ (.A(\z80.tv80s.i_tv80_core.F[4] ),
    .B(_0836_),
    .Y(_0838_));
 sky130_fd_sc_hd__or2_1 _3701_ (.A(\z80.tv80s.i_tv80_core.BusA[3] ),
    .B(\z80.tv80s.i_tv80_core.F[4] ),
    .X(_0839_));
 sky130_fd_sc_hd__mux2_1 _3702_ (.A0(_0838_),
    .A1(_0839_),
    .S(\z80.tv80s.i_tv80_core.BusA[1] ),
    .X(_0840_));
 sky130_fd_sc_hd__a2bb2o_1 _3703_ (.A1_N(_0790_),
    .A2_N(_0840_),
    .B1(_0828_),
    .B2(_0763_),
    .X(_0841_));
 sky130_fd_sc_hd__nor2_1 _3704_ (.A(_0835_),
    .B(_0841_),
    .Y(_0842_));
 sky130_fd_sc_hd__inv_2 _3705_ (.A(_0842_),
    .Y(_0843_));
 sky130_fd_sc_hd__mux2_1 _3706_ (.A0(\z80.tv80s.di_reg[1] ),
    .A1(_0843_),
    .S(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(_0844_));
 sky130_fd_sc_hd__mux2_4 _3707_ (.A0(_0844_),
    .A1(net701),
    .S(_0761_),
    .X(_0845_));
 sky130_fd_sc_hd__a21o_1 _3708_ (.A1(net74),
    .A2(_0845_),
    .B1(_0677_),
    .X(_0846_));
 sky130_fd_sc_hd__nand2_1 _3709_ (.A(net126),
    .B(_2917_),
    .Y(_0847_));
 sky130_fd_sc_hd__o311a_1 _3710_ (.A1(_2942_),
    .A2(_0393_),
    .A3(_0416_),
    .B1(_0682_),
    .C1(_0847_),
    .X(_0848_));
 sky130_fd_sc_hd__nand2_1 _3711_ (.A(_0466_),
    .B(_0616_),
    .Y(_0849_));
 sky130_fd_sc_hd__a221oi_4 _3712_ (.A1(_0684_),
    .A2(_0848_),
    .B1(_0849_),
    .B2(_2885_),
    .C1(net115),
    .Y(_0850_));
 sky130_fd_sc_hd__nand2_1 _3713_ (.A(_2843_),
    .B(_2935_),
    .Y(_0851_));
 sky130_fd_sc_hd__a21o_1 _3714_ (.A1(_0701_),
    .A2(_0851_),
    .B1(_2837_),
    .X(_0852_));
 sky130_fd_sc_hd__nor2_1 _3715_ (.A(net127),
    .B(net150),
    .Y(_0853_));
 sky130_fd_sc_hd__a21o_1 _3716_ (.A1(net126),
    .A2(_0385_),
    .B1(net148),
    .X(_0854_));
 sky130_fd_sc_hd__a31o_2 _3717_ (.A1(net107),
    .A2(_0852_),
    .A3(_0854_),
    .B1(_0850_),
    .X(_0855_));
 sky130_fd_sc_hd__inv_4 _3718_ (.A(net77),
    .Y(_0856_));
 sky130_fd_sc_hd__o311a_1 _3719_ (.A1(_0711_),
    .A2(net75),
    .A3(_0723_),
    .B1(_0724_),
    .C1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ),
    .X(_0857_));
 sky130_fd_sc_hd__o311a_1 _3720_ (.A1(_0711_),
    .A2(net75),
    .A3(_0723_),
    .B1(_0724_),
    .C1(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][1] ),
    .X(_0858_));
 sky130_fd_sc_hd__a211o_1 _3721_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ),
    .A2(net70),
    .B1(_0857_),
    .C1(net71),
    .X(_0859_));
 sky130_fd_sc_hd__a211o_1 _3722_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][1] ),
    .A2(net70),
    .B1(_0858_),
    .C1(net72),
    .X(_0860_));
 sky130_fd_sc_hd__a21o_1 _3723_ (.A1(_0859_),
    .A2(_0860_),
    .B1(net65),
    .X(_0861_));
 sky130_fd_sc_hd__mux2_1 _3724_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][1] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][1] ),
    .S(net70),
    .X(_0862_));
 sky130_fd_sc_hd__o311a_1 _3725_ (.A1(_0711_),
    .A2(net75),
    .A3(_0723_),
    .B1(_0724_),
    .C1(_2720_),
    .X(_0863_));
 sky130_fd_sc_hd__a211oi_1 _3726_ (.A1(_2721_),
    .A2(net70),
    .B1(_0863_),
    .C1(net72),
    .Y(_0864_));
 sky130_fd_sc_hd__a211o_1 _3727_ (.A1(net72),
    .A2(_0862_),
    .B1(_0864_),
    .C1(_0717_),
    .X(_0865_));
 sky130_fd_sc_hd__nand2_1 _3728_ (.A(_0861_),
    .B(_0865_),
    .Y(_0866_));
 sky130_fd_sc_hd__inv_2 _3729_ (.A(_0866_),
    .Y(_0867_));
 sky130_fd_sc_hd__and3_1 _3730_ (.A(net77),
    .B(_0861_),
    .C(_0865_),
    .X(_0868_));
 sky130_fd_sc_hd__a21o_1 _3731_ (.A1(_0861_),
    .A2(_0865_),
    .B1(net77),
    .X(_0869_));
 sky130_fd_sc_hd__nand2b_1 _3732_ (.A_N(_0868_),
    .B(_0869_),
    .Y(_0870_));
 sky130_fd_sc_hd__nor2_1 _3733_ (.A(_0760_),
    .B(_0870_),
    .Y(_0871_));
 sky130_fd_sc_hd__a21o_1 _3734_ (.A1(_0760_),
    .A2(_0870_),
    .B1(net74),
    .X(_0872_));
 sky130_fd_sc_hd__o21bai_1 _3735_ (.A1(_0871_),
    .A2(_0872_),
    .B1_N(_0846_),
    .Y(_0873_));
 sky130_fd_sc_hd__o21a_1 _3736_ (.A1(net228),
    .A2(net89),
    .B1(_0676_),
    .X(_0874_));
 sky130_fd_sc_hd__a22o_2 _3737_ (.A1(net90),
    .A2(net876),
    .B1(_0873_),
    .B2(_0874_),
    .X(_0875_));
 sky130_fd_sc_hd__mux2_1 _3738_ (.A0(net408),
    .A1(_0875_),
    .S(_0729_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _3739_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ),
    .S(net85),
    .X(_0876_));
 sky130_fd_sc_hd__mux2_1 _3740_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ),
    .S(net82),
    .X(_0877_));
 sky130_fd_sc_hd__mux2_1 _3741_ (.A0(_0876_),
    .A1(_0877_),
    .S(net79),
    .X(_0878_));
 sky130_fd_sc_hd__o221a_1 _3742_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ),
    .A2(net140),
    .B1(net85),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ),
    .C1(net81),
    .X(_0879_));
 sky130_fd_sc_hd__o221a_1 _3743_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ),
    .A2(net140),
    .B1(net85),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ),
    .C1(net79),
    .X(_0880_));
 sky130_fd_sc_hd__or3_1 _3744_ (.A(_0809_),
    .B(_0879_),
    .C(_0880_),
    .X(_0881_));
 sky130_fd_sc_hd__o21a_1 _3745_ (.A1(_0808_),
    .A2(_0878_),
    .B1(_0881_),
    .X(_0882_));
 sky130_fd_sc_hd__a21o_1 _3746_ (.A1(_0759_),
    .A2(_0869_),
    .B1(_0868_),
    .X(_0883_));
 sky130_fd_sc_hd__mux2_1 _3747_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ),
    .S(net69),
    .X(_0884_));
 sky130_fd_sc_hd__nor2_1 _3748_ (.A(net71),
    .B(_0884_),
    .Y(_0885_));
 sky130_fd_sc_hd__mux2_1 _3749_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ),
    .S(net69),
    .X(_0886_));
 sky130_fd_sc_hd__o21ai_1 _3750_ (.A1(net72),
    .A2(_0886_),
    .B1(_0717_),
    .Y(_0887_));
 sky130_fd_sc_hd__mux2_1 _3751_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ),
    .S(net69),
    .X(_0888_));
 sky130_fd_sc_hd__mux2_1 _3752_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ),
    .S(net69),
    .X(_0889_));
 sky130_fd_sc_hd__mux2_1 _3753_ (.A0(_0888_),
    .A1(_0889_),
    .S(net71),
    .X(_0890_));
 sky130_fd_sc_hd__o2bb2a_2 _3754_ (.A1_N(net65),
    .A2_N(_0890_),
    .B1(_0887_),
    .B2(_0885_),
    .X(_0891_));
 sky130_fd_sc_hd__inv_2 _3755_ (.A(_0891_),
    .Y(_0892_));
 sky130_fd_sc_hd__nor2_1 _3756_ (.A(_0856_),
    .B(_0891_),
    .Y(_0893_));
 sky130_fd_sc_hd__xnor2_2 _3757_ (.A(net77),
    .B(_0891_),
    .Y(_0894_));
 sky130_fd_sc_hd__nand2_1 _3758_ (.A(_0883_),
    .B(_0894_),
    .Y(_0895_));
 sky130_fd_sc_hd__or2_1 _3759_ (.A(_0883_),
    .B(_0894_),
    .X(_0896_));
 sky130_fd_sc_hd__nor2_1 _3760_ (.A(net108),
    .B(\z80.tv80s.i_tv80_core.BusB[2] ),
    .Y(_0897_));
 sky130_fd_sc_hd__nor2_1 _3761_ (.A(net154),
    .B(_2726_),
    .Y(_0898_));
 sky130_fd_sc_hd__o21ai_1 _3762_ (.A1(_0897_),
    .A2(_0898_),
    .B1(\z80.tv80s.i_tv80_core.BusA[2] ),
    .Y(_0899_));
 sky130_fd_sc_hd__nand2_1 _3763_ (.A(net108),
    .B(_0899_),
    .Y(_0900_));
 sky130_fd_sc_hd__or3_1 _3764_ (.A(\z80.tv80s.i_tv80_core.BusA[2] ),
    .B(_0897_),
    .C(_0898_),
    .X(_0901_));
 sky130_fd_sc_hd__and2_1 _3765_ (.A(_0899_),
    .B(_0901_),
    .X(_0902_));
 sky130_fd_sc_hd__a21bo_1 _3766_ (.A1(_0822_),
    .A2(_0823_),
    .B1_N(_0819_),
    .X(_0903_));
 sky130_fd_sc_hd__xnor2_1 _3767_ (.A(_0902_),
    .B(_0903_),
    .Y(_0904_));
 sky130_fd_sc_hd__a22o_1 _3768_ (.A1(_0764_),
    .A2(_0900_),
    .B1(_0902_),
    .B2(_0778_),
    .X(_0905_));
 sky130_fd_sc_hd__o21ba_1 _3769_ (.A1(_0776_),
    .A2(_0904_),
    .B1_N(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__a31o_1 _3770_ (.A1(_2725_),
    .A2(_0776_),
    .A3(_0897_),
    .B1(_0906_),
    .X(_0907_));
 sky130_fd_sc_hd__mux2_1 _3771_ (.A0(\z80.tv80s.i_tv80_core.F[1] ),
    .A1(_2724_),
    .S(_0838_),
    .X(_0908_));
 sky130_fd_sc_hd__xor2_1 _3772_ (.A(\z80.tv80s.i_tv80_core.BusA[1] ),
    .B(\z80.tv80s.i_tv80_core.BusA[2] ),
    .X(_0909_));
 sky130_fd_sc_hd__xnor2_2 _3773_ (.A(_0908_),
    .B(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__mux2_1 _3774_ (.A0(\z80.tv80s.i_tv80_core.BusB[2] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[6] ),
    .S(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .X(_0911_));
 sky130_fd_sc_hd__mux2_1 _3775_ (.A0(\z80.tv80s.i_tv80_core.BusA[1] ),
    .A1(\z80.tv80s.i_tv80_core.BusA[3] ),
    .S(net129),
    .X(_0912_));
 sky130_fd_sc_hd__a221o_1 _3776_ (.A1(_0786_),
    .A2(_0911_),
    .B1(_0912_),
    .B2(_0791_),
    .C1(_0763_),
    .X(_0913_));
 sky130_fd_sc_hd__nor2_1 _3777_ (.A(net127),
    .B(_2761_),
    .Y(_0914_));
 sky130_fd_sc_hd__nor2_1 _3778_ (.A(_0794_),
    .B(_0914_),
    .Y(_0915_));
 sky130_fd_sc_hd__a211o_1 _3779_ (.A1(_0785_),
    .A2(_0914_),
    .B1(_0915_),
    .C1(_0784_),
    .X(_0916_));
 sky130_fd_sc_hd__a22o_1 _3780_ (.A1(_0789_),
    .A2(_0910_),
    .B1(_0916_),
    .B2(\z80.tv80s.i_tv80_core.BusB[2] ),
    .X(_0917_));
 sky130_fd_sc_hd__a211o_1 _3781_ (.A1(_0784_),
    .A2(_0914_),
    .B1(_0917_),
    .C1(_0913_),
    .X(_0918_));
 sky130_fd_sc_hd__a21bo_1 _3782_ (.A1(_0763_),
    .A2(_0907_),
    .B1_N(_0918_),
    .X(_0919_));
 sky130_fd_sc_hd__mux2_1 _3783_ (.A0(_2735_),
    .A1(_0919_),
    .S(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(_0920_));
 sky130_fd_sc_hd__mux2_2 _3784_ (.A0(_0920_),
    .A1(_2726_),
    .S(_0761_),
    .X(_0921_));
 sky130_fd_sc_hd__inv_2 _3785_ (.A(_0921_),
    .Y(_0922_));
 sky130_fd_sc_hd__o21ai_1 _3786_ (.A1(_0736_),
    .A2(_0921_),
    .B1(net89),
    .Y(_0923_));
 sky130_fd_sc_hd__a31o_1 _3787_ (.A1(_0736_),
    .A2(_0895_),
    .A3(_0896_),
    .B1(_0923_),
    .X(_0924_));
 sky130_fd_sc_hd__o21a_1 _3788_ (.A1(net224),
    .A2(net89),
    .B1(_0676_),
    .X(_0925_));
 sky130_fd_sc_hd__a22o_2 _3789_ (.A1(net90),
    .A2(_0882_),
    .B1(_0924_),
    .B2(_0925_),
    .X(_0926_));
 sky130_fd_sc_hd__mux2_1 _3790_ (.A0(net457),
    .A1(_0926_),
    .S(_0729_),
    .X(_0038_));
 sky130_fd_sc_hd__a22o_1 _3791_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][3] ),
    .A2(_0738_),
    .B1(_0740_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][3] ),
    .X(_0927_));
 sky130_fd_sc_hd__a22o_1 _3792_ (.A1(net329),
    .A2(_0750_),
    .B1(_0752_),
    .B2(net380),
    .X(_0928_));
 sky130_fd_sc_hd__and4_1 _3793_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ),
    .B(net65),
    .C(_0722_),
    .D(_0725_),
    .X(_0929_));
 sky130_fd_sc_hd__and4_1 _3794_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ),
    .B(net65),
    .C(_0722_),
    .D(_0726_),
    .X(_0930_));
 sky130_fd_sc_hd__and4_1 _3795_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][3] ),
    .B(_0717_),
    .C(_0722_),
    .D(_0726_),
    .X(_0931_));
 sky130_fd_sc_hd__a2111o_1 _3796_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ),
    .A2(_0727_),
    .B1(_0929_),
    .C1(_0930_),
    .D1(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__or3_2 _3797_ (.A(_0927_),
    .B(_0928_),
    .C(_0932_),
    .X(_0933_));
 sky130_fd_sc_hd__or4_1 _3798_ (.A(net77),
    .B(_0927_),
    .C(_0928_),
    .D(_0932_),
    .X(_0934_));
 sky130_fd_sc_hd__o31a_1 _3799_ (.A1(_0927_),
    .A2(_0928_),
    .A3(_0932_),
    .B1(net77),
    .X(_0935_));
 sky130_fd_sc_hd__xnor2_1 _3800_ (.A(net77),
    .B(_0933_),
    .Y(_0936_));
 sky130_fd_sc_hd__a21oi_1 _3801_ (.A1(_0883_),
    .A2(_0894_),
    .B1(_0893_),
    .Y(_0937_));
 sky130_fd_sc_hd__xnor2_1 _3802_ (.A(_0936_),
    .B(_0937_),
    .Y(_0938_));
 sky130_fd_sc_hd__nor2_1 _3803_ (.A(net74),
    .B(_0938_),
    .Y(_0939_));
 sky130_fd_sc_hd__nor2_1 _3804_ (.A(net108),
    .B(\z80.tv80s.i_tv80_core.BusB[3] ),
    .Y(_0940_));
 sky130_fd_sc_hd__nor2_1 _3805_ (.A(net154),
    .B(_2727_),
    .Y(_0941_));
 sky130_fd_sc_hd__o21a_1 _3806_ (.A1(_0940_),
    .A2(_0941_),
    .B1(\z80.tv80s.i_tv80_core.BusA[3] ),
    .X(_0942_));
 sky130_fd_sc_hd__or2_1 _3807_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[1] ),
    .B(_0942_),
    .X(_0943_));
 sky130_fd_sc_hd__nor3_1 _3808_ (.A(\z80.tv80s.i_tv80_core.BusA[3] ),
    .B(_0940_),
    .C(_0941_),
    .Y(_0944_));
 sky130_fd_sc_hd__nor2_1 _3809_ (.A(_0942_),
    .B(_0944_),
    .Y(_0945_));
 sky130_fd_sc_hd__a21bo_1 _3810_ (.A1(_0902_),
    .A2(_0903_),
    .B1_N(_0899_),
    .X(_0946_));
 sky130_fd_sc_hd__or2_1 _3811_ (.A(_0945_),
    .B(_0946_),
    .X(_0947_));
 sky130_fd_sc_hd__a21oi_1 _3812_ (.A1(_0945_),
    .A2(_0946_),
    .B1(_0776_),
    .Y(_0948_));
 sky130_fd_sc_hd__a22o_1 _3813_ (.A1(_0764_),
    .A2(_0943_),
    .B1(_0945_),
    .B2(_0778_),
    .X(_0949_));
 sky130_fd_sc_hd__a21o_1 _3814_ (.A1(_0947_),
    .A2(_0948_),
    .B1(_0949_),
    .X(_0950_));
 sky130_fd_sc_hd__o41a_2 _3815_ (.A1(net108),
    .A2(\z80.tv80s.i_tv80_core.BusA[3] ),
    .A3(\z80.tv80s.i_tv80_core.BusB[3] ),
    .A4(_0777_),
    .B1(_0950_),
    .X(_0951_));
 sky130_fd_sc_hd__a21o_1 _3816_ (.A1(\z80.tv80s.i_tv80_core.BusA[1] ),
    .A2(\z80.tv80s.i_tv80_core.BusA[2] ),
    .B1(\z80.tv80s.i_tv80_core.BusA[3] ),
    .X(_0952_));
 sky130_fd_sc_hd__a31oi_1 _3817_ (.A1(\z80.tv80s.i_tv80_core.BusA[1] ),
    .A2(\z80.tv80s.i_tv80_core.BusA[2] ),
    .A3(\z80.tv80s.i_tv80_core.BusA[3] ),
    .B1(_0838_),
    .Y(_0953_));
 sky130_fd_sc_hd__or3_1 _3818_ (.A(\z80.tv80s.i_tv80_core.BusA[1] ),
    .B(\z80.tv80s.i_tv80_core.BusA[2] ),
    .C(\z80.tv80s.i_tv80_core.BusA[3] ),
    .X(_0954_));
 sky130_fd_sc_hd__a21o_1 _3819_ (.A1(_0837_),
    .A2(_0954_),
    .B1(\z80.tv80s.i_tv80_core.F[1] ),
    .X(_0955_));
 sky130_fd_sc_hd__nand2_1 _3820_ (.A(_0839_),
    .B(_0955_),
    .Y(_0956_));
 sky130_fd_sc_hd__a31o_1 _3821_ (.A1(\z80.tv80s.i_tv80_core.F[1] ),
    .A2(_0952_),
    .A3(_0953_),
    .B1(_0956_),
    .X(_0957_));
 sky130_fd_sc_hd__mux2_1 _3822_ (.A0(\z80.tv80s.i_tv80_core.BusB[3] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[7] ),
    .S(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .X(_0958_));
 sky130_fd_sc_hd__mux2_1 _3823_ (.A0(\z80.tv80s.i_tv80_core.BusA[2] ),
    .A1(\z80.tv80s.i_tv80_core.BusA[4] ),
    .S(net129),
    .X(_0959_));
 sky130_fd_sc_hd__and2_1 _3824_ (.A(_0791_),
    .B(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__a2bb2o_1 _3825_ (.A1_N(_0790_),
    .A2_N(_0957_),
    .B1(_0958_),
    .B2(_0786_),
    .X(_0961_));
 sky130_fd_sc_hd__mux2_1 _3826_ (.A0(_0795_),
    .A1(_0785_),
    .S(_0581_),
    .X(_0962_));
 sky130_fd_sc_hd__or2_1 _3827_ (.A(\z80.tv80s.i_tv80_core.BusB[3] ),
    .B(_0581_),
    .X(_0963_));
 sky130_fd_sc_hd__a221o_1 _3828_ (.A1(net790),
    .A2(_0962_),
    .B1(_0963_),
    .B2(_0784_),
    .C1(_0960_),
    .X(_0964_));
 sky130_fd_sc_hd__a211oi_2 _3829_ (.A1(_0763_),
    .A2(_0951_),
    .B1(_0961_),
    .C1(_0964_),
    .Y(_0965_));
 sky130_fd_sc_hd__mux2_1 _3830_ (.A0(_2734_),
    .A1(_0965_),
    .S(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(_0966_));
 sky130_fd_sc_hd__mux2_2 _3831_ (.A0(_0966_),
    .A1(_2727_),
    .S(_0761_),
    .X(_0967_));
 sky130_fd_sc_hd__inv_2 _3832_ (.A(_0967_),
    .Y(_0968_));
 sky130_fd_sc_hd__o21ai_1 _3833_ (.A1(_0736_),
    .A2(_0967_),
    .B1(net89),
    .Y(_0969_));
 sky130_fd_sc_hd__o221a_1 _3834_ (.A1(net236),
    .A2(net89),
    .B1(_0939_),
    .B2(_0969_),
    .C1(_0676_),
    .X(_0970_));
 sky130_fd_sc_hd__mux4_2 _3835_ (.A0(net414),
    .A1(net380),
    .A2(net454),
    .A3(net329),
    .S0(net81),
    .S1(net82),
    .X(_0971_));
 sky130_fd_sc_hd__a21o_2 _3836_ (.A1(net90),
    .A2(_0971_),
    .B1(_0970_),
    .X(_0972_));
 sky130_fd_sc_hd__mux2_1 _3837_ (.A0(net439),
    .A1(_0972_),
    .S(_0729_),
    .X(_0039_));
 sky130_fd_sc_hd__nand2_1 _3838_ (.A(\z80.tv80s.i_tv80_core.F[1] ),
    .B(\z80.tv80s.i_tv80_core.F[4] ),
    .Y(_0973_));
 sky130_fd_sc_hd__o22a_1 _3839_ (.A1(\z80.tv80s.i_tv80_core.F[1] ),
    .A2(_0837_),
    .B1(_0952_),
    .B2(_0973_),
    .X(_0974_));
 sky130_fd_sc_hd__xor2_2 _3840_ (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .B(_0974_),
    .X(_0975_));
 sky130_fd_sc_hd__a21o_1 _3841_ (.A1(\z80.tv80s.i_tv80_core.BusB[4] ),
    .A2(_0783_),
    .B1(_0409_),
    .X(_0976_));
 sky130_fd_sc_hd__o21a_1 _3842_ (.A1(_0410_),
    .A2(_0785_),
    .B1(\z80.tv80s.i_tv80_core.BusB[4] ),
    .X(_0977_));
 sky130_fd_sc_hd__o21a_1 _3843_ (.A1(_0784_),
    .A2(_0977_),
    .B1(_0976_),
    .X(_0978_));
 sky130_fd_sc_hd__mux2_1 _3844_ (.A0(\z80.tv80s.i_tv80_core.BusA[3] ),
    .A1(\z80.tv80s.i_tv80_core.BusA[5] ),
    .S(net129),
    .X(_0979_));
 sky130_fd_sc_hd__a221o_1 _3845_ (.A1(\z80.tv80s.i_tv80_core.BusA[4] ),
    .A2(_0786_),
    .B1(_0791_),
    .B2(_0979_),
    .C1(_0978_),
    .X(_0980_));
 sky130_fd_sc_hd__o21ba_1 _3846_ (.A1(_0790_),
    .A2(_0975_),
    .B1_N(_0980_),
    .X(_0981_));
 sky130_fd_sc_hd__nor2_1 _3847_ (.A(net108),
    .B(\z80.tv80s.i_tv80_core.BusB[4] ),
    .Y(_0982_));
 sky130_fd_sc_hd__or3b_1 _3848_ (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .B(_0777_),
    .C_N(_0982_),
    .X(_0983_));
 sky130_fd_sc_hd__nor2_1 _3849_ (.A(net154),
    .B(_2728_),
    .Y(_0984_));
 sky130_fd_sc_hd__o21ai_1 _3850_ (.A1(_0982_),
    .A2(_0984_),
    .B1(\z80.tv80s.i_tv80_core.BusA[4] ),
    .Y(_0985_));
 sky130_fd_sc_hd__or3_1 _3851_ (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .B(_0982_),
    .C(_0984_),
    .X(_0986_));
 sky130_fd_sc_hd__and2_1 _3852_ (.A(_0985_),
    .B(_0986_),
    .X(_0987_));
 sky130_fd_sc_hd__a21o_1 _3853_ (.A1(_0945_),
    .A2(_0946_),
    .B1(_0942_),
    .X(_0988_));
 sky130_fd_sc_hd__or2_1 _3854_ (.A(_0987_),
    .B(_0988_),
    .X(_0989_));
 sky130_fd_sc_hd__nand2_1 _3855_ (.A(_0987_),
    .B(_0988_),
    .Y(_0990_));
 sky130_fd_sc_hd__nand2_1 _3856_ (.A(net108),
    .B(_0985_),
    .Y(_0991_));
 sky130_fd_sc_hd__a22o_1 _3857_ (.A1(_0778_),
    .A2(_0987_),
    .B1(_0991_),
    .B2(_0764_),
    .X(_0992_));
 sky130_fd_sc_hd__a31o_1 _3858_ (.A1(_0777_),
    .A2(_0989_),
    .A3(_0990_),
    .B1(_0992_),
    .X(_0993_));
 sky130_fd_sc_hd__nand2_1 _3859_ (.A(_0983_),
    .B(_0993_),
    .Y(_0994_));
 sky130_fd_sc_hd__inv_2 _3860_ (.A(_0994_),
    .Y(_0995_));
 sky130_fd_sc_hd__o21a_1 _3861_ (.A1(_0762_),
    .A2(_0994_),
    .B1(_0981_),
    .X(_0996_));
 sky130_fd_sc_hd__mux2_1 _3862_ (.A0(_2736_),
    .A1(_0996_),
    .S(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(_0997_));
 sky130_fd_sc_hd__mux2_2 _3863_ (.A0(_0997_),
    .A1(_2728_),
    .S(_0761_),
    .X(_0998_));
 sky130_fd_sc_hd__inv_2 _3864_ (.A(_0998_),
    .Y(_0999_));
 sky130_fd_sc_hd__o21ai_2 _3865_ (.A1(_0736_),
    .A2(_0998_),
    .B1(_0678_),
    .Y(_1000_));
 sky130_fd_sc_hd__a311o_1 _3866_ (.A1(_0883_),
    .A2(_0894_),
    .A3(_0934_),
    .B1(_0935_),
    .C1(_0893_),
    .X(_1001_));
 sky130_fd_sc_hd__a22o_1 _3867_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][4] ),
    .A2(_0738_),
    .B1(_0740_),
    .B2(net313),
    .X(_1002_));
 sky130_fd_sc_hd__a22o_1 _3868_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ),
    .A2(_0742_),
    .B1(_0744_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ),
    .X(_1003_));
 sky130_fd_sc_hd__mux2_1 _3869_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][4] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][4] ),
    .S(_0726_),
    .X(_1004_));
 sky130_fd_sc_hd__mux2_1 _3870_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ),
    .S(_0726_),
    .X(_1005_));
 sky130_fd_sc_hd__o21a_1 _3871_ (.A1(_0721_),
    .A2(_1005_),
    .B1(_0717_),
    .X(_1006_));
 sky130_fd_sc_hd__o21a_1 _3872_ (.A1(_0722_),
    .A2(_1004_),
    .B1(_1006_),
    .X(_1007_));
 sky130_fd_sc_hd__or3_2 _3873_ (.A(_1002_),
    .B(_1003_),
    .C(_1007_),
    .X(_1008_));
 sky130_fd_sc_hd__and2_1 _3874_ (.A(net77),
    .B(_1008_),
    .X(_1009_));
 sky130_fd_sc_hd__xnor2_1 _3875_ (.A(_0856_),
    .B(_1008_),
    .Y(_1010_));
 sky130_fd_sc_hd__xnor2_1 _3876_ (.A(_1001_),
    .B(_1010_),
    .Y(_1011_));
 sky130_fd_sc_hd__nor2_1 _3877_ (.A(net74),
    .B(_1011_),
    .Y(_1012_));
 sky130_fd_sc_hd__o22a_1 _3878_ (.A1(net230),
    .A2(net89),
    .B1(_1000_),
    .B2(_1012_),
    .X(_1013_));
 sky130_fd_sc_hd__mux4_1 _3879_ (.A0(net313),
    .A1(net337),
    .A2(net422),
    .A3(net277),
    .S0(net80),
    .S1(net83),
    .X(_1014_));
 sky130_fd_sc_hd__mux2_2 _3880_ (.A0(_1013_),
    .A1(_1014_),
    .S(net90),
    .X(_1015_));
 sky130_fd_sc_hd__mux2_1 _3881_ (.A0(net372),
    .A1(_1015_),
    .S(_0729_),
    .X(_0040_));
 sky130_fd_sc_hd__a22o_1 _3882_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][5] ),
    .A2(_0750_),
    .B1(_0752_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][5] ),
    .X(_1016_));
 sky130_fd_sc_hd__a22o_1 _3883_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ),
    .A2(_0727_),
    .B1(_0754_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ),
    .X(_1017_));
 sky130_fd_sc_hd__mux2_1 _3884_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][5] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][5] ),
    .S(_0726_),
    .X(_1018_));
 sky130_fd_sc_hd__mux2_1 _3885_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][5] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ),
    .S(_0726_),
    .X(_1019_));
 sky130_fd_sc_hd__o21a_1 _3886_ (.A1(_0721_),
    .A2(_1019_),
    .B1(_0718_),
    .X(_1020_));
 sky130_fd_sc_hd__o21ai_1 _3887_ (.A1(_0722_),
    .A2(_1018_),
    .B1(_1020_),
    .Y(_1021_));
 sky130_fd_sc_hd__or3b_4 _3888_ (.A(_1016_),
    .B(_1017_),
    .C_N(_1021_),
    .X(_1022_));
 sky130_fd_sc_hd__nand2_1 _3889_ (.A(net77),
    .B(_1022_),
    .Y(_1023_));
 sky130_fd_sc_hd__xnor2_1 _3890_ (.A(_0856_),
    .B(_1022_),
    .Y(_1024_));
 sky130_fd_sc_hd__a21o_1 _3891_ (.A1(_1001_),
    .A2(_1010_),
    .B1(_1009_),
    .X(_1025_));
 sky130_fd_sc_hd__xnor2_1 _3892_ (.A(_1024_),
    .B(_1025_),
    .Y(_1026_));
 sky130_fd_sc_hd__nor2_1 _3893_ (.A(net74),
    .B(_1026_),
    .Y(_1027_));
 sky130_fd_sc_hd__nor2_1 _3894_ (.A(_2723_),
    .B(\z80.tv80s.i_tv80_core.BusB[5] ),
    .Y(_1028_));
 sky130_fd_sc_hd__and2_1 _3895_ (.A(net108),
    .B(\z80.tv80s.i_tv80_core.BusB[5] ),
    .X(_1029_));
 sky130_fd_sc_hd__o21a_1 _3896_ (.A1(_1028_),
    .A2(_1029_),
    .B1(\z80.tv80s.i_tv80_core.BusA[5] ),
    .X(_1030_));
 sky130_fd_sc_hd__nor3_1 _3897_ (.A(\z80.tv80s.i_tv80_core.BusA[5] ),
    .B(_1028_),
    .C(_1029_),
    .Y(_1031_));
 sky130_fd_sc_hd__nor2_1 _3898_ (.A(_1030_),
    .B(_1031_),
    .Y(_1032_));
 sky130_fd_sc_hd__nand2_1 _3899_ (.A(_0985_),
    .B(_0990_),
    .Y(_1033_));
 sky130_fd_sc_hd__nand2_1 _3900_ (.A(_1032_),
    .B(_1033_),
    .Y(_1034_));
 sky130_fd_sc_hd__o21a_1 _3901_ (.A1(_1032_),
    .A2(_1033_),
    .B1(_0777_),
    .X(_1035_));
 sky130_fd_sc_hd__o21a_1 _3902_ (.A1(\z80.tv80s.i_tv80_core.ALU_Op_r[1] ),
    .A2(_1030_),
    .B1(_0764_),
    .X(_1036_));
 sky130_fd_sc_hd__a221o_1 _3903_ (.A1(_0778_),
    .A2(_1032_),
    .B1(_1034_),
    .B2(_1035_),
    .C1(_1036_),
    .X(_1037_));
 sky130_fd_sc_hd__o41a_2 _3904_ (.A1(_2723_),
    .A2(\z80.tv80s.i_tv80_core.BusA[5] ),
    .A3(\z80.tv80s.i_tv80_core.BusB[5] ),
    .A4(_0777_),
    .B1(_1037_),
    .X(_1038_));
 sky130_fd_sc_hd__and2_1 _3905_ (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .B(_0836_),
    .X(_1039_));
 sky130_fd_sc_hd__nor2_1 _3906_ (.A(\z80.tv80s.i_tv80_core.BusA[5] ),
    .B(_1039_),
    .Y(_1040_));
 sky130_fd_sc_hd__o31a_1 _3907_ (.A1(\z80.tv80s.i_tv80_core.BusA[5] ),
    .A2(\z80.tv80s.i_tv80_core.BusA[6] ),
    .A3(_1039_),
    .B1(net139),
    .X(_1041_));
 sky130_fd_sc_hd__nor2_1 _3908_ (.A(\z80.tv80s.i_tv80_core.F[0] ),
    .B(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__or2_2 _3909_ (.A(\z80.tv80s.i_tv80_core.F[0] ),
    .B(_1041_),
    .X(_1043_));
 sky130_fd_sc_hd__and3_1 _3910_ (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .B(\z80.tv80s.i_tv80_core.BusA[5] ),
    .C(_0836_),
    .X(_1044_));
 sky130_fd_sc_hd__or2_1 _3911_ (.A(_1040_),
    .B(_1044_),
    .X(_1045_));
 sky130_fd_sc_hd__or3_1 _3912_ (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .B(_0838_),
    .C(_0952_),
    .X(_1046_));
 sky130_fd_sc_hd__or2_1 _3913_ (.A(\z80.tv80s.i_tv80_core.BusA[5] ),
    .B(_1046_),
    .X(_1047_));
 sky130_fd_sc_hd__xor2_1 _3914_ (.A(\z80.tv80s.i_tv80_core.BusA[5] ),
    .B(_1046_),
    .X(_1048_));
 sky130_fd_sc_hd__mux2_1 _3915_ (.A0(_1045_),
    .A1(_1048_),
    .S(\z80.tv80s.i_tv80_core.F[1] ),
    .X(_1049_));
 sky130_fd_sc_hd__xnor2_2 _3916_ (.A(_1043_),
    .B(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__inv_2 _3917_ (.A(_1050_),
    .Y(_1051_));
 sky130_fd_sc_hd__a22o_1 _3918_ (.A1(\z80.tv80s.i_tv80_core.BusA[5] ),
    .A2(_0786_),
    .B1(_0789_),
    .B2(_1050_),
    .X(_1052_));
 sky130_fd_sc_hd__mux2_1 _3919_ (.A0(\z80.tv80s.i_tv80_core.BusA[4] ),
    .A1(\z80.tv80s.i_tv80_core.BusA[6] ),
    .S(net129),
    .X(_1053_));
 sky130_fd_sc_hd__and2_1 _3920_ (.A(_0791_),
    .B(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__nor2_1 _3921_ (.A(_0411_),
    .B(_0794_),
    .Y(_1055_));
 sky130_fd_sc_hd__a211o_1 _3922_ (.A1(_0411_),
    .A2(_0785_),
    .B1(_1055_),
    .C1(_0784_),
    .X(_1056_));
 sky130_fd_sc_hd__a221o_1 _3923_ (.A1(_0411_),
    .A2(_0784_),
    .B1(_1056_),
    .B2(\z80.tv80s.i_tv80_core.BusB[5] ),
    .C1(_1054_),
    .X(_1057_));
 sky130_fd_sc_hd__a211o_1 _3924_ (.A1(_0763_),
    .A2(_1038_),
    .B1(_1052_),
    .C1(_1057_),
    .X(_1058_));
 sky130_fd_sc_hd__mux2_1 _3925_ (.A0(\z80.tv80s.di_reg[5] ),
    .A1(_1058_),
    .S(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(_1059_));
 sky130_fd_sc_hd__mux2_4 _3926_ (.A0(_1059_),
    .A1(net605),
    .S(_0761_),
    .X(_1060_));
 sky130_fd_sc_hd__a21o_1 _3927_ (.A1(net74),
    .A2(_1060_),
    .B1(_0677_),
    .X(_1061_));
 sky130_fd_sc_hd__o22a_1 _3928_ (.A1(net234),
    .A2(net89),
    .B1(_1027_),
    .B2(_1061_),
    .X(_1062_));
 sky130_fd_sc_hd__mux4_1 _3929_ (.A0(net364),
    .A1(net315),
    .A2(net321),
    .A3(net433),
    .S0(net81),
    .S1(net82),
    .X(_1063_));
 sky130_fd_sc_hd__mux2_2 _3930_ (.A0(_1062_),
    .A1(_1063_),
    .S(net90),
    .X(_1064_));
 sky130_fd_sc_hd__mux2_1 _3931_ (.A0(net449),
    .A1(_1064_),
    .S(_0729_),
    .X(_0041_));
 sky130_fd_sc_hd__xor2_1 _3932_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[1] ),
    .B(\z80.tv80s.i_tv80_core.BusB[6] ),
    .X(_1065_));
 sky130_fd_sc_hd__and2_1 _3933_ (.A(\z80.tv80s.i_tv80_core.BusA[6] ),
    .B(_1065_),
    .X(_1066_));
 sky130_fd_sc_hd__nor2_1 _3934_ (.A(\z80.tv80s.i_tv80_core.BusA[6] ),
    .B(_1065_),
    .Y(_1067_));
 sky130_fd_sc_hd__nor2_1 _3935_ (.A(_1066_),
    .B(_1067_),
    .Y(_1068_));
 sky130_fd_sc_hd__a21o_1 _3936_ (.A1(_1032_),
    .A2(_1033_),
    .B1(_1030_),
    .X(_1069_));
 sky130_fd_sc_hd__a21oi_1 _3937_ (.A1(_1068_),
    .A2(_1069_),
    .B1(_0776_),
    .Y(_1070_));
 sky130_fd_sc_hd__o21a_1 _3938_ (.A1(_1068_),
    .A2(_1069_),
    .B1(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__or2_1 _3939_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[1] ),
    .B(_1066_),
    .X(_1072_));
 sky130_fd_sc_hd__a221o_1 _3940_ (.A1(_0778_),
    .A2(_1068_),
    .B1(_1072_),
    .B2(_0764_),
    .C1(_1071_),
    .X(_1073_));
 sky130_fd_sc_hd__o41a_2 _3941_ (.A1(net108),
    .A2(\z80.tv80s.i_tv80_core.BusA[6] ),
    .A3(\z80.tv80s.i_tv80_core.BusB[6] ),
    .A4(_0777_),
    .B1(_1073_),
    .X(_1074_));
 sky130_fd_sc_hd__xnor2_1 _3942_ (.A(\z80.tv80s.i_tv80_core.BusA[6] ),
    .B(_1044_),
    .Y(_1075_));
 sky130_fd_sc_hd__a21o_1 _3943_ (.A1(_1043_),
    .A2(_1045_),
    .B1(_1075_),
    .X(_1076_));
 sky130_fd_sc_hd__nand2_1 _3944_ (.A(_1045_),
    .B(_1075_),
    .Y(_1077_));
 sky130_fd_sc_hd__o21ai_1 _3945_ (.A1(_1042_),
    .A2(_1077_),
    .B1(_1076_),
    .Y(_1078_));
 sky130_fd_sc_hd__xor2_1 _3946_ (.A(\z80.tv80s.i_tv80_core.BusA[6] ),
    .B(_1047_),
    .X(_1079_));
 sky130_fd_sc_hd__nor2_1 _3947_ (.A(_1042_),
    .B(_1048_),
    .Y(_1080_));
 sky130_fd_sc_hd__xnor2_1 _3948_ (.A(_1079_),
    .B(_1080_),
    .Y(_1081_));
 sky130_fd_sc_hd__mux2_1 _3949_ (.A0(_1078_),
    .A1(_1081_),
    .S(\z80.tv80s.i_tv80_core.F[1] ),
    .X(_1082_));
 sky130_fd_sc_hd__nor2_1 _3950_ (.A(_2891_),
    .B(_0794_),
    .Y(_1083_));
 sky130_fd_sc_hd__mux2_1 _3951_ (.A0(\z80.tv80s.i_tv80_core.BusA[5] ),
    .A1(net139),
    .S(net129),
    .X(_1084_));
 sky130_fd_sc_hd__a221o_1 _3952_ (.A1(\z80.tv80s.i_tv80_core.BusA[6] ),
    .A2(_0786_),
    .B1(_0791_),
    .B2(_1084_),
    .C1(_0763_),
    .X(_1085_));
 sky130_fd_sc_hd__a211o_1 _3953_ (.A1(_2891_),
    .A2(_0785_),
    .B1(_1083_),
    .C1(_0784_),
    .X(_1086_));
 sky130_fd_sc_hd__a22o_1 _3954_ (.A1(_2891_),
    .A2(_0784_),
    .B1(_1086_),
    .B2(\z80.tv80s.i_tv80_core.BusB[6] ),
    .X(_1087_));
 sky130_fd_sc_hd__a211o_1 _3955_ (.A1(_0789_),
    .A2(_1082_),
    .B1(_1085_),
    .C1(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__o21ai_1 _3956_ (.A1(_0762_),
    .A2(_1074_),
    .B1(_1088_),
    .Y(_1089_));
 sky130_fd_sc_hd__mux2_1 _3957_ (.A0(_2737_),
    .A1(_1089_),
    .S(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(_1090_));
 sky130_fd_sc_hd__mux2_4 _3958_ (.A0(_1090_),
    .A1(_2729_),
    .S(_0761_),
    .X(_1091_));
 sky130_fd_sc_hd__inv_2 _3959_ (.A(_1091_),
    .Y(_1092_));
 sky130_fd_sc_hd__o21ai_2 _3960_ (.A1(_0736_),
    .A2(_1091_),
    .B1(_0678_),
    .Y(_1093_));
 sky130_fd_sc_hd__mux2_1 _3961_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][6] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][6] ),
    .S(net69),
    .X(_1094_));
 sky130_fd_sc_hd__mux2_1 _3962_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ),
    .S(net69),
    .X(_1095_));
 sky130_fd_sc_hd__mux2_1 _3963_ (.A0(_1094_),
    .A1(_1095_),
    .S(net71),
    .X(_1096_));
 sky130_fd_sc_hd__o311a_1 _3964_ (.A1(_0711_),
    .A2(net75),
    .A3(_0723_),
    .B1(_0724_),
    .C1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][6] ),
    .X(_1097_));
 sky130_fd_sc_hd__a211o_1 _3965_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][6] ),
    .A2(net70),
    .B1(_1097_),
    .C1(net71),
    .X(_1098_));
 sky130_fd_sc_hd__o311a_1 _3966_ (.A1(_0711_),
    .A2(net75),
    .A3(_0723_),
    .B1(_0724_),
    .C1(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ),
    .X(_1099_));
 sky130_fd_sc_hd__a211o_1 _3967_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][6] ),
    .A2(net70),
    .B1(_1099_),
    .C1(net72),
    .X(_1100_));
 sky130_fd_sc_hd__and3_1 _3968_ (.A(_0717_),
    .B(_1098_),
    .C(_1100_),
    .X(_1101_));
 sky130_fd_sc_hd__a21o_2 _3969_ (.A1(net65),
    .A2(_1096_),
    .B1(_1101_),
    .X(_1102_));
 sky130_fd_sc_hd__xnor2_1 _3970_ (.A(net77),
    .B(_1102_),
    .Y(_1103_));
 sky130_fd_sc_hd__o21ai_1 _3971_ (.A1(net77),
    .A2(_1022_),
    .B1(_1025_),
    .Y(_1104_));
 sky130_fd_sc_hd__o21a_1 _3972_ (.A1(_1008_),
    .A2(_1022_),
    .B1(net77),
    .X(_1105_));
 sky130_fd_sc_hd__a21oi_1 _3973_ (.A1(_1023_),
    .A2(_1104_),
    .B1(_1103_),
    .Y(_1106_));
 sky130_fd_sc_hd__and3_1 _3974_ (.A(_1023_),
    .B(_1103_),
    .C(_1104_),
    .X(_1107_));
 sky130_fd_sc_hd__or2_1 _3975_ (.A(_1106_),
    .B(_1107_),
    .X(_1108_));
 sky130_fd_sc_hd__nor2_1 _3976_ (.A(net74),
    .B(_1108_),
    .Y(_1109_));
 sky130_fd_sc_hd__o22a_1 _3977_ (.A1(net218),
    .A2(net89),
    .B1(_1093_),
    .B2(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__mux4_2 _3978_ (.A0(net477),
    .A1(net501),
    .A2(net378),
    .A3(net396),
    .S0(net81),
    .S1(net82),
    .X(_1111_));
 sky130_fd_sc_hd__mux2_2 _3979_ (.A0(_1110_),
    .A1(_1111_),
    .S(net90),
    .X(_1112_));
 sky130_fd_sc_hd__mux2_1 _3980_ (.A0(net488),
    .A1(_1112_),
    .S(_0729_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _3981_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][7] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][7] ),
    .S(net69),
    .X(_1113_));
 sky130_fd_sc_hd__mux2_1 _3982_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][7] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][7] ),
    .S(net69),
    .X(_1114_));
 sky130_fd_sc_hd__mux2_1 _3983_ (.A0(_1113_),
    .A1(_1114_),
    .S(net71),
    .X(_1115_));
 sky130_fd_sc_hd__o311a_1 _3984_ (.A1(_0711_),
    .A2(net75),
    .A3(_0723_),
    .B1(_0724_),
    .C1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][7] ),
    .X(_1116_));
 sky130_fd_sc_hd__a211o_1 _3985_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][7] ),
    .A2(net70),
    .B1(_1116_),
    .C1(net71),
    .X(_1117_));
 sky130_fd_sc_hd__o311a_1 _3986_ (.A1(_0711_),
    .A2(net75),
    .A3(_0723_),
    .B1(_0724_),
    .C1(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][7] ),
    .X(_1118_));
 sky130_fd_sc_hd__a211o_1 _3987_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ),
    .A2(net70),
    .B1(_1118_),
    .C1(net72),
    .X(_1119_));
 sky130_fd_sc_hd__and3_1 _3988_ (.A(net65),
    .B(_1117_),
    .C(_1119_),
    .X(_1120_));
 sky130_fd_sc_hd__a21o_1 _3989_ (.A1(_0717_),
    .A2(_1115_),
    .B1(_1120_),
    .X(_1121_));
 sky130_fd_sc_hd__xnor2_1 _3990_ (.A(_0856_),
    .B(_1121_),
    .Y(_1122_));
 sky130_fd_sc_hd__a21o_1 _3991_ (.A1(net77),
    .A2(_1102_),
    .B1(_1106_),
    .X(_1123_));
 sky130_fd_sc_hd__xnor2_1 _3992_ (.A(_1122_),
    .B(_1123_),
    .Y(_1124_));
 sky130_fd_sc_hd__nor2_1 _3993_ (.A(net74),
    .B(_1124_),
    .Y(_1125_));
 sky130_fd_sc_hd__a21o_1 _3994_ (.A1(_1068_),
    .A2(_1069_),
    .B1(_1066_),
    .X(_1126_));
 sky130_fd_sc_hd__xor2_1 _3995_ (.A(net139),
    .B(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__xor2_1 _3996_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[1] ),
    .B(\z80.tv80s.i_tv80_core.BusB[7] ),
    .X(_1128_));
 sky130_fd_sc_hd__or2_1 _3997_ (.A(_1127_),
    .B(_1128_),
    .X(_1129_));
 sky130_fd_sc_hd__nand2_1 _3998_ (.A(_1127_),
    .B(_1128_),
    .Y(_1130_));
 sky130_fd_sc_hd__or2_1 _3999_ (.A(net139),
    .B(\z80.tv80s.i_tv80_core.BusB[7] ),
    .X(_1131_));
 sky130_fd_sc_hd__nand2_1 _4000_ (.A(net139),
    .B(\z80.tv80s.i_tv80_core.BusB[7] ),
    .Y(_1132_));
 sky130_fd_sc_hd__nand2_1 _4001_ (.A(net108),
    .B(_1132_),
    .Y(_1133_));
 sky130_fd_sc_hd__a32o_1 _4002_ (.A1(_0778_),
    .A2(_1131_),
    .A3(_1132_),
    .B1(_1133_),
    .B2(_0764_),
    .X(_1134_));
 sky130_fd_sc_hd__a31o_1 _4003_ (.A1(_0777_),
    .A2(_1129_),
    .A3(_1130_),
    .B1(_1134_),
    .X(_1135_));
 sky130_fd_sc_hd__o41a_2 _4004_ (.A1(net108),
    .A2(net139),
    .A3(\z80.tv80s.i_tv80_core.BusB[7] ),
    .A4(_0777_),
    .B1(_1135_),
    .X(_1136_));
 sky130_fd_sc_hd__nand2_1 _4005_ (.A(_1043_),
    .B(_1077_),
    .Y(_1137_));
 sky130_fd_sc_hd__xor2_1 _4006_ (.A(net139),
    .B(\z80.tv80s.i_tv80_core.BusA[6] ),
    .X(_1138_));
 sky130_fd_sc_hd__mux2_1 _4007_ (.A0(net139),
    .A1(_1138_),
    .S(_1044_),
    .X(_1139_));
 sky130_fd_sc_hd__xnor2_1 _4008_ (.A(_1137_),
    .B(_1139_),
    .Y(_1140_));
 sky130_fd_sc_hd__or3_1 _4009_ (.A(net139),
    .B(\z80.tv80s.i_tv80_core.BusA[6] ),
    .C(_1047_),
    .X(_1141_));
 sky130_fd_sc_hd__o21ai_1 _4010_ (.A1(\z80.tv80s.i_tv80_core.BusA[6] ),
    .A2(_1047_),
    .B1(net139),
    .Y(_1142_));
 sky130_fd_sc_hd__nand2_1 _4011_ (.A(_1141_),
    .B(_1142_),
    .Y(_1143_));
 sky130_fd_sc_hd__nor2_1 _4012_ (.A(_1048_),
    .B(_1079_),
    .Y(_1144_));
 sky130_fd_sc_hd__nor2_1 _4013_ (.A(_1143_),
    .B(_1144_),
    .Y(_1145_));
 sky130_fd_sc_hd__or2_1 _4014_ (.A(_1042_),
    .B(_1144_),
    .X(_1146_));
 sky130_fd_sc_hd__a22o_1 _4015_ (.A1(_1043_),
    .A2(_1145_),
    .B1(_1146_),
    .B2(_1143_),
    .X(_1147_));
 sky130_fd_sc_hd__mux2_1 _4016_ (.A0(_1140_),
    .A1(_1147_),
    .S(\z80.tv80s.i_tv80_core.F[1] ),
    .X(_1148_));
 sky130_fd_sc_hd__and2_1 _4017_ (.A(\z80.tv80s.i_tv80_core.BusB[7] ),
    .B(_2861_),
    .X(_1149_));
 sky130_fd_sc_hd__a22o_1 _4018_ (.A1(net139),
    .A2(_0786_),
    .B1(_0789_),
    .B2(_1148_),
    .X(_1150_));
 sky130_fd_sc_hd__a31o_1 _4019_ (.A1(net625),
    .A2(_2861_),
    .A3(_0785_),
    .B1(_1150_),
    .X(_1151_));
 sky130_fd_sc_hd__nand2_1 _4020_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .B(_2861_),
    .Y(_1152_));
 sky130_fd_sc_hd__or2_1 _4021_ (.A(\z80.tv80s.i_tv80_core.BusB[7] ),
    .B(_2861_),
    .X(_1153_));
 sky130_fd_sc_hd__and2_1 _4022_ (.A(net129),
    .B(\z80.tv80s.i_tv80_core.BusA[0] ),
    .X(_1154_));
 sky130_fd_sc_hd__a22o_1 _4023_ (.A1(net119),
    .A2(\z80.tv80s.i_tv80_core.BusA[6] ),
    .B1(_2750_),
    .B2(_1154_),
    .X(_1155_));
 sky130_fd_sc_hd__a221o_2 _4024_ (.A1(net139),
    .A2(_0411_),
    .B1(_0581_),
    .B2(\z80.tv80s.i_tv80_core.F[0] ),
    .C1(_1155_),
    .X(_1156_));
 sky130_fd_sc_hd__a32o_1 _4025_ (.A1(_0783_),
    .A2(_1152_),
    .A3(_1153_),
    .B1(_1156_),
    .B2(_0791_),
    .X(_1157_));
 sky130_fd_sc_hd__a211o_1 _4026_ (.A1(_0763_),
    .A2(_1136_),
    .B1(_1151_),
    .C1(_1157_),
    .X(_1158_));
 sky130_fd_sc_hd__mux2_1 _4027_ (.A0(\z80.tv80s.di_reg[7] ),
    .A1(_1158_),
    .S(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(_1159_));
 sky130_fd_sc_hd__and2b_1 _4028_ (.A_N(_0761_),
    .B(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__a21oi_2 _4029_ (.A1(net625),
    .A2(_0761_),
    .B1(_1160_),
    .Y(_1161_));
 sky130_fd_sc_hd__inv_2 _4030_ (.A(_1161_),
    .Y(_1162_));
 sky130_fd_sc_hd__o21ai_2 _4031_ (.A1(_0736_),
    .A2(_1161_),
    .B1(_0678_),
    .Y(_1163_));
 sky130_fd_sc_hd__o22a_1 _4032_ (.A1(net220),
    .A2(net89),
    .B1(_1125_),
    .B2(_1163_),
    .X(_1164_));
 sky130_fd_sc_hd__mux4_1 _4033_ (.A0(net385),
    .A1(net275),
    .A2(net323),
    .A3(net293),
    .S0(net81),
    .S1(net82),
    .X(_1165_));
 sky130_fd_sc_hd__mux2_2 _4034_ (.A0(_1164_),
    .A1(_1165_),
    .S(net90),
    .X(_1166_));
 sky130_fd_sc_hd__mux2_1 _4035_ (.A0(net335),
    .A1(_1166_),
    .S(_0729_),
    .X(_0043_));
 sky130_fd_sc_hd__nor2_1 _4036_ (.A(net117),
    .B(_2891_),
    .Y(_1167_));
 sky130_fd_sc_hd__o31a_1 _4037_ (.A1(net95),
    .A2(_2909_),
    .A3(_1167_),
    .B1(net166),
    .X(_1168_));
 sky130_fd_sc_hd__and3_1 _4038_ (.A(net146),
    .B(_2752_),
    .C(net94),
    .X(_1169_));
 sky130_fd_sc_hd__and2_1 _4039_ (.A(_2786_),
    .B(_2812_),
    .X(_1170_));
 sky130_fd_sc_hd__or2_1 _4040_ (.A(_2817_),
    .B(_1170_),
    .X(_1171_));
 sky130_fd_sc_hd__a21oi_2 _4041_ (.A1(net94),
    .A2(_0431_),
    .B1(_2835_),
    .Y(_1172_));
 sky130_fd_sc_hd__or4_2 _4042_ (.A(net96),
    .B(_1169_),
    .C(_1171_),
    .D(_1172_),
    .X(_1173_));
 sky130_fd_sc_hd__and3_1 _4043_ (.A(_2760_),
    .B(_2773_),
    .C(_0385_),
    .X(_1174_));
 sky130_fd_sc_hd__nor2_1 _4044_ (.A(_2892_),
    .B(_0430_),
    .Y(_1175_));
 sky130_fd_sc_hd__or2_1 _4045_ (.A(_2934_),
    .B(_1175_),
    .X(_1176_));
 sky130_fd_sc_hd__nor2_1 _4046_ (.A(_2928_),
    .B(_0597_),
    .Y(_1177_));
 sky130_fd_sc_hd__a21o_1 _4047_ (.A1(_2939_),
    .A2(_1167_),
    .B1(_1177_),
    .X(_1178_));
 sky130_fd_sc_hd__or4b_1 _4048_ (.A(_1173_),
    .B(_1174_),
    .C(_1178_),
    .D_N(_1176_),
    .X(_1179_));
 sky130_fd_sc_hd__a21o_1 _4049_ (.A1(_2852_),
    .A2(_1173_),
    .B1(net125),
    .X(_1180_));
 sky130_fd_sc_hd__a32o_1 _4050_ (.A1(_1168_),
    .A2(_1179_),
    .A3(_1180_),
    .B1(net163),
    .B2(net134),
    .X(_1181_));
 sky130_fd_sc_hd__or3_2 _4051_ (.A(net151),
    .B(_2767_),
    .C(_2852_),
    .X(_1182_));
 sky130_fd_sc_hd__inv_2 _4052_ (.A(_1182_),
    .Y(_1183_));
 sky130_fd_sc_hd__and2_1 _4053_ (.A(_1167_),
    .B(_1183_),
    .X(_1184_));
 sky130_fd_sc_hd__and3_1 _4054_ (.A(net126),
    .B(_2896_),
    .C(_0589_),
    .X(_1185_));
 sky130_fd_sc_hd__a21o_1 _4055_ (.A1(_2703_),
    .A2(_1185_),
    .B1(_1184_),
    .X(_1186_));
 sky130_fd_sc_hd__nor2_2 _4056_ (.A(_2852_),
    .B(_2865_),
    .Y(_1187_));
 sky130_fd_sc_hd__o21ai_1 _4057_ (.A1(_2840_),
    .A2(_0431_),
    .B1(_0470_),
    .Y(_1188_));
 sky130_fd_sc_hd__or2_1 _4058_ (.A(_1187_),
    .B(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__a211o_1 _4059_ (.A1(net125),
    .A2(_1186_),
    .B1(_1189_),
    .C1(net105),
    .X(_1190_));
 sky130_fd_sc_hd__o21a_4 _4060_ (.A1(net107),
    .A2(_1181_),
    .B1(_1190_),
    .X(_1191_));
 sky130_fd_sc_hd__and4_1 _4061_ (.A(net122),
    .B(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ),
    .C(_2790_),
    .D(_1183_),
    .X(_1192_));
 sky130_fd_sc_hd__a2111o_1 _4062_ (.A1(_2818_),
    .A2(_1185_),
    .B1(_1192_),
    .C1(net105),
    .D1(_0618_),
    .X(_1193_));
 sky130_fd_sc_hd__o21ai_1 _4063_ (.A1(_2702_),
    .A2(net117),
    .B1(_1177_),
    .Y(_1194_));
 sky130_fd_sc_hd__a21oi_1 _4064_ (.A1(_1176_),
    .A2(_1194_),
    .B1(_2703_),
    .Y(_1195_));
 sky130_fd_sc_hd__o21a_1 _4065_ (.A1(net145),
    .A2(_0471_),
    .B1(_0419_),
    .X(_1196_));
 sky130_fd_sc_hd__a31o_1 _4066_ (.A1(net126),
    .A2(_2878_),
    .A3(_0589_),
    .B1(_1196_),
    .X(_1197_));
 sky130_fd_sc_hd__a41o_1 _4067_ (.A1(net122),
    .A2(net146),
    .A3(_2790_),
    .A4(_2939_),
    .B1(_0612_),
    .X(_1198_));
 sky130_fd_sc_hd__a311o_1 _4068_ (.A1(_2773_),
    .A2(_2818_),
    .A3(_0385_),
    .B1(_1173_),
    .C1(_1198_),
    .X(_1199_));
 sky130_fd_sc_hd__or3_1 _4069_ (.A(_1195_),
    .B(_1197_),
    .C(_1199_),
    .X(_1200_));
 sky130_fd_sc_hd__nand2_1 _4070_ (.A(net117),
    .B(net94),
    .Y(_1201_));
 sky130_fd_sc_hd__a31o_1 _4071_ (.A1(net122),
    .A2(_2790_),
    .A3(_1201_),
    .B1(_2852_),
    .X(_1202_));
 sky130_fd_sc_hd__a32o_1 _4072_ (.A1(net164),
    .A2(_1200_),
    .A3(_1202_),
    .B1(net163),
    .B2(net132),
    .X(_1203_));
 sky130_fd_sc_hd__o22a_4 _4073_ (.A1(_1188_),
    .A2(_1193_),
    .B1(_1203_),
    .B2(net107),
    .X(_1204_));
 sky130_fd_sc_hd__or4b_1 _4074_ (.A(\z80.tv80s.i_tv80_core.XY_Ind ),
    .B(_0443_),
    .C(_1191_),
    .D_N(_1204_),
    .X(_1205_));
 sky130_fd_sc_hd__mux2_1 _4075_ (.A0(\z80.tv80s.i_tv80_core.XY_State[1] ),
    .A1(\z80.tv80s.i_tv80_core.Alternate ),
    .S(_1205_),
    .X(_1206_));
 sky130_fd_sc_hd__mux2_1 _4076_ (.A0(net244),
    .A1(_1206_),
    .S(net109),
    .X(_0044_));
 sky130_fd_sc_hd__or2_2 _4077_ (.A(net142),
    .B(net163),
    .X(_1207_));
 sky130_fd_sc_hd__o21ai_1 _4078_ (.A1(net116),
    .A2(_0498_),
    .B1(_1176_),
    .Y(_1208_));
 sky130_fd_sc_hd__a22o_1 _4079_ (.A1(_2939_),
    .A2(_2940_),
    .B1(_0599_),
    .B2(net148),
    .X(_1209_));
 sky130_fd_sc_hd__a211o_1 _4080_ (.A1(_2760_),
    .A2(_0612_),
    .B1(_1208_),
    .C1(_1209_),
    .X(_1210_));
 sky130_fd_sc_hd__a22o_1 _4081_ (.A1(net145),
    .A2(_2769_),
    .B1(_0396_),
    .B2(_0398_),
    .X(_1211_));
 sky130_fd_sc_hd__a311o_1 _4082_ (.A1(net125),
    .A2(_2925_),
    .A3(_2936_),
    .B1(_1169_),
    .C1(net96),
    .X(_1212_));
 sky130_fd_sc_hd__a21o_1 _4083_ (.A1(net133),
    .A2(_1172_),
    .B1(_1212_),
    .X(_1213_));
 sky130_fd_sc_hd__or3_1 _4084_ (.A(_1210_),
    .B(_1211_),
    .C(_1213_),
    .X(_1214_));
 sky130_fd_sc_hd__or2_1 _4085_ (.A(net148),
    .B(_2892_),
    .X(_1215_));
 sky130_fd_sc_hd__a31o_1 _4086_ (.A1(net134),
    .A2(_2860_),
    .A3(_1215_),
    .B1(net95),
    .X(_1216_));
 sky130_fd_sc_hd__a21o_1 _4087_ (.A1(_0392_),
    .A2(_0590_),
    .B1(_0618_),
    .X(_1217_));
 sky130_fd_sc_hd__a22o_1 _4088_ (.A1(net148),
    .A2(_2890_),
    .B1(_1217_),
    .B2(_2703_),
    .X(_1218_));
 sky130_fd_sc_hd__a221o_1 _4089_ (.A1(_2844_),
    .A2(_2936_),
    .B1(_1218_),
    .B2(net125),
    .C1(_1189_),
    .X(_1219_));
 sky130_fd_sc_hd__a32o_1 _4090_ (.A1(net167),
    .A2(_1214_),
    .A3(_1216_),
    .B1(_1219_),
    .B2(net107),
    .X(_1220_));
 sky130_fd_sc_hd__a22o_4 _4091_ (.A1(net134),
    .A2(_1207_),
    .B1(_1220_),
    .B2(_2697_),
    .X(_1221_));
 sky130_fd_sc_hd__a31o_1 _4092_ (.A1(_2768_),
    .A2(_2936_),
    .A3(_0423_),
    .B1(_1196_),
    .X(_1222_));
 sky130_fd_sc_hd__a211o_1 _4093_ (.A1(_2818_),
    .A2(_0612_),
    .B1(_1209_),
    .C1(_1222_),
    .X(_1223_));
 sky130_fd_sc_hd__and4b_1 _4094_ (.A_N(_2774_),
    .B(net96),
    .C(_1215_),
    .D(net132),
    .X(_1224_));
 sky130_fd_sc_hd__a21o_1 _4095_ (.A1(_2702_),
    .A2(net146),
    .B1(net149),
    .X(_1225_));
 sky130_fd_sc_hd__a32o_1 _4096_ (.A1(net122),
    .A2(_2925_),
    .A3(_1225_),
    .B1(_2936_),
    .B2(_2829_),
    .X(_1226_));
 sky130_fd_sc_hd__a2111o_1 _4097_ (.A1(net131),
    .A2(_1172_),
    .B1(_1224_),
    .C1(_1226_),
    .D1(_1169_),
    .X(_1227_));
 sky130_fd_sc_hd__a211o_1 _4098_ (.A1(_0392_),
    .A2(_0593_),
    .B1(_1211_),
    .C1(_1227_),
    .X(_1228_));
 sky130_fd_sc_hd__or3_1 _4099_ (.A(_0681_),
    .B(_1223_),
    .C(_1228_),
    .X(_1229_));
 sky130_fd_sc_hd__a32o_1 _4100_ (.A1(net122),
    .A2(net148),
    .A3(_2890_),
    .B1(_0430_),
    .B2(_2844_),
    .X(_1230_));
 sky130_fd_sc_hd__a211o_1 _4101_ (.A1(_2818_),
    .A2(_1217_),
    .B1(_1230_),
    .C1(_1189_),
    .X(_1231_));
 sky130_fd_sc_hd__a22o_1 _4102_ (.A1(net167),
    .A2(_1229_),
    .B1(_1231_),
    .B2(net107),
    .X(_1232_));
 sky130_fd_sc_hd__a22o_4 _4103_ (.A1(net132),
    .A2(_1207_),
    .B1(_1232_),
    .B2(_2697_),
    .X(_1233_));
 sky130_fd_sc_hd__or4b_1 _4104_ (.A(\z80.tv80s.i_tv80_core.XY_Ind ),
    .B(_0443_),
    .C(_1221_),
    .D_N(_1233_),
    .X(_1234_));
 sky130_fd_sc_hd__mux2_1 _4105_ (.A0(net576),
    .A1(\z80.tv80s.i_tv80_core.Alternate ),
    .S(_1234_),
    .X(_1235_));
 sky130_fd_sc_hd__mux2_1 _4106_ (.A0(net584),
    .A1(_1235_),
    .S(net109),
    .X(_0045_));
 sky130_fd_sc_hd__nor2_4 _4107_ (.A(_0709_),
    .B(_0753_),
    .Y(_1236_));
 sky130_fd_sc_hd__mux2_1 _4108_ (.A0(net303),
    .A1(_0807_),
    .S(_1236_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _4109_ (.A0(net308),
    .A1(_0875_),
    .S(_1236_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _4110_ (.A0(net311),
    .A1(_0926_),
    .S(_1236_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _4111_ (.A0(net380),
    .A1(_0972_),
    .S(_1236_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _4112_ (.A0(net337),
    .A1(_1015_),
    .S(_1236_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _4113_ (.A0(net315),
    .A1(_1064_),
    .S(_1236_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _4114_ (.A0(net501),
    .A1(_1112_),
    .S(_1236_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _4115_ (.A0(net275),
    .A1(_1166_),
    .S(_1236_),
    .X(_0053_));
 sky130_fd_sc_hd__nand2_2 _4116_ (.A(net164),
    .B(_2814_),
    .Y(_1237_));
 sky130_fd_sc_hd__and3_2 _4117_ (.A(net166),
    .B(_2800_),
    .C(_2820_),
    .X(_1238_));
 sky130_fd_sc_hd__nand2_1 _4118_ (.A(net166),
    .B(_2822_),
    .Y(_1239_));
 sky130_fd_sc_hd__nand2_1 _4119_ (.A(net88),
    .B(net86),
    .Y(_1240_));
 sky130_fd_sc_hd__a21oi_1 _4120_ (.A1(net104),
    .A2(_1240_),
    .B1(net555),
    .Y(_1241_));
 sky130_fd_sc_hd__or2_1 _4121_ (.A(net555),
    .B(_1240_),
    .X(_1242_));
 sky130_fd_sc_hd__a22o_1 _4122_ (.A1(net741),
    .A2(_1241_),
    .B1(_1242_),
    .B2(net576),
    .X(_1243_));
 sky130_fd_sc_hd__mux2_1 _4123_ (.A0(net169),
    .A1(_1243_),
    .S(net109),
    .X(_0054_));
 sky130_fd_sc_hd__or4_1 _4124_ (.A(net117),
    .B(net148),
    .C(_2839_),
    .D(net106),
    .X(_1244_));
 sky130_fd_sc_hd__or3_1 _4125_ (.A(_2886_),
    .B(_0448_),
    .C(_1175_),
    .X(_1245_));
 sky130_fd_sc_hd__or3b_1 _4126_ (.A(net115),
    .B(_1245_),
    .C_N(_0634_),
    .X(_1246_));
 sky130_fd_sc_hd__a21oi_1 _4127_ (.A1(_1244_),
    .A2(_1246_),
    .B1(net155),
    .Y(_1247_));
 sky130_fd_sc_hd__a21o_1 _4128_ (.A1(net155),
    .A2(net543),
    .B1(_1247_),
    .X(_0055_));
 sky130_fd_sc_hd__nand2b_1 _4129_ (.A_N(net382),
    .B(net413),
    .Y(_1248_));
 sky130_fd_sc_hd__a2111o_1 _4130_ (.A1(\z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ),
    .A2(\z80.tv80s.i_tv80_core.Read_To_Reg_r[2] ),
    .B1(\z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ),
    .C1(_0672_),
    .D1(_1248_),
    .X(_1249_));
 sky130_fd_sc_hd__a41o_4 _4131_ (.A1(_0676_),
    .A2(_0678_),
    .A3(_0708_),
    .A4(_1249_),
    .B1(net157),
    .X(_1250_));
 sky130_fd_sc_hd__nor2_4 _4132_ (.A(_0728_),
    .B(_1250_),
    .Y(_1251_));
 sky130_fd_sc_hd__mux4_1 _4133_ (.A0(net362),
    .A1(net368),
    .A2(net456),
    .A3(net386),
    .S0(net83),
    .S1(net80),
    .X(_1252_));
 sky130_fd_sc_hd__and2b_1 _4134_ (.A_N(_1103_),
    .B(_1122_),
    .X(_1253_));
 sky130_fd_sc_hd__and4_1 _4135_ (.A(_1001_),
    .B(_1010_),
    .C(_1024_),
    .D(_1253_),
    .X(_1254_));
 sky130_fd_sc_hd__o21a_1 _4136_ (.A1(_1102_),
    .A2(_1121_),
    .B1(net77),
    .X(_1255_));
 sky130_fd_sc_hd__a211o_1 _4137_ (.A1(_1105_),
    .A2(_1253_),
    .B1(_1254_),
    .C1(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__o22a_1 _4138_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][0] ),
    .A2(_0751_),
    .B1(_0753_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][0] ),
    .X(_1257_));
 sky130_fd_sc_hd__o221a_1 _4139_ (.A1(net368),
    .A2(_0739_),
    .B1(_0741_),
    .B2(net362),
    .C1(_1257_),
    .X(_1258_));
 sky130_fd_sc_hd__o22a_1 _4140_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ),
    .A2(_0728_),
    .B1(_0743_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ),
    .X(_1259_));
 sky130_fd_sc_hd__o221a_1 _4141_ (.A1(net487),
    .A2(_0745_),
    .B1(_0755_),
    .B2(net339),
    .C1(_1259_),
    .X(_1260_));
 sky130_fd_sc_hd__nand2_2 _4142_ (.A(_1258_),
    .B(_1260_),
    .Y(_1261_));
 sky130_fd_sc_hd__inv_2 _4143_ (.A(_1261_),
    .Y(_1262_));
 sky130_fd_sc_hd__xnor2_1 _4144_ (.A(_0856_),
    .B(_1261_),
    .Y(_1263_));
 sky130_fd_sc_hd__and2b_1 _4145_ (.A_N(_1263_),
    .B(_1256_),
    .X(_1264_));
 sky130_fd_sc_hd__and2b_1 _4146_ (.A_N(_1256_),
    .B(_1263_),
    .X(_1265_));
 sky130_fd_sc_hd__or2_1 _4147_ (.A(_1264_),
    .B(_1265_),
    .X(_1266_));
 sky130_fd_sc_hd__o21ai_1 _4148_ (.A1(net74),
    .A2(_1266_),
    .B1(_0804_),
    .Y(_1267_));
 sky130_fd_sc_hd__o21a_1 _4149_ (.A1(net238),
    .A2(_0678_),
    .B1(_0676_),
    .X(_1268_));
 sky130_fd_sc_hd__a22o_2 _4150_ (.A1(net91),
    .A2(_1252_),
    .B1(_1267_),
    .B2(_1268_),
    .X(_1269_));
 sky130_fd_sc_hd__mux2_1 _4151_ (.A0(net394),
    .A1(_1269_),
    .S(_1251_),
    .X(_0056_));
 sky130_fd_sc_hd__a22o_1 _4152_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][1] ),
    .A2(_0738_),
    .B1(_0740_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][1] ),
    .X(_1270_));
 sky130_fd_sc_hd__a221o_1 _4153_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][1] ),
    .A2(_0750_),
    .B1(_0752_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][1] ),
    .C1(_1270_),
    .X(_1271_));
 sky130_fd_sc_hd__a22o_1 _4154_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ),
    .A2(_0727_),
    .B1(_0742_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ),
    .X(_1272_));
 sky130_fd_sc_hd__a221o_1 _4155_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ),
    .A2(_0744_),
    .B1(_0754_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ),
    .C1(_1272_),
    .X(_1273_));
 sky130_fd_sc_hd__nor2_2 _4156_ (.A(_1271_),
    .B(_1273_),
    .Y(_1274_));
 sky130_fd_sc_hd__inv_2 _4157_ (.A(_1274_),
    .Y(_1275_));
 sky130_fd_sc_hd__nor2_1 _4158_ (.A(_0856_),
    .B(_1274_),
    .Y(_1276_));
 sky130_fd_sc_hd__xnor2_1 _4159_ (.A(net78),
    .B(_1274_),
    .Y(_1277_));
 sky130_fd_sc_hd__a21oi_1 _4160_ (.A1(net78),
    .A2(_1262_),
    .B1(_1264_),
    .Y(_1278_));
 sky130_fd_sc_hd__xor2_1 _4161_ (.A(_1277_),
    .B(_1278_),
    .X(_1279_));
 sky130_fd_sc_hd__nor2_1 _4162_ (.A(net74),
    .B(_1279_),
    .Y(_1280_));
 sky130_fd_sc_hd__o221a_1 _4163_ (.A1(net253),
    .A2(_0678_),
    .B1(_0846_),
    .B2(_1280_),
    .C1(_0676_),
    .X(_1281_));
 sky130_fd_sc_hd__mux4_1 _4164_ (.A0(net455),
    .A1(net295),
    .A2(net418),
    .A3(net279),
    .S0(net80),
    .S1(net83),
    .X(_1282_));
 sky130_fd_sc_hd__a21o_2 _4165_ (.A1(net91),
    .A2(_1282_),
    .B1(_1281_),
    .X(_1283_));
 sky130_fd_sc_hd__mux2_1 _4166_ (.A0(net426),
    .A1(_1283_),
    .S(_1251_),
    .X(_0057_));
 sky130_fd_sc_hd__a22o_1 _4167_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][2] ),
    .A2(_0738_),
    .B1(_0740_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][2] ),
    .X(_1284_));
 sky130_fd_sc_hd__a221o_1 _4168_ (.A1(net283),
    .A2(_0750_),
    .B1(_0752_),
    .B2(net271),
    .C1(_1284_),
    .X(_1285_));
 sky130_fd_sc_hd__a22o_1 _4169_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ),
    .A2(_0727_),
    .B1(_0742_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ),
    .X(_1286_));
 sky130_fd_sc_hd__a221o_1 _4170_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ),
    .A2(_0744_),
    .B1(_0754_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ),
    .C1(_1286_),
    .X(_1287_));
 sky130_fd_sc_hd__or2_2 _4171_ (.A(_1285_),
    .B(_1287_),
    .X(_1288_));
 sky130_fd_sc_hd__nand2_1 _4172_ (.A(net78),
    .B(_1288_),
    .Y(_1289_));
 sky130_fd_sc_hd__xnor2_2 _4173_ (.A(_0856_),
    .B(_1288_),
    .Y(_1290_));
 sky130_fd_sc_hd__and2b_1 _4174_ (.A_N(_1263_),
    .B(_1277_),
    .X(_1291_));
 sky130_fd_sc_hd__a221o_1 _4175_ (.A1(net78),
    .A2(_1262_),
    .B1(_1291_),
    .B2(_1256_),
    .C1(_1276_),
    .X(_1292_));
 sky130_fd_sc_hd__xnor2_1 _4176_ (.A(_1290_),
    .B(_1292_),
    .Y(_1293_));
 sky130_fd_sc_hd__nor2_1 _4177_ (.A(net74),
    .B(_1293_),
    .Y(_1294_));
 sky130_fd_sc_hd__o221a_1 _4178_ (.A1(net232),
    .A2(net89),
    .B1(_0923_),
    .B2(_1294_),
    .C1(_0676_),
    .X(_1295_));
 sky130_fd_sc_hd__mux4_1 _4179_ (.A0(net317),
    .A1(net271),
    .A2(net403),
    .A3(net283),
    .S0(net80),
    .S1(net84),
    .X(_1296_));
 sky130_fd_sc_hd__a21o_2 _4180_ (.A1(net91),
    .A2(_1296_),
    .B1(_1295_),
    .X(_1297_));
 sky130_fd_sc_hd__mux2_1 _4181_ (.A0(net360),
    .A1(_1297_),
    .S(_1251_),
    .X(_0058_));
 sky130_fd_sc_hd__a22o_1 _4182_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][3] ),
    .A2(_0750_),
    .B1(_0752_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][3] ),
    .X(_1298_));
 sky130_fd_sc_hd__a221o_1 _4183_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][3] ),
    .A2(_0738_),
    .B1(_0740_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][3] ),
    .C1(_1298_),
    .X(_1299_));
 sky130_fd_sc_hd__a22o_1 _4184_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ),
    .A2(_0727_),
    .B1(_0742_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ),
    .X(_1300_));
 sky130_fd_sc_hd__a221o_1 _4185_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ),
    .A2(_0744_),
    .B1(_0754_),
    .B2(net390),
    .C1(_1300_),
    .X(_1301_));
 sky130_fd_sc_hd__or2_2 _4186_ (.A(_1299_),
    .B(_1301_),
    .X(_1302_));
 sky130_fd_sc_hd__xnor2_1 _4187_ (.A(_0856_),
    .B(_1302_),
    .Y(_1303_));
 sky130_fd_sc_hd__a21bo_1 _4188_ (.A1(_1290_),
    .A2(_1292_),
    .B1_N(_1289_),
    .X(_1304_));
 sky130_fd_sc_hd__xnor2_1 _4189_ (.A(_1303_),
    .B(_1304_),
    .Y(_1305_));
 sky130_fd_sc_hd__nor2_1 _4190_ (.A(net74),
    .B(_1305_),
    .Y(_1306_));
 sky130_fd_sc_hd__o22a_1 _4191_ (.A1(net226),
    .A2(net89),
    .B1(_0969_),
    .B2(_1306_),
    .X(_1307_));
 sky130_fd_sc_hd__mux4_1 _4192_ (.A0(net465),
    .A1(net376),
    .A2(net503),
    .A3(net299),
    .S0(net80),
    .S1(net84),
    .X(_1308_));
 sky130_fd_sc_hd__mux2_2 _4193_ (.A0(_1307_),
    .A1(_1308_),
    .S(net91),
    .X(_1309_));
 sky130_fd_sc_hd__mux2_1 _4194_ (.A0(net341),
    .A1(_1309_),
    .S(_1251_),
    .X(_0059_));
 sky130_fd_sc_hd__and2_1 _4195_ (.A(_1290_),
    .B(_1303_),
    .X(_1310_));
 sky130_fd_sc_hd__o41a_1 _4196_ (.A1(_1262_),
    .A2(_1275_),
    .A3(_1288_),
    .A4(_1302_),
    .B1(net78),
    .X(_1311_));
 sky130_fd_sc_hd__a31oi_2 _4197_ (.A1(_1256_),
    .A2(_1291_),
    .A3(_1310_),
    .B1(_1311_),
    .Y(_1312_));
 sky130_fd_sc_hd__a22o_1 _4198_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][4] ),
    .A2(_0738_),
    .B1(_0740_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][4] ),
    .X(_1313_));
 sky130_fd_sc_hd__a221o_1 _4199_ (.A1(net287),
    .A2(_0750_),
    .B1(_0752_),
    .B2(net285),
    .C1(_1313_),
    .X(_1314_));
 sky130_fd_sc_hd__a22o_1 _4200_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ),
    .A2(_0727_),
    .B1(_0742_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ),
    .X(_1315_));
 sky130_fd_sc_hd__a221o_1 _4201_ (.A1(net482),
    .A2(_0744_),
    .B1(_0754_),
    .B2(net423),
    .C1(_1315_),
    .X(_1316_));
 sky130_fd_sc_hd__nor2_1 _4202_ (.A(_1314_),
    .B(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__inv_2 _4203_ (.A(_1317_),
    .Y(_1318_));
 sky130_fd_sc_hd__or2_1 _4204_ (.A(_0856_),
    .B(_1317_),
    .X(_1319_));
 sky130_fd_sc_hd__nand2_1 _4205_ (.A(_0856_),
    .B(_1317_),
    .Y(_1320_));
 sky130_fd_sc_hd__nand2_1 _4206_ (.A(_1319_),
    .B(_1320_),
    .Y(_1321_));
 sky130_fd_sc_hd__xnor2_1 _4207_ (.A(_1312_),
    .B(_1321_),
    .Y(_1322_));
 sky130_fd_sc_hd__nor2_1 _4208_ (.A(net74),
    .B(_1322_),
    .Y(_1323_));
 sky130_fd_sc_hd__o22a_1 _4209_ (.A1(net246),
    .A2(net89),
    .B1(_1000_),
    .B2(_1323_),
    .X(_1324_));
 sky130_fd_sc_hd__mux4_1 _4210_ (.A0(net451),
    .A1(net285),
    .A2(net388),
    .A3(net287),
    .S0(net80),
    .S1(net83),
    .X(_1325_));
 sky130_fd_sc_hd__mux2_2 _4211_ (.A0(_1324_),
    .A1(_1325_),
    .S(net91),
    .X(_1326_));
 sky130_fd_sc_hd__mux2_1 _4212_ (.A0(net358),
    .A1(_1326_),
    .S(_1251_),
    .X(_0060_));
 sky130_fd_sc_hd__a22o_1 _4213_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][5] ),
    .A2(_0750_),
    .B1(_0752_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][5] ),
    .X(_1327_));
 sky130_fd_sc_hd__a221o_1 _4214_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][5] ),
    .A2(_0738_),
    .B1(_0740_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][5] ),
    .C1(_1327_),
    .X(_1328_));
 sky130_fd_sc_hd__a22o_1 _4215_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ),
    .A2(_0727_),
    .B1(_0742_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ),
    .X(_1329_));
 sky130_fd_sc_hd__a221o_1 _4216_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ),
    .A2(_0744_),
    .B1(_0754_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ),
    .C1(_1329_),
    .X(_1330_));
 sky130_fd_sc_hd__or2_2 _4217_ (.A(_1328_),
    .B(_1330_),
    .X(_1331_));
 sky130_fd_sc_hd__nand2_1 _4218_ (.A(net78),
    .B(_1331_),
    .Y(_1332_));
 sky130_fd_sc_hd__or2_1 _4219_ (.A(net78),
    .B(_1331_),
    .X(_1333_));
 sky130_fd_sc_hd__nand2_1 _4220_ (.A(_1332_),
    .B(_1333_),
    .Y(_1334_));
 sky130_fd_sc_hd__o21a_1 _4221_ (.A1(_1312_),
    .A2(_1321_),
    .B1(_1319_),
    .X(_1335_));
 sky130_fd_sc_hd__xnor2_1 _4222_ (.A(_1334_),
    .B(_1335_),
    .Y(_1336_));
 sky130_fd_sc_hd__nor2_1 _4223_ (.A(net74),
    .B(_1336_),
    .Y(_1337_));
 sky130_fd_sc_hd__o22a_1 _4224_ (.A1(net248),
    .A2(net89),
    .B1(_1061_),
    .B2(_1337_),
    .X(_1338_));
 sky130_fd_sc_hd__mux4_1 _4225_ (.A0(net470),
    .A1(net392),
    .A2(net445),
    .A3(net289),
    .S0(net80),
    .S1(net83),
    .X(_1339_));
 sky130_fd_sc_hd__mux2_2 _4226_ (.A0(_1338_),
    .A1(_1339_),
    .S(net91),
    .X(_1340_));
 sky130_fd_sc_hd__mux2_1 _4227_ (.A0(net354),
    .A1(_1340_),
    .S(_1251_),
    .X(_0061_));
 sky130_fd_sc_hd__a22o_1 _4228_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][6] ),
    .A2(_0738_),
    .B1(_0740_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][6] ),
    .X(_1341_));
 sky130_fd_sc_hd__a221o_1 _4229_ (.A1(net281),
    .A2(_0750_),
    .B1(_0752_),
    .B2(net297),
    .C1(_1341_),
    .X(_1342_));
 sky130_fd_sc_hd__a22o_1 _4230_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ),
    .A2(_0727_),
    .B1(_0742_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ),
    .X(_1343_));
 sky130_fd_sc_hd__a221o_1 _4231_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ),
    .A2(_0744_),
    .B1(_0754_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ),
    .C1(_1343_),
    .X(_1344_));
 sky130_fd_sc_hd__nor2_1 _4232_ (.A(_1342_),
    .B(_1344_),
    .Y(_1345_));
 sky130_fd_sc_hd__inv_2 _4233_ (.A(_1345_),
    .Y(_1346_));
 sky130_fd_sc_hd__xnor2_1 _4234_ (.A(net77),
    .B(_1345_),
    .Y(_1347_));
 sky130_fd_sc_hd__o311a_1 _4235_ (.A1(_1312_),
    .A2(_1321_),
    .A3(_1334_),
    .B1(_1332_),
    .C1(_1319_),
    .X(_1348_));
 sky130_fd_sc_hd__and2b_1 _4236_ (.A_N(_1348_),
    .B(_1347_),
    .X(_1349_));
 sky130_fd_sc_hd__and2b_1 _4237_ (.A_N(_1347_),
    .B(_1348_),
    .X(_1350_));
 sky130_fd_sc_hd__or2_1 _4238_ (.A(_1349_),
    .B(_1350_),
    .X(_1351_));
 sky130_fd_sc_hd__nor2_1 _4239_ (.A(_0737_),
    .B(_1351_),
    .Y(_1352_));
 sky130_fd_sc_hd__o22a_1 _4240_ (.A1(net222),
    .A2(net89),
    .B1(_1093_),
    .B2(_1352_),
    .X(_1353_));
 sky130_fd_sc_hd__mux4_1 _4241_ (.A0(net471),
    .A1(net297),
    .A2(net350),
    .A3(net281),
    .S0(net81),
    .S1(net84),
    .X(_1354_));
 sky130_fd_sc_hd__mux2_2 _4242_ (.A0(_1353_),
    .A1(_1354_),
    .S(net91),
    .X(_1355_));
 sky130_fd_sc_hd__mux2_1 _4243_ (.A0(net374),
    .A1(_1355_),
    .S(_1251_),
    .X(_0062_));
 sky130_fd_sc_hd__a21o_1 _4244_ (.A1(net77),
    .A2(_1346_),
    .B1(_1349_),
    .X(_1356_));
 sky130_fd_sc_hd__a22o_1 _4245_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][7] ),
    .A2(_0738_),
    .B1(_0740_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][7] ),
    .X(_1357_));
 sky130_fd_sc_hd__a221o_1 _4246_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][7] ),
    .A2(_0750_),
    .B1(_0752_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][7] ),
    .C1(_1357_),
    .X(_1358_));
 sky130_fd_sc_hd__a22o_1 _4247_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][7] ),
    .A2(_0727_),
    .B1(_0742_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][7] ),
    .X(_1359_));
 sky130_fd_sc_hd__a221o_1 _4248_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][7] ),
    .A2(_0744_),
    .B1(_0754_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][7] ),
    .C1(_1359_),
    .X(_1360_));
 sky130_fd_sc_hd__or2_1 _4249_ (.A(_1358_),
    .B(_1360_),
    .X(_1361_));
 sky130_fd_sc_hd__xnor2_1 _4250_ (.A(_0856_),
    .B(_1361_),
    .Y(_1362_));
 sky130_fd_sc_hd__xnor2_1 _4251_ (.A(_1356_),
    .B(_1362_),
    .Y(_1363_));
 sky130_fd_sc_hd__o21bai_1 _4252_ (.A1(_0737_),
    .A2(_1363_),
    .B1_N(_1163_),
    .Y(_1364_));
 sky130_fd_sc_hd__o21a_1 _4253_ (.A1(net242),
    .A2(net89),
    .B1(_0676_),
    .X(_1365_));
 sky130_fd_sc_hd__mux2_1 _4254_ (.A0(net370),
    .A1(net327),
    .S(net84),
    .X(_1366_));
 sky130_fd_sc_hd__mux2_1 _4255_ (.A0(net467),
    .A1(net431),
    .S(net84),
    .X(_1367_));
 sky130_fd_sc_hd__mux2_1 _4256_ (.A0(_1366_),
    .A1(_1367_),
    .S(net79),
    .X(_1368_));
 sky130_fd_sc_hd__o221a_1 _4257_ (.A1(net428),
    .A2(net141),
    .B1(net84),
    .B2(net459),
    .C1(net80),
    .X(_1369_));
 sky130_fd_sc_hd__o221a_1 _4258_ (.A1(net511),
    .A2(net141),
    .B1(net84),
    .B2(net495),
    .C1(net79),
    .X(_1370_));
 sky130_fd_sc_hd__or3_1 _4259_ (.A(_0809_),
    .B(_1369_),
    .C(_1370_),
    .X(_1371_));
 sky130_fd_sc_hd__o21a_1 _4260_ (.A1(_0808_),
    .A2(_1368_),
    .B1(_1371_),
    .X(_1372_));
 sky130_fd_sc_hd__a22o_2 _4261_ (.A1(_1364_),
    .A2(_1365_),
    .B1(_1372_),
    .B2(net91),
    .X(_1373_));
 sky130_fd_sc_hd__mux2_1 _4262_ (.A0(net428),
    .A1(_1373_),
    .S(_1251_),
    .X(_0063_));
 sky130_fd_sc_hd__nor2_4 _4263_ (.A(_0753_),
    .B(_1250_),
    .Y(_1374_));
 sky130_fd_sc_hd__mux2_1 _4264_ (.A0(net456),
    .A1(_1269_),
    .S(_1374_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _4265_ (.A0(net295),
    .A1(_1283_),
    .S(_1374_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _4266_ (.A0(net271),
    .A1(_1297_),
    .S(_1374_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _4267_ (.A0(net376),
    .A1(_1309_),
    .S(_1374_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _4268_ (.A0(net285),
    .A1(_1326_),
    .S(_1374_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _4269_ (.A0(net392),
    .A1(_1340_),
    .S(_1374_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _4270_ (.A0(net297),
    .A1(_1355_),
    .S(_1374_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _4271_ (.A0(net370),
    .A1(_1373_),
    .S(_1374_),
    .X(_0071_));
 sky130_fd_sc_hd__or2_1 _4272_ (.A(net109),
    .B(net162),
    .X(_1375_));
 sky130_fd_sc_hd__o31a_1 _4273_ (.A1(net155),
    .A2(_0440_),
    .A3(_1242_),
    .B1(_1375_),
    .X(_0072_));
 sky130_fd_sc_hd__nor2_4 _4274_ (.A(_0751_),
    .B(_1250_),
    .Y(_1376_));
 sky130_fd_sc_hd__mux2_1 _4275_ (.A0(net386),
    .A1(_1269_),
    .S(_1376_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _4276_ (.A0(net279),
    .A1(_1283_),
    .S(_1376_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _4277_ (.A0(net283),
    .A1(_1297_),
    .S(_1376_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _4278_ (.A0(net299),
    .A1(_1309_),
    .S(_1376_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _4279_ (.A0(net287),
    .A1(_1326_),
    .S(_1376_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _4280_ (.A0(net289),
    .A1(_1340_),
    .S(_1376_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _4281_ (.A0(net281),
    .A1(_1355_),
    .S(_1376_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _4282_ (.A0(net327),
    .A1(_1373_),
    .S(_1376_),
    .X(_0080_));
 sky130_fd_sc_hd__or2_4 _4283_ (.A(_0745_),
    .B(_1250_),
    .X(_1377_));
 sky130_fd_sc_hd__mux2_1 _4284_ (.A0(_1269_),
    .A1(net487),
    .S(_1377_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _4285_ (.A0(_1283_),
    .A1(net500),
    .S(_1377_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _4286_ (.A0(_1297_),
    .A1(net441),
    .S(_1377_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _4287_ (.A0(_1309_),
    .A1(net492),
    .S(_1377_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _4288_ (.A0(_1326_),
    .A1(net482),
    .S(_1377_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _4289_ (.A0(_1340_),
    .A1(net383),
    .S(_1377_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _4290_ (.A0(_1355_),
    .A1(net499),
    .S(_1377_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _4291_ (.A0(_1373_),
    .A1(net495),
    .S(_1377_),
    .X(_0088_));
 sky130_fd_sc_hd__or2_4 _4292_ (.A(_0709_),
    .B(_0745_),
    .X(_1378_));
 sky130_fd_sc_hd__mux2_1 _4293_ (.A0(_0807_),
    .A1(net513),
    .S(_1378_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _4294_ (.A0(_0875_),
    .A1(net538),
    .S(_1378_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _4295_ (.A0(_0926_),
    .A1(net476),
    .S(_1378_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _4296_ (.A0(_0972_),
    .A1(net356),
    .S(_1378_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _4297_ (.A0(_1015_),
    .A1(net479),
    .S(_1378_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _4298_ (.A0(_1064_),
    .A1(net404),
    .S(_1378_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _4299_ (.A0(_1112_),
    .A1(net437),
    .S(_1378_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _4300_ (.A0(_1166_),
    .A1(net458),
    .S(_1378_),
    .X(_0096_));
 sky130_fd_sc_hd__or2_4 _4301_ (.A(_0741_),
    .B(_1250_),
    .X(_1379_));
 sky130_fd_sc_hd__mux2_1 _4302_ (.A0(_1269_),
    .A1(net362),
    .S(_1379_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _4303_ (.A0(_1283_),
    .A1(net455),
    .S(_1379_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _4304_ (.A0(_1297_),
    .A1(net317),
    .S(_1379_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _4305_ (.A0(_1309_),
    .A1(net465),
    .S(_1379_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _4306_ (.A0(_1326_),
    .A1(net451),
    .S(_1379_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _4307_ (.A0(_1340_),
    .A1(net470),
    .S(_1379_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _4308_ (.A0(_1355_),
    .A1(net471),
    .S(_1379_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _4309_ (.A0(_1373_),
    .A1(net467),
    .S(_1379_),
    .X(_0104_));
 sky130_fd_sc_hd__or2_4 _4310_ (.A(_0709_),
    .B(_0739_),
    .X(_1380_));
 sky130_fd_sc_hd__mux2_1 _4311_ (.A0(_0807_),
    .A1(net434),
    .S(_1380_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _4312_ (.A0(_0875_),
    .A1(net366),
    .S(_1380_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _4313_ (.A0(_0926_),
    .A1(net345),
    .S(_1380_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _4314_ (.A0(_0972_),
    .A1(net454),
    .S(_1380_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _4315_ (.A0(_1015_),
    .A1(net422),
    .S(_1380_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _4316_ (.A0(_1064_),
    .A1(net321),
    .S(_1380_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _4317_ (.A0(_1112_),
    .A1(net378),
    .S(_1380_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _4318_ (.A0(_1166_),
    .A1(net323),
    .S(_1380_),
    .X(_0112_));
 sky130_fd_sc_hd__or2_4 _4319_ (.A(_0709_),
    .B(_0741_),
    .X(_1381_));
 sky130_fd_sc_hd__mux2_1 _4320_ (.A0(_0807_),
    .A1(net406),
    .S(_1381_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _4321_ (.A0(_0875_),
    .A1(net307),
    .S(_1381_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _4322_ (.A0(_0926_),
    .A1(net305),
    .S(_1381_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _4323_ (.A0(_0972_),
    .A1(net414),
    .S(_1381_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _4324_ (.A0(_1015_),
    .A1(net313),
    .S(_1381_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _4325_ (.A0(_1064_),
    .A1(net364),
    .S(_1381_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _4326_ (.A0(_1112_),
    .A1(net477),
    .S(_1381_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _4327_ (.A0(_1166_),
    .A1(net385),
    .S(_1381_),
    .X(_0120_));
 sky130_fd_sc_hd__or2_4 _4328_ (.A(_0709_),
    .B(_0743_),
    .X(_1382_));
 sky130_fd_sc_hd__mux2_1 _4329_ (.A0(_0807_),
    .A1(net509),
    .S(_1382_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _4330_ (.A0(_0875_),
    .A1(net522),
    .S(_1382_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _4331_ (.A0(_0926_),
    .A1(net402),
    .S(_1382_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _4332_ (.A0(_0972_),
    .A1(net411),
    .S(_1382_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _4333_ (.A0(_1015_),
    .A1(net481),
    .S(_1382_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _4334_ (.A0(_1064_),
    .A1(net319),
    .S(_1382_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _4335_ (.A0(_1112_),
    .A1(net331),
    .S(_1382_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _4336_ (.A0(_1166_),
    .A1(net480),
    .S(_1382_),
    .X(_0128_));
 sky130_fd_sc_hd__nor2_4 _4337_ (.A(_0709_),
    .B(_0755_),
    .Y(_1383_));
 sky130_fd_sc_hd__mux2_1 _4338_ (.A0(net347),
    .A1(_0807_),
    .S(_1383_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _4339_ (.A0(net425),
    .A1(_0875_),
    .S(_1383_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _4340_ (.A0(net436),
    .A1(_0926_),
    .S(_1383_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _4341_ (.A0(net325),
    .A1(_0972_),
    .S(_1383_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _4342_ (.A0(net416),
    .A1(_1015_),
    .S(_1383_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _4343_ (.A0(net352),
    .A1(_1064_),
    .S(_1383_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _4344_ (.A0(net502),
    .A1(_1112_),
    .S(_1383_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _4345_ (.A0(net444),
    .A1(_1166_),
    .S(_1383_),
    .X(_0136_));
 sky130_fd_sc_hd__or2_4 _4346_ (.A(_0743_),
    .B(_1250_),
    .X(_1384_));
 sky130_fd_sc_hd__mux2_1 _4347_ (.A0(_1269_),
    .A1(net484),
    .S(_1384_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _4348_ (.A0(_1283_),
    .A1(net494),
    .S(_1384_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _4349_ (.A0(_1297_),
    .A1(net430),
    .S(_1384_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _4350_ (.A0(_1309_),
    .A1(net506),
    .S(_1384_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _4351_ (.A0(_1326_),
    .A1(net483),
    .S(_1384_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _4352_ (.A0(_1340_),
    .A1(net447),
    .S(_1384_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _4353_ (.A0(_1355_),
    .A1(net463),
    .S(_1384_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _4354_ (.A0(_1373_),
    .A1(net511),
    .S(_1384_),
    .X(_0144_));
 sky130_fd_sc_hd__or2_4 _4355_ (.A(_0739_),
    .B(_1250_),
    .X(_1385_));
 sky130_fd_sc_hd__mux2_1 _4356_ (.A0(_1269_),
    .A1(net368),
    .S(_1385_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _4357_ (.A0(_1283_),
    .A1(net418),
    .S(_1385_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _4358_ (.A0(_1297_),
    .A1(net403),
    .S(_1385_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _4359_ (.A0(_1309_),
    .A1(net503),
    .S(_1385_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _4360_ (.A0(_1326_),
    .A1(net388),
    .S(_1385_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _4361_ (.A0(_1340_),
    .A1(net445),
    .S(_1385_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _4362_ (.A0(_1355_),
    .A1(net350),
    .S(_1385_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _4363_ (.A0(_1373_),
    .A1(net431),
    .S(_1385_),
    .X(_0152_));
 sky130_fd_sc_hd__nor2_4 _4364_ (.A(_0755_),
    .B(_1250_),
    .Y(_1386_));
 sky130_fd_sc_hd__mux2_1 _4365_ (.A0(net339),
    .A1(_1269_),
    .S(_1386_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _4366_ (.A0(net469),
    .A1(_1283_),
    .S(_1386_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _4367_ (.A0(net472),
    .A1(_1297_),
    .S(_1386_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _4368_ (.A0(net390),
    .A1(_1309_),
    .S(_1386_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _4369_ (.A0(net423),
    .A1(_1326_),
    .S(_1386_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _4370_ (.A0(net400),
    .A1(_1340_),
    .S(_1386_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _4371_ (.A0(net442),
    .A1(_1355_),
    .S(_1386_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _4372_ (.A0(net459),
    .A1(_1373_),
    .S(_1386_),
    .X(_0160_));
 sky130_fd_sc_hd__o22a_1 _4373_ (.A1(_0542_),
    .A2(_0550_),
    .B1(_0585_),
    .B2(net836),
    .X(_0161_));
 sky130_fd_sc_hd__or2_4 _4374_ (.A(net55),
    .B(net102),
    .X(_1387_));
 sky130_fd_sc_hd__inv_2 _4375_ (.A(_1387_),
    .Y(_1388_));
 sky130_fd_sc_hd__nor2_4 _4376_ (.A(net158),
    .B(_1387_),
    .Y(_1389_));
 sky130_fd_sc_hd__nor2_1 _4377_ (.A(\z80.tv80s.i_tv80_core.No_BTR ),
    .B(_0607_),
    .Y(_1390_));
 sky130_fd_sc_hd__mux2_1 _4378_ (.A0(net269),
    .A1(_1390_),
    .S(net53),
    .X(_0162_));
 sky130_fd_sc_hd__a31o_1 _4379_ (.A1(net131),
    .A2(net130),
    .A3(_2774_),
    .B1(_2800_),
    .X(_1391_));
 sky130_fd_sc_hd__a21oi_1 _4380_ (.A1(net146),
    .A2(_1391_),
    .B1(_2797_),
    .Y(_1392_));
 sky130_fd_sc_hd__nor2_1 _4381_ (.A(_2766_),
    .B(_1392_),
    .Y(_1393_));
 sky130_fd_sc_hd__a21oi_2 _4382_ (.A1(net144),
    .A2(_2805_),
    .B1(net146),
    .Y(_1394_));
 sky130_fd_sc_hd__a31oi_2 _4383_ (.A1(net125),
    .A2(net122),
    .A3(net146),
    .B1(_1394_),
    .Y(_1395_));
 sky130_fd_sc_hd__a32o_1 _4384_ (.A1(net126),
    .A2(_2878_),
    .A3(_0472_),
    .B1(_0430_),
    .B2(_2885_),
    .X(_1396_));
 sky130_fd_sc_hd__nor2_1 _4385_ (.A(_2928_),
    .B(_1394_),
    .Y(_1397_));
 sky130_fd_sc_hd__a221o_1 _4386_ (.A1(_2773_),
    .A2(_1395_),
    .B1(_1397_),
    .B2(net116),
    .C1(_1393_),
    .X(_1398_));
 sky130_fd_sc_hd__a21o_1 _4387_ (.A1(net130),
    .A2(_1201_),
    .B1(net95),
    .X(_1399_));
 sky130_fd_sc_hd__o311ai_2 _4388_ (.A1(_1173_),
    .A2(_1396_),
    .A3(_1398_),
    .B1(_1399_),
    .C1(net165),
    .Y(_1400_));
 sky130_fd_sc_hd__o211a_1 _4389_ (.A1(net118),
    .A2(_1182_),
    .B1(_0403_),
    .C1(_2857_),
    .X(_1401_));
 sky130_fd_sc_hd__nor2_1 _4390_ (.A(_2712_),
    .B(_2806_),
    .Y(_1402_));
 sky130_fd_sc_hd__nor2_1 _4391_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .B(_2805_),
    .Y(_1403_));
 sky130_fd_sc_hd__or3b_1 _4392_ (.A(_1402_),
    .B(_1403_),
    .C_N(_1185_),
    .X(_1404_));
 sky130_fd_sc_hd__o211a_1 _4393_ (.A1(net117),
    .A2(_1401_),
    .B1(_1404_),
    .C1(_0470_),
    .X(_1405_));
 sky130_fd_sc_hd__o221a_4 _4394_ (.A1(_2699_),
    .A2(_2708_),
    .B1(net105),
    .B2(_1405_),
    .C1(_1400_),
    .X(_1406_));
 sky130_fd_sc_hd__inv_2 _4395_ (.A(_1406_),
    .Y(_1407_));
 sky130_fd_sc_hd__a22o_1 _4396_ (.A1(net128),
    .A2(_2777_),
    .B1(_0396_),
    .B2(_2765_),
    .X(_1408_));
 sky130_fd_sc_hd__a31o_1 _4397_ (.A1(net128),
    .A2(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .A3(_2781_),
    .B1(_1408_),
    .X(_1409_));
 sky130_fd_sc_hd__or3_1 _4398_ (.A(net118),
    .B(net145),
    .C(_2778_),
    .X(_1410_));
 sky130_fd_sc_hd__a32o_2 _4399_ (.A1(net165),
    .A2(_1409_),
    .A3(_1410_),
    .B1(_0377_),
    .B2(_1187_),
    .X(_1411_));
 sky130_fd_sc_hd__o21a_1 _4400_ (.A1(_1407_),
    .A2(_1411_),
    .B1(_0518_),
    .X(_1412_));
 sky130_fd_sc_hd__mux2_1 _4401_ (.A0(net382),
    .A1(_1412_),
    .S(net112),
    .X(_0163_));
 sky130_fd_sc_hd__o21a_1 _4402_ (.A1(_1191_),
    .A2(_1411_),
    .B1(_0518_),
    .X(_1413_));
 sky130_fd_sc_hd__mux2_1 _4403_ (.A0(net679),
    .A1(_1413_),
    .S(net112),
    .X(_0164_));
 sky130_fd_sc_hd__o21a_1 _4404_ (.A1(_1204_),
    .A2(_1411_),
    .B1(_0518_),
    .X(_1414_));
 sky130_fd_sc_hd__mux2_1 _4405_ (.A0(net542),
    .A1(_1414_),
    .S(net112),
    .X(_0165_));
 sky130_fd_sc_hd__nor2_1 _4406_ (.A(_2806_),
    .B(_0431_),
    .Y(_1415_));
 sky130_fd_sc_hd__a32o_1 _4407_ (.A1(_2773_),
    .A2(_2805_),
    .A3(_0385_),
    .B1(_1415_),
    .B2(_2927_),
    .X(_1416_));
 sky130_fd_sc_hd__a21o_1 _4408_ (.A1(_2805_),
    .A2(_1185_),
    .B1(_1187_),
    .X(_1417_));
 sky130_fd_sc_hd__a22o_2 _4409_ (.A1(net164),
    .A2(_1416_),
    .B1(_1417_),
    .B2(net107),
    .X(_1418_));
 sky130_fd_sc_hd__nor2_1 _4410_ (.A(net158),
    .B(_1411_),
    .Y(_1419_));
 sky130_fd_sc_hd__a32o_1 _4411_ (.A1(_0518_),
    .A2(_1418_),
    .A3(_1419_),
    .B1(net635),
    .B2(net158),
    .X(_0166_));
 sky130_fd_sc_hd__nor2_1 _4412_ (.A(_2835_),
    .B(_2859_),
    .Y(_1420_));
 sky130_fd_sc_hd__or4_1 _4413_ (.A(_2833_),
    .B(_2867_),
    .C(_2887_),
    .D(_1420_),
    .X(_1421_));
 sky130_fd_sc_hd__a22o_1 _4414_ (.A1(_2868_),
    .A2(_2869_),
    .B1(_1421_),
    .B2(net150),
    .X(_1422_));
 sky130_fd_sc_hd__and2_1 _4415_ (.A(net163),
    .B(_1422_),
    .X(_1423_));
 sky130_fd_sc_hd__or3_1 _4416_ (.A(_1169_),
    .B(_1171_),
    .C(_1208_),
    .X(_1424_));
 sky130_fd_sc_hd__or3_1 _4417_ (.A(_2766_),
    .B(_2771_),
    .C(_0384_),
    .X(_1425_));
 sky130_fd_sc_hd__or4b_1 _4418_ (.A(_2851_),
    .B(_1172_),
    .C(_1178_),
    .D_N(_1425_),
    .X(_1426_));
 sky130_fd_sc_hd__o31a_1 _4419_ (.A1(_1197_),
    .A2(_1424_),
    .A3(_1426_),
    .B1(_1168_),
    .X(_1427_));
 sky130_fd_sc_hd__a221o_1 _4420_ (.A1(net148),
    .A2(_2844_),
    .B1(_0379_),
    .B2(_0396_),
    .C1(_0618_),
    .X(_1428_));
 sky130_fd_sc_hd__o31a_1 _4421_ (.A1(_1184_),
    .A2(_1185_),
    .A3(_1428_),
    .B1(net107),
    .X(_1429_));
 sky130_fd_sc_hd__o41a_1 _4422_ (.A1(_1411_),
    .A2(_1423_),
    .A3(_1427_),
    .A4(_1429_),
    .B1(_0518_),
    .X(_1430_));
 sky130_fd_sc_hd__mux2_1 _4423_ (.A0(net413),
    .A1(_1430_),
    .S(net112),
    .X(_0167_));
 sky130_fd_sc_hd__or4_1 _4424_ (.A(_2773_),
    .B(_2823_),
    .C(_2831_),
    .D(_0447_),
    .X(_1431_));
 sky130_fd_sc_hd__a211o_1 _4425_ (.A1(_2787_),
    .A2(_2812_),
    .B1(_2913_),
    .C1(_2943_),
    .X(_1432_));
 sky130_fd_sc_hd__or4_1 _4426_ (.A(_2770_),
    .B(_2815_),
    .C(_0448_),
    .D(_0628_),
    .X(_1433_));
 sky130_fd_sc_hd__or4_1 _4427_ (.A(_2931_),
    .B(_0495_),
    .C(_1432_),
    .D(_1433_),
    .X(_1434_));
 sky130_fd_sc_hd__or3_1 _4428_ (.A(_2878_),
    .B(_2886_),
    .C(_0625_),
    .X(_1435_));
 sky130_fd_sc_hd__or3_1 _4429_ (.A(_1431_),
    .B(_1434_),
    .C(_1435_),
    .X(_1436_));
 sky130_fd_sc_hd__a221o_1 _4430_ (.A1(_2920_),
    .A2(_0384_),
    .B1(_0431_),
    .B2(_2789_),
    .C1(_1436_),
    .X(_1437_));
 sky130_fd_sc_hd__a21o_1 _4431_ (.A1(net94),
    .A2(_0480_),
    .B1(_0481_),
    .X(_1438_));
 sky130_fd_sc_hd__o211a_1 _4432_ (.A1(net95),
    .A2(_2865_),
    .B1(_0380_),
    .C1(_2857_),
    .X(_1439_));
 sky130_fd_sc_hd__or4_1 _4433_ (.A(_2845_),
    .B(_2856_),
    .C(_0379_),
    .D(_1187_),
    .X(_1440_));
 sky130_fd_sc_hd__o221a_1 _4434_ (.A1(net150),
    .A2(_2843_),
    .B1(_2857_),
    .B2(_0385_),
    .C1(_1440_),
    .X(_1441_));
 sky130_fd_sc_hd__nor2_1 _4435_ (.A(net106),
    .B(_1441_),
    .Y(_1442_));
 sky130_fd_sc_hd__a221o_1 _4436_ (.A1(net166),
    .A2(_1437_),
    .B1(_1438_),
    .B2(net163),
    .C1(_1442_),
    .X(_1443_));
 sky130_fd_sc_hd__a22o_1 _4437_ (.A1(_0377_),
    .A2(_0435_),
    .B1(_1170_),
    .B2(net165),
    .X(_1444_));
 sky130_fd_sc_hd__a21o_1 _4438_ (.A1(net121),
    .A2(_1443_),
    .B1(_1444_),
    .X(_1445_));
 sky130_fd_sc_hd__or2_1 _4439_ (.A(_2916_),
    .B(_2939_),
    .X(_1446_));
 sky130_fd_sc_hd__a221o_1 _4440_ (.A1(_2834_),
    .A2(net94),
    .B1(_0480_),
    .B2(_1446_),
    .C1(_0577_),
    .X(_1447_));
 sky130_fd_sc_hd__a21bo_1 _4441_ (.A1(net119),
    .A2(_0480_),
    .B1_N(_1447_),
    .X(_1448_));
 sky130_fd_sc_hd__a311o_1 _4442_ (.A1(net150),
    .A2(_2835_),
    .A3(_2852_),
    .B1(_2859_),
    .C1(_0853_),
    .X(_1449_));
 sky130_fd_sc_hd__a21oi_1 _4443_ (.A1(_1448_),
    .A2(_1449_),
    .B1(_2708_),
    .Y(_1450_));
 sky130_fd_sc_hd__o31a_1 _4444_ (.A1(_2856_),
    .A2(_0379_),
    .A3(_1439_),
    .B1(net126),
    .X(_1451_));
 sky130_fd_sc_hd__nor2_1 _4445_ (.A(net126),
    .B(_2857_),
    .Y(_1452_));
 sky130_fd_sc_hd__nor2_1 _4446_ (.A(_2839_),
    .B(_0431_),
    .Y(_1453_));
 sky130_fd_sc_hd__a2111o_1 _4447_ (.A1(net116),
    .A2(_2844_),
    .B1(_0434_),
    .C1(_1451_),
    .D1(_1452_),
    .X(_1454_));
 sky130_fd_sc_hd__o311a_1 _4448_ (.A1(net126),
    .A2(_0618_),
    .A3(_1453_),
    .B1(_1454_),
    .C1(net107),
    .X(_1455_));
 sky130_fd_sc_hd__a22o_1 _4449_ (.A1(net117),
    .A2(_2920_),
    .B1(_1436_),
    .B2(net128),
    .X(_1456_));
 sky130_fd_sc_hd__a211o_1 _4450_ (.A1(net166),
    .A2(_1456_),
    .B1(_1455_),
    .C1(_1450_),
    .X(_1457_));
 sky130_fd_sc_hd__and4bb_1 _4451_ (.A_N(net155),
    .B_N(_1445_),
    .C(net144),
    .D(\z80.tv80s.i_tv80_core.ISet[1] ),
    .X(_1458_));
 sky130_fd_sc_hd__a22o_1 _4452_ (.A1(net160),
    .A2(net409),
    .B1(_1457_),
    .B2(_1458_),
    .X(_0168_));
 sky130_fd_sc_hd__a22o_1 _4453_ (.A1(net155),
    .A2(net711),
    .B1(_0563_),
    .B2(_0612_),
    .X(_0169_));
 sky130_fd_sc_hd__a22o_1 _4454_ (.A1(\z80.tv80s.i_tv80_core.NMICycle ),
    .A2(_0650_),
    .B1(_0654_),
    .B2(net504),
    .X(_0170_));
 sky130_fd_sc_hd__o21a_1 _4455_ (.A1(net155),
    .A2(_0520_),
    .B1(net749),
    .X(_0171_));
 sky130_fd_sc_hd__a21bo_1 _4456_ (.A1(net746),
    .A2(_0650_),
    .B1_N(_0661_),
    .X(_0172_));
 sky130_fd_sc_hd__or2_1 _4457_ (.A(_0543_),
    .B(_0550_),
    .X(_1459_));
 sky130_fd_sc_hd__a32o_1 _4458_ (.A1(_2703_),
    .A2(_0548_),
    .A3(_0549_),
    .B1(_1459_),
    .B2(net507),
    .X(_0173_));
 sky130_fd_sc_hd__a32o_1 _4459_ (.A1(_2805_),
    .A2(_0548_),
    .A3(_0549_),
    .B1(_1459_),
    .B2(net576),
    .X(_0174_));
 sky130_fd_sc_hd__and4_1 _4460_ (.A(net164),
    .B(net110),
    .C(_2884_),
    .D(net101),
    .X(_1460_));
 sky130_fd_sc_hd__xnor2_1 _4461_ (.A(_2718_),
    .B(_1460_),
    .Y(_0175_));
 sky130_fd_sc_hd__a2111o_1 _4462_ (.A1(net116),
    .A2(_2931_),
    .B1(_2943_),
    .C1(_0420_),
    .D1(_2914_),
    .X(_1461_));
 sky130_fd_sc_hd__a22o_1 _4463_ (.A1(_0473_),
    .A2(_0556_),
    .B1(_1461_),
    .B2(net145),
    .X(_1462_));
 sky130_fd_sc_hd__o21ai_1 _4464_ (.A1(net149),
    .A2(_2895_),
    .B1(_2897_),
    .Y(_1463_));
 sky130_fd_sc_hd__a32o_2 _4465_ (.A1(net145),
    .A2(net107),
    .A3(_1463_),
    .B1(_1462_),
    .B2(net164),
    .X(_1464_));
 sky130_fd_sc_hd__nand2_4 _4466_ (.A(net136),
    .B(_1464_),
    .Y(_1465_));
 sky130_fd_sc_hd__mux4_1 _4467_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ),
    .S0(net162),
    .S1(net153),
    .X(_1466_));
 sky130_fd_sc_hd__mux4_1 _4468_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][0] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ),
    .S0(net162),
    .S1(net153),
    .X(_1467_));
 sky130_fd_sc_hd__mux2_4 _4469_ (.A0(_1467_),
    .A1(_1466_),
    .S(net169),
    .X(_1468_));
 sky130_fd_sc_hd__and2b_1 _4470_ (.A_N(net137),
    .B(\z80.tv80s.i_tv80_core.SP[0] ),
    .X(_1469_));
 sky130_fd_sc_hd__a31o_1 _4471_ (.A1(net137),
    .A2(\z80.tv80s.di_reg[0] ),
    .A3(_1468_),
    .B1(_1469_),
    .X(_1470_));
 sky130_fd_sc_hd__nor2_1 _4472_ (.A(\z80.tv80s.di_reg[0] ),
    .B(_1468_),
    .Y(_1471_));
 sky130_fd_sc_hd__a21oi_1 _4473_ (.A1(net137),
    .A2(_1471_),
    .B1(_1470_),
    .Y(_1472_));
 sky130_fd_sc_hd__and2_4 _4474_ (.A(net555),
    .B(net136),
    .X(_1473_));
 sky130_fd_sc_hd__nand2_2 _4475_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ),
    .B(net136),
    .Y(_1474_));
 sky130_fd_sc_hd__nor2_1 _4476_ (.A(net103),
    .B(_1474_),
    .Y(_1475_));
 sky130_fd_sc_hd__a211o_1 _4477_ (.A1(net746),
    .A2(net517),
    .B1(net619),
    .C1(net519),
    .X(_1476_));
 sky130_fd_sc_hd__nand2_1 _4478_ (.A(net746),
    .B(net263),
    .Y(_1477_));
 sky130_fd_sc_hd__and3_4 _4479_ (.A(_0545_),
    .B(_1476_),
    .C(_1477_),
    .X(_1478_));
 sky130_fd_sc_hd__mux2_1 _4480_ (.A0(net744),
    .A1(net1),
    .S(_1478_),
    .X(_1479_));
 sky130_fd_sc_hd__a22o_1 _4481_ (.A1(_1472_),
    .A2(_1475_),
    .B1(_1479_),
    .B2(net103),
    .X(_1480_));
 sky130_fd_sc_hd__mux2_1 _4482_ (.A0(\z80.tv80s.di_reg[0] ),
    .A1(_1480_),
    .S(_1465_),
    .X(_1481_));
 sky130_fd_sc_hd__or3_1 _4483_ (.A(_2933_),
    .B(_0448_),
    .C(_0632_),
    .X(_1482_));
 sky130_fd_sc_hd__or3_2 _4484_ (.A(_2943_),
    .B(_0627_),
    .C(_1482_),
    .X(_1483_));
 sky130_fd_sc_hd__nand2_1 _4485_ (.A(net131),
    .B(net165),
    .Y(_1484_));
 sky130_fd_sc_hd__or4_1 _4486_ (.A(_2753_),
    .B(_2828_),
    .C(_0587_),
    .D(_1484_),
    .X(_1485_));
 sky130_fd_sc_hd__nor3_2 _4487_ (.A(_1435_),
    .B(_1483_),
    .C(_1485_),
    .Y(_1486_));
 sky130_fd_sc_hd__nand2_2 _4488_ (.A(_0545_),
    .B(_1486_),
    .Y(_1487_));
 sky130_fd_sc_hd__and2_4 _4489_ (.A(_1474_),
    .B(_1487_),
    .X(_1488_));
 sky130_fd_sc_hd__a31o_1 _4490_ (.A1(net101),
    .A2(_1465_),
    .A3(_1488_),
    .B1(net157),
    .X(_1489_));
 sky130_fd_sc_hd__a22o_1 _4491_ (.A1(net109),
    .A2(_1481_),
    .B1(_1489_),
    .B2(net744),
    .X(_0176_));
 sky130_fd_sc_hd__a311o_4 _4492_ (.A1(net107),
    .A2(_0852_),
    .A3(_0854_),
    .B1(_0850_),
    .C1(net136),
    .X(_1490_));
 sky130_fd_sc_hd__nand2_1 _4493_ (.A(net137),
    .B(_2732_),
    .Y(_1491_));
 sky130_fd_sc_hd__mux4_1 _4494_ (.A0(net349),
    .A1(net408),
    .A2(net308),
    .A3(net425),
    .S0(net162),
    .S1(net153),
    .X(_1492_));
 sky130_fd_sc_hd__mux4_1 _4495_ (.A0(net366),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ),
    .A2(net307),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ),
    .S0(net162),
    .S1(net153),
    .X(_1493_));
 sky130_fd_sc_hd__mux2_2 _4496_ (.A0(_1493_),
    .A1(_1492_),
    .S(net169),
    .X(_1494_));
 sky130_fd_sc_hd__mux2_1 _4497_ (.A0(\z80.tv80s.i_tv80_core.SP[1] ),
    .A1(_1494_),
    .S(net136),
    .X(_1495_));
 sky130_fd_sc_hd__and3_1 _4498_ (.A(_1490_),
    .B(_1491_),
    .C(_1495_),
    .X(_1496_));
 sky130_fd_sc_hd__a21o_1 _4499_ (.A1(_1490_),
    .A2(_1491_),
    .B1(_1495_),
    .X(_1497_));
 sky130_fd_sc_hd__and2b_1 _4500_ (.A_N(_1496_),
    .B(_1497_),
    .X(_1498_));
 sky130_fd_sc_hd__xor2_1 _4501_ (.A(_1470_),
    .B(_1498_),
    .X(_1499_));
 sky130_fd_sc_hd__a22o_1 _4502_ (.A1(net765),
    .A2(_1488_),
    .B1(_1499_),
    .B2(_1473_),
    .X(_1500_));
 sky130_fd_sc_hd__mux2_1 _4503_ (.A0(net765),
    .A1(net2),
    .S(_1478_),
    .X(_1501_));
 sky130_fd_sc_hd__mux2_1 _4504_ (.A0(_1500_),
    .A1(_1501_),
    .S(net103),
    .X(_1502_));
 sky130_fd_sc_hd__mux2_1 _4505_ (.A0(\z80.tv80s.di_reg[1] ),
    .A1(_1502_),
    .S(_1465_),
    .X(_1503_));
 sky130_fd_sc_hd__mux2_1 _4506_ (.A0(net765),
    .A1(_1503_),
    .S(net109),
    .X(_0177_));
 sky130_fd_sc_hd__nand2_1 _4507_ (.A(net137),
    .B(_2735_),
    .Y(_1504_));
 sky130_fd_sc_hd__mux4_1 _4508_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ),
    .S0(net153),
    .S1(net162),
    .X(_1505_));
 sky130_fd_sc_hd__mux4_1 _4509_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ),
    .S0(net153),
    .S1(net162),
    .X(_1506_));
 sky130_fd_sc_hd__mux2_2 _4510_ (.A0(_1506_),
    .A1(_1505_),
    .S(net169),
    .X(_1507_));
 sky130_fd_sc_hd__mux2_1 _4511_ (.A0(\z80.tv80s.i_tv80_core.SP[2] ),
    .A1(_1507_),
    .S(net137),
    .X(_1508_));
 sky130_fd_sc_hd__and3_1 _4512_ (.A(_1490_),
    .B(_1504_),
    .C(_1508_),
    .X(_1509_));
 sky130_fd_sc_hd__a21o_1 _4513_ (.A1(_1490_),
    .A2(_1504_),
    .B1(_1508_),
    .X(_1510_));
 sky130_fd_sc_hd__nand2b_1 _4514_ (.A_N(_1509_),
    .B(_1510_),
    .Y(_1511_));
 sky130_fd_sc_hd__a21o_1 _4515_ (.A1(_1470_),
    .A2(_1497_),
    .B1(_1496_),
    .X(_1512_));
 sky130_fd_sc_hd__xnor2_1 _4516_ (.A(_1511_),
    .B(_1512_),
    .Y(_1513_));
 sky130_fd_sc_hd__a22o_1 _4517_ (.A1(net759),
    .A2(_1488_),
    .B1(_1513_),
    .B2(_1473_),
    .X(_1514_));
 sky130_fd_sc_hd__mux2_1 _4518_ (.A0(net759),
    .A1(net3),
    .S(_1478_),
    .X(_1515_));
 sky130_fd_sc_hd__mux2_1 _4519_ (.A0(_1514_),
    .A1(_1515_),
    .S(net103),
    .X(_1516_));
 sky130_fd_sc_hd__mux2_1 _4520_ (.A0(\z80.tv80s.di_reg[2] ),
    .A1(_1516_),
    .S(_1465_),
    .X(_1517_));
 sky130_fd_sc_hd__mux2_1 _4521_ (.A0(net759),
    .A1(_1517_),
    .S(net109),
    .X(_0178_));
 sky130_fd_sc_hd__nand2_1 _4522_ (.A(net137),
    .B(_2734_),
    .Y(_1518_));
 sky130_fd_sc_hd__mux4_1 _4523_ (.A0(net329),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][3] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][3] ),
    .S0(net153),
    .S1(net162),
    .X(_1519_));
 sky130_fd_sc_hd__mux4_1 _4524_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][3] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][3] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ),
    .S0(net153),
    .S1(net162),
    .X(_1520_));
 sky130_fd_sc_hd__mux2_2 _4525_ (.A0(_1520_),
    .A1(_1519_),
    .S(net169),
    .X(_1521_));
 sky130_fd_sc_hd__mux2_1 _4526_ (.A0(\z80.tv80s.i_tv80_core.SP[3] ),
    .A1(_1521_),
    .S(net137),
    .X(_1522_));
 sky130_fd_sc_hd__nand3_1 _4527_ (.A(_1490_),
    .B(_1518_),
    .C(_1522_),
    .Y(_1523_));
 sky130_fd_sc_hd__a21o_1 _4528_ (.A1(_1490_),
    .A2(_1518_),
    .B1(_1522_),
    .X(_1524_));
 sky130_fd_sc_hd__nand2_1 _4529_ (.A(_1523_),
    .B(_1524_),
    .Y(_1525_));
 sky130_fd_sc_hd__a21o_1 _4530_ (.A1(_1510_),
    .A2(_1512_),
    .B1(_1509_),
    .X(_1526_));
 sky130_fd_sc_hd__xnor2_1 _4531_ (.A(_1525_),
    .B(_1526_),
    .Y(_1527_));
 sky130_fd_sc_hd__mux2_1 _4532_ (.A0(net129),
    .A1(net757),
    .S(_1487_),
    .X(_1528_));
 sky130_fd_sc_hd__mux2_1 _4533_ (.A0(_1527_),
    .A1(_1528_),
    .S(_1474_),
    .X(_1529_));
 sky130_fd_sc_hd__mux2_1 _4534_ (.A0(net757),
    .A1(net4),
    .S(_1478_),
    .X(_1530_));
 sky130_fd_sc_hd__mux2_1 _4535_ (.A0(_1529_),
    .A1(_1530_),
    .S(net103),
    .X(_1531_));
 sky130_fd_sc_hd__mux2_1 _4536_ (.A0(\z80.tv80s.di_reg[3] ),
    .A1(_1531_),
    .S(_1465_),
    .X(_1532_));
 sky130_fd_sc_hd__mux2_1 _4537_ (.A0(net757),
    .A1(_1532_),
    .S(net112),
    .X(_0179_));
 sky130_fd_sc_hd__nand2_1 _4538_ (.A(net137),
    .B(_2736_),
    .Y(_1533_));
 sky130_fd_sc_hd__mux4_1 _4539_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][4] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][4] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ),
    .S0(net153),
    .S1(net162),
    .X(_1534_));
 sky130_fd_sc_hd__mux4_1 _4540_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][4] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][4] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ),
    .S0(net152),
    .S1(net161),
    .X(_1535_));
 sky130_fd_sc_hd__mux2_2 _4541_ (.A0(_1535_),
    .A1(_1534_),
    .S(net169),
    .X(_1536_));
 sky130_fd_sc_hd__mux2_1 _4542_ (.A0(\z80.tv80s.i_tv80_core.SP[4] ),
    .A1(_1536_),
    .S(net137),
    .X(_1537_));
 sky130_fd_sc_hd__nand3_1 _4543_ (.A(_1490_),
    .B(_1533_),
    .C(_1537_),
    .Y(_1538_));
 sky130_fd_sc_hd__a21o_1 _4544_ (.A1(_1490_),
    .A2(_1533_),
    .B1(_1537_),
    .X(_1539_));
 sky130_fd_sc_hd__nand2_1 _4545_ (.A(_1538_),
    .B(_1539_),
    .Y(_1540_));
 sky130_fd_sc_hd__a21bo_1 _4546_ (.A1(_1524_),
    .A2(_1526_),
    .B1_N(_1523_),
    .X(_1541_));
 sky130_fd_sc_hd__xnor2_2 _4547_ (.A(_1540_),
    .B(_1541_),
    .Y(_1542_));
 sky130_fd_sc_hd__mux2_1 _4548_ (.A0(net125),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .S(_1487_),
    .X(_1543_));
 sky130_fd_sc_hd__mux2_1 _4549_ (.A0(_1542_),
    .A1(_1543_),
    .S(_1474_),
    .X(_1544_));
 sky130_fd_sc_hd__mux2_1 _4550_ (.A0(net763),
    .A1(net5),
    .S(_1478_),
    .X(_1545_));
 sky130_fd_sc_hd__mux2_1 _4551_ (.A0(_1544_),
    .A1(_1545_),
    .S(net103),
    .X(_1546_));
 sky130_fd_sc_hd__mux2_1 _4552_ (.A0(\z80.tv80s.di_reg[4] ),
    .A1(_1546_),
    .S(_1465_),
    .X(_1547_));
 sky130_fd_sc_hd__mux2_1 _4553_ (.A0(net763),
    .A1(_1547_),
    .S(net112),
    .X(_0180_));
 sky130_fd_sc_hd__nand2b_1 _4554_ (.A_N(\z80.tv80s.di_reg[5] ),
    .B(net137),
    .Y(_1548_));
 sky130_fd_sc_hd__mux4_1 _4555_ (.A0(net433),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][5] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ),
    .S0(net153),
    .S1(net162),
    .X(_1549_));
 sky130_fd_sc_hd__mux4_1 _4556_ (.A0(net321),
    .A1(net364),
    .A2(net319),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ),
    .S0(net153),
    .S1(net162),
    .X(_1550_));
 sky130_fd_sc_hd__mux2_2 _4557_ (.A0(_1550_),
    .A1(_1549_),
    .S(net169),
    .X(_1551_));
 sky130_fd_sc_hd__mux2_1 _4558_ (.A0(\z80.tv80s.i_tv80_core.SP[5] ),
    .A1(_1551_),
    .S(net137),
    .X(_1552_));
 sky130_fd_sc_hd__nand3_1 _4559_ (.A(_1490_),
    .B(_1548_),
    .C(_1552_),
    .Y(_1553_));
 sky130_fd_sc_hd__a21o_1 _4560_ (.A1(_1490_),
    .A2(_1548_),
    .B1(_1552_),
    .X(_1554_));
 sky130_fd_sc_hd__nand2_1 _4561_ (.A(_1553_),
    .B(_1554_),
    .Y(_1555_));
 sky130_fd_sc_hd__a21bo_1 _4562_ (.A1(_1539_),
    .A2(_1541_),
    .B1_N(_1538_),
    .X(_1556_));
 sky130_fd_sc_hd__xnor2_1 _4563_ (.A(_1555_),
    .B(_1556_),
    .Y(_1557_));
 sky130_fd_sc_hd__mux2_1 _4564_ (.A0(net122),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .S(_1487_),
    .X(_1558_));
 sky130_fd_sc_hd__mux2_1 _4565_ (.A0(_1557_),
    .A1(_1558_),
    .S(_1474_),
    .X(_1559_));
 sky130_fd_sc_hd__mux2_1 _4566_ (.A0(net776),
    .A1(net6),
    .S(_1478_),
    .X(_1560_));
 sky130_fd_sc_hd__mux2_1 _4567_ (.A0(_1559_),
    .A1(_1560_),
    .S(net103),
    .X(_1561_));
 sky130_fd_sc_hd__mux2_1 _4568_ (.A0(\z80.tv80s.di_reg[5] ),
    .A1(_1561_),
    .S(_1465_),
    .X(_1562_));
 sky130_fd_sc_hd__mux2_1 _4569_ (.A0(net776),
    .A1(_1562_),
    .S(net112),
    .X(_0181_));
 sky130_fd_sc_hd__nand2_1 _4570_ (.A(net137),
    .B(_2737_),
    .Y(_1563_));
 sky130_fd_sc_hd__mux4_1 _4571_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][6] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][6] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][6] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ),
    .S0(net153),
    .S1(net162),
    .X(_1564_));
 sky130_fd_sc_hd__mux4_1 _4572_ (.A0(net378),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][6] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ),
    .S0(net153),
    .S1(net162),
    .X(_1565_));
 sky130_fd_sc_hd__mux2_2 _4573_ (.A0(_1565_),
    .A1(_1564_),
    .S(net169),
    .X(_1566_));
 sky130_fd_sc_hd__mux2_1 _4574_ (.A0(\z80.tv80s.i_tv80_core.SP[6] ),
    .A1(_1566_),
    .S(net137),
    .X(_1567_));
 sky130_fd_sc_hd__and3_1 _4575_ (.A(_1490_),
    .B(_1563_),
    .C(_1567_),
    .X(_1568_));
 sky130_fd_sc_hd__a21o_1 _4576_ (.A1(_1490_),
    .A2(_1563_),
    .B1(_1567_),
    .X(_1569_));
 sky130_fd_sc_hd__nand2b_1 _4577_ (.A_N(_1568_),
    .B(_1569_),
    .Y(_1570_));
 sky130_fd_sc_hd__a21bo_1 _4578_ (.A1(_1554_),
    .A2(_1556_),
    .B1_N(_1553_),
    .X(_1571_));
 sky130_fd_sc_hd__xnor2_1 _4579_ (.A(_1570_),
    .B(_1571_),
    .Y(_1572_));
 sky130_fd_sc_hd__a22o_1 _4580_ (.A1(net769),
    .A2(_1488_),
    .B1(_1572_),
    .B2(_1473_),
    .X(_1573_));
 sky130_fd_sc_hd__mux2_1 _4581_ (.A0(net769),
    .A1(net7),
    .S(_1478_),
    .X(_1574_));
 sky130_fd_sc_hd__mux2_1 _4582_ (.A0(_1573_),
    .A1(_1574_),
    .S(net102),
    .X(_1575_));
 sky130_fd_sc_hd__mux2_1 _4583_ (.A0(\z80.tv80s.di_reg[6] ),
    .A1(_1575_),
    .S(_1465_),
    .X(_1576_));
 sky130_fd_sc_hd__mux2_1 _4584_ (.A0(net769),
    .A1(_1576_),
    .S(net112),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_2 _4585_ (.A0(net78),
    .A1(\z80.tv80s.di_reg[7] ),
    .S(net137),
    .X(_1577_));
 sky130_fd_sc_hd__mux4_1 _4586_ (.A0(net293),
    .A1(net275),
    .A2(net335),
    .A3(net444),
    .S0(net153),
    .S1(net162),
    .X(_1578_));
 sky130_fd_sc_hd__mux4_1 _4587_ (.A0(net323),
    .A1(net385),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][7] ),
    .S0(net153),
    .S1(net162),
    .X(_1579_));
 sky130_fd_sc_hd__mux2_2 _4588_ (.A0(_1579_),
    .A1(_1578_),
    .S(net169),
    .X(_1580_));
 sky130_fd_sc_hd__mux2_1 _4589_ (.A0(\z80.tv80s.i_tv80_core.SP[7] ),
    .A1(_1580_),
    .S(net137),
    .X(_1581_));
 sky130_fd_sc_hd__and2_1 _4590_ (.A(net73),
    .B(_1581_),
    .X(_1582_));
 sky130_fd_sc_hd__or2_1 _4591_ (.A(net73),
    .B(_1581_),
    .X(_1583_));
 sky130_fd_sc_hd__nand2b_1 _4592_ (.A_N(_1582_),
    .B(_1583_),
    .Y(_1584_));
 sky130_fd_sc_hd__a21o_1 _4593_ (.A1(_1569_),
    .A2(_1571_),
    .B1(_1568_),
    .X(_1585_));
 sky130_fd_sc_hd__xnor2_1 _4594_ (.A(_1584_),
    .B(_1585_),
    .Y(_1586_));
 sky130_fd_sc_hd__a22o_1 _4595_ (.A1(net751),
    .A2(_1488_),
    .B1(_1586_),
    .B2(_1473_),
    .X(_1587_));
 sky130_fd_sc_hd__mux2_1 _4596_ (.A0(net751),
    .A1(net8),
    .S(_1478_),
    .X(_1588_));
 sky130_fd_sc_hd__mux2_1 _4597_ (.A0(_1587_),
    .A1(_1588_),
    .S(net102),
    .X(_1589_));
 sky130_fd_sc_hd__mux2_1 _4598_ (.A0(\z80.tv80s.di_reg[7] ),
    .A1(_1589_),
    .S(_1465_),
    .X(_1590_));
 sky130_fd_sc_hd__mux2_1 _4599_ (.A0(net751),
    .A1(_1590_),
    .S(net111),
    .X(_0183_));
 sky130_fd_sc_hd__mux4_1 _4600_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][0] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ),
    .S0(net161),
    .S1(net152),
    .X(_1591_));
 sky130_fd_sc_hd__mux4_1 _4601_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][0] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ),
    .S0(net161),
    .S1(net152),
    .X(_1592_));
 sky130_fd_sc_hd__mux2_2 _4602_ (.A0(_1592_),
    .A1(_1591_),
    .S(net169),
    .X(_1593_));
 sky130_fd_sc_hd__mux2_1 _4603_ (.A0(\z80.tv80s.i_tv80_core.SP[8] ),
    .A1(_1593_),
    .S(net138),
    .X(_1594_));
 sky130_fd_sc_hd__nand2_2 _4604_ (.A(net73),
    .B(_1594_),
    .Y(_1595_));
 sky130_fd_sc_hd__or2_1 _4605_ (.A(net73),
    .B(_1594_),
    .X(_1596_));
 sky130_fd_sc_hd__nand2_1 _4606_ (.A(_1595_),
    .B(_1596_),
    .Y(_1597_));
 sky130_fd_sc_hd__a21oi_1 _4607_ (.A1(_1583_),
    .A2(_1585_),
    .B1(_1582_),
    .Y(_1598_));
 sky130_fd_sc_hd__or2_1 _4608_ (.A(_1597_),
    .B(_1598_),
    .X(_1599_));
 sky130_fd_sc_hd__nand2_1 _4609_ (.A(_1597_),
    .B(_1598_),
    .Y(_1600_));
 sky130_fd_sc_hd__and2_1 _4610_ (.A(_1599_),
    .B(_1600_),
    .X(_1601_));
 sky130_fd_sc_hd__and3_1 _4611_ (.A(_1475_),
    .B(_1599_),
    .C(_1600_),
    .X(_1602_));
 sky130_fd_sc_hd__or2_1 _4612_ (.A(net102),
    .B(_1488_),
    .X(_1603_));
 sky130_fd_sc_hd__nor3_1 _4613_ (.A(_0627_),
    .B(_0632_),
    .C(_0634_),
    .Y(_1604_));
 sky130_fd_sc_hd__or4_1 _4614_ (.A(_2773_),
    .B(_2812_),
    .C(_0628_),
    .D(_0635_),
    .X(_1605_));
 sky130_fd_sc_hd__or4_1 _4615_ (.A(_2815_),
    .B(_2817_),
    .C(_2823_),
    .D(_1605_),
    .X(_1606_));
 sky130_fd_sc_hd__nor2_1 _4616_ (.A(_0625_),
    .B(_1606_),
    .Y(_1607_));
 sky130_fd_sc_hd__and4bb_2 _4617_ (.A_N(_2831_),
    .B_N(_0447_),
    .C(_1604_),
    .D(_1607_),
    .X(_1608_));
 sky130_fd_sc_hd__and3_1 _4618_ (.A(_2896_),
    .B(net107),
    .C(_0396_),
    .X(_1609_));
 sky130_fd_sc_hd__o21a_4 _4619_ (.A1(_1608_),
    .A2(_1609_),
    .B1(net136),
    .X(_1610_));
 sky130_fd_sc_hd__o21ai_4 _4620_ (.A1(_1608_),
    .A2(_1609_),
    .B1(net136),
    .Y(_1611_));
 sky130_fd_sc_hd__a211o_1 _4621_ (.A1(net607),
    .A2(_1603_),
    .B1(_1610_),
    .C1(_1602_),
    .X(_1612_));
 sky130_fd_sc_hd__a21oi_1 _4622_ (.A1(_2733_),
    .A2(_1610_),
    .B1(net156),
    .Y(_1613_));
 sky130_fd_sc_hd__a22o_1 _4623_ (.A1(net156),
    .A2(net607),
    .B1(_1612_),
    .B2(_1613_),
    .X(_0184_));
 sky130_fd_sc_hd__mux4_1 _4624_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][1] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][1] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ),
    .S0(net152),
    .S1(net161),
    .X(_1614_));
 sky130_fd_sc_hd__mux4_1 _4625_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][1] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][1] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ),
    .S0(net152),
    .S1(net161),
    .X(_1615_));
 sky130_fd_sc_hd__mux2_2 _4626_ (.A0(_1615_),
    .A1(_1614_),
    .S(net169),
    .X(_1616_));
 sky130_fd_sc_hd__mux2_1 _4627_ (.A0(\z80.tv80s.i_tv80_core.SP[9] ),
    .A1(_1616_),
    .S(net138),
    .X(_1617_));
 sky130_fd_sc_hd__nor2_1 _4628_ (.A(net73),
    .B(_1617_),
    .Y(_1618_));
 sky130_fd_sc_hd__nand2_1 _4629_ (.A(net73),
    .B(_1617_),
    .Y(_1619_));
 sky130_fd_sc_hd__and2b_1 _4630_ (.A_N(_1618_),
    .B(_1619_),
    .X(_1620_));
 sky130_fd_sc_hd__nand2_1 _4631_ (.A(_1595_),
    .B(_1599_),
    .Y(_1621_));
 sky130_fd_sc_hd__xor2_1 _4632_ (.A(_1620_),
    .B(_1621_),
    .X(_1622_));
 sky130_fd_sc_hd__a22o_1 _4633_ (.A1(net671),
    .A2(_1488_),
    .B1(_1622_),
    .B2(_1473_),
    .X(_1623_));
 sky130_fd_sc_hd__a21o_1 _4634_ (.A1(net671),
    .A2(net102),
    .B1(_1610_),
    .X(_1624_));
 sky130_fd_sc_hd__a21oi_1 _4635_ (.A1(net100),
    .A2(_1623_),
    .B1(_1624_),
    .Y(_1625_));
 sky130_fd_sc_hd__a21oi_1 _4636_ (.A1(_2732_),
    .A2(_1610_),
    .B1(_1625_),
    .Y(_1626_));
 sky130_fd_sc_hd__mux2_1 _4637_ (.A0(net671),
    .A1(_1626_),
    .S(net111),
    .X(_0185_));
 sky130_fd_sc_hd__mux4_1 _4638_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][2] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ),
    .S0(net152),
    .S1(net161),
    .X(_1627_));
 sky130_fd_sc_hd__mux4_1 _4639_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][2] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ),
    .S0(net152),
    .S1(net161),
    .X(_1628_));
 sky130_fd_sc_hd__mux2_2 _4640_ (.A0(_1628_),
    .A1(_1627_),
    .S(net169),
    .X(_1629_));
 sky130_fd_sc_hd__mux2_1 _4641_ (.A0(\z80.tv80s.i_tv80_core.SP[10] ),
    .A1(_1629_),
    .S(net138),
    .X(_1630_));
 sky130_fd_sc_hd__nand2_1 _4642_ (.A(net73),
    .B(_1630_),
    .Y(_1631_));
 sky130_fd_sc_hd__or2_1 _4643_ (.A(net73),
    .B(_1630_),
    .X(_1632_));
 sky130_fd_sc_hd__nand2_1 _4644_ (.A(_1631_),
    .B(_1632_),
    .Y(_1633_));
 sky130_fd_sc_hd__o31a_1 _4645_ (.A1(_1597_),
    .A2(_1598_),
    .A3(_1618_),
    .B1(_1619_),
    .X(_1634_));
 sky130_fd_sc_hd__a21oi_1 _4646_ (.A1(_1595_),
    .A2(_1634_),
    .B1(_1633_),
    .Y(_1635_));
 sky130_fd_sc_hd__and3_1 _4647_ (.A(_1595_),
    .B(_1633_),
    .C(_1634_),
    .X(_1636_));
 sky130_fd_sc_hd__nor2_1 _4648_ (.A(_1635_),
    .B(_1636_),
    .Y(_1637_));
 sky130_fd_sc_hd__a22o_1 _4649_ (.A1(net737),
    .A2(_1488_),
    .B1(_1637_),
    .B2(_1473_),
    .X(_1638_));
 sky130_fd_sc_hd__a21o_1 _4650_ (.A1(net737),
    .A2(net102),
    .B1(_1610_),
    .X(_1639_));
 sky130_fd_sc_hd__a21oi_1 _4651_ (.A1(net100),
    .A2(_1638_),
    .B1(_1639_),
    .Y(_1640_));
 sky130_fd_sc_hd__a21oi_1 _4652_ (.A1(_2735_),
    .A2(_1610_),
    .B1(_1640_),
    .Y(_1641_));
 sky130_fd_sc_hd__mux2_1 _4653_ (.A0(net737),
    .A1(_1641_),
    .S(net111),
    .X(_0186_));
 sky130_fd_sc_hd__mux4_1 _4654_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][3] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][3] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][3] ),
    .S0(net152),
    .S1(net161),
    .X(_1642_));
 sky130_fd_sc_hd__mux4_1 _4655_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][3] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][3] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ),
    .S0(net152),
    .S1(net161),
    .X(_1643_));
 sky130_fd_sc_hd__mux2_2 _4656_ (.A0(_1643_),
    .A1(_1642_),
    .S(net169),
    .X(_1644_));
 sky130_fd_sc_hd__mux2_1 _4657_ (.A0(\z80.tv80s.i_tv80_core.SP[11] ),
    .A1(_1644_),
    .S(net138),
    .X(_1645_));
 sky130_fd_sc_hd__nor2_1 _4658_ (.A(net73),
    .B(_1645_),
    .Y(_1646_));
 sky130_fd_sc_hd__nand2_1 _4659_ (.A(net73),
    .B(_1645_),
    .Y(_1647_));
 sky130_fd_sc_hd__and2b_1 _4660_ (.A_N(_1646_),
    .B(_1647_),
    .X(_1648_));
 sky130_fd_sc_hd__a21o_1 _4661_ (.A1(net73),
    .A2(_1630_),
    .B1(_1635_),
    .X(_1649_));
 sky130_fd_sc_hd__xor2_1 _4662_ (.A(_1648_),
    .B(_1649_),
    .X(_1650_));
 sky130_fd_sc_hd__a22o_1 _4663_ (.A1(net697),
    .A2(_1488_),
    .B1(_1650_),
    .B2(_1473_),
    .X(_1651_));
 sky130_fd_sc_hd__a21o_1 _4664_ (.A1(net697),
    .A2(net102),
    .B1(_1610_),
    .X(_1652_));
 sky130_fd_sc_hd__a21oi_1 _4665_ (.A1(net100),
    .A2(_1651_),
    .B1(_1652_),
    .Y(_1653_));
 sky130_fd_sc_hd__a21oi_1 _4666_ (.A1(_2734_),
    .A2(_1610_),
    .B1(_1653_),
    .Y(_1654_));
 sky130_fd_sc_hd__mux2_1 _4667_ (.A0(net697),
    .A1(_1654_),
    .S(net111),
    .X(_0187_));
 sky130_fd_sc_hd__mux4_1 _4668_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][4] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][4] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][4] ),
    .S0(net152),
    .S1(net161),
    .X(_1655_));
 sky130_fd_sc_hd__mux4_1 _4669_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][4] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][4] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][4] ),
    .S0(net152),
    .S1(net161),
    .X(_1656_));
 sky130_fd_sc_hd__mux2_2 _4670_ (.A0(_1656_),
    .A1(_1655_),
    .S(net169),
    .X(_1657_));
 sky130_fd_sc_hd__mux2_1 _4671_ (.A0(\z80.tv80s.i_tv80_core.SP[12] ),
    .A1(_1657_),
    .S(net138),
    .X(_1658_));
 sky130_fd_sc_hd__nand2_1 _4672_ (.A(net73),
    .B(_1658_),
    .Y(_1659_));
 sky130_fd_sc_hd__or2_1 _4673_ (.A(net73),
    .B(_1658_),
    .X(_1660_));
 sky130_fd_sc_hd__nand2_1 _4674_ (.A(_1659_),
    .B(_1660_),
    .Y(_1661_));
 sky130_fd_sc_hd__a211o_1 _4675_ (.A1(_1595_),
    .A2(_1634_),
    .B1(_1646_),
    .C1(_1633_),
    .X(_1662_));
 sky130_fd_sc_hd__and3_1 _4676_ (.A(_1631_),
    .B(_1647_),
    .C(_1662_),
    .X(_1663_));
 sky130_fd_sc_hd__xor2_1 _4677_ (.A(_1661_),
    .B(_1663_),
    .X(_1664_));
 sky130_fd_sc_hd__a22o_1 _4678_ (.A1(net718),
    .A2(_1488_),
    .B1(_1664_),
    .B2(_1473_),
    .X(_1665_));
 sky130_fd_sc_hd__a21o_1 _4679_ (.A1(net718),
    .A2(net102),
    .B1(_1610_),
    .X(_1666_));
 sky130_fd_sc_hd__a21oi_1 _4680_ (.A1(net100),
    .A2(_1665_),
    .B1(_1666_),
    .Y(_1667_));
 sky130_fd_sc_hd__a21oi_1 _4681_ (.A1(_2736_),
    .A2(_1610_),
    .B1(_1667_),
    .Y(_1668_));
 sky130_fd_sc_hd__mux2_1 _4682_ (.A0(net718),
    .A1(_1668_),
    .S(net111),
    .X(_0188_));
 sky130_fd_sc_hd__mux4_1 _4683_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][5] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][5] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ),
    .S0(net152),
    .S1(net161),
    .X(_1669_));
 sky130_fd_sc_hd__mux4_1 _4684_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][5] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][5] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ),
    .S0(net152),
    .S1(net161),
    .X(_1670_));
 sky130_fd_sc_hd__mux2_2 _4685_ (.A0(_1670_),
    .A1(_1669_),
    .S(net169),
    .X(_1671_));
 sky130_fd_sc_hd__mux2_1 _4686_ (.A0(\z80.tv80s.i_tv80_core.SP[13] ),
    .A1(_1671_),
    .S(net138),
    .X(_1672_));
 sky130_fd_sc_hd__nor2_1 _4687_ (.A(net73),
    .B(_1672_),
    .Y(_1673_));
 sky130_fd_sc_hd__nand2_1 _4688_ (.A(net73),
    .B(_1672_),
    .Y(_1674_));
 sky130_fd_sc_hd__nand2b_1 _4689_ (.A_N(_1673_),
    .B(_1674_),
    .Y(_1675_));
 sky130_fd_sc_hd__o21ai_1 _4690_ (.A1(_1661_),
    .A2(_1663_),
    .B1(_1659_),
    .Y(_1676_));
 sky130_fd_sc_hd__xnor2_1 _4691_ (.A(_1675_),
    .B(_1676_),
    .Y(_1677_));
 sky130_fd_sc_hd__a221o_1 _4692_ (.A1(net727),
    .A2(_1603_),
    .B1(_1677_),
    .B2(_1475_),
    .C1(_1610_),
    .X(_1678_));
 sky130_fd_sc_hd__o21a_1 _4693_ (.A1(\z80.tv80s.di_reg[5] ),
    .A2(_1611_),
    .B1(_1678_),
    .X(_1679_));
 sky130_fd_sc_hd__mux2_1 _4694_ (.A0(net727),
    .A1(_1679_),
    .S(net111),
    .X(_0189_));
 sky130_fd_sc_hd__mux4_1 _4695_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][6] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][6] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ),
    .S0(net152),
    .S1(net161),
    .X(_1680_));
 sky130_fd_sc_hd__mux4_1 _4696_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][6] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][6] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ),
    .S0(net152),
    .S1(net161),
    .X(_1681_));
 sky130_fd_sc_hd__mux2_2 _4697_ (.A0(_1681_),
    .A1(_1680_),
    .S(net169),
    .X(_1682_));
 sky130_fd_sc_hd__mux2_1 _4698_ (.A0(\z80.tv80s.i_tv80_core.SP[14] ),
    .A1(_1682_),
    .S(net138),
    .X(_1683_));
 sky130_fd_sc_hd__nand2_1 _4699_ (.A(net73),
    .B(_1683_),
    .Y(_1684_));
 sky130_fd_sc_hd__or2_1 _4700_ (.A(_1577_),
    .B(_1683_),
    .X(_1685_));
 sky130_fd_sc_hd__nand2_1 _4701_ (.A(_1684_),
    .B(_1685_),
    .Y(_1686_));
 sky130_fd_sc_hd__a311o_1 _4702_ (.A1(_1631_),
    .A2(_1647_),
    .A3(_1662_),
    .B1(_1673_),
    .C1(_1661_),
    .X(_1687_));
 sky130_fd_sc_hd__and3_1 _4703_ (.A(_1659_),
    .B(_1674_),
    .C(_1687_),
    .X(_1688_));
 sky130_fd_sc_hd__a31o_1 _4704_ (.A1(_1659_),
    .A2(_1674_),
    .A3(_1687_),
    .B1(_1686_),
    .X(_1689_));
 sky130_fd_sc_hd__xor2_1 _4705_ (.A(_1686_),
    .B(_1688_),
    .X(_1690_));
 sky130_fd_sc_hd__a22o_1 _4706_ (.A1(net640),
    .A2(_1488_),
    .B1(_1690_),
    .B2(_1473_),
    .X(_1691_));
 sky130_fd_sc_hd__a21o_1 _4707_ (.A1(net640),
    .A2(net102),
    .B1(_1610_),
    .X(_1692_));
 sky130_fd_sc_hd__a21o_1 _4708_ (.A1(net100),
    .A2(_1691_),
    .B1(_1692_),
    .X(_1693_));
 sky130_fd_sc_hd__o21a_1 _4709_ (.A1(\z80.tv80s.di_reg[6] ),
    .A2(_1611_),
    .B1(_1693_),
    .X(_1694_));
 sky130_fd_sc_hd__mux2_1 _4710_ (.A0(net640),
    .A1(_1694_),
    .S(net111),
    .X(_0190_));
 sky130_fd_sc_hd__mux4_1 _4711_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][7] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][7] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][7] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][7] ),
    .S0(\z80.tv80s.i_tv80_core.RegAddrC[0] ),
    .S1(\z80.tv80s.i_tv80_core.RegAddrC[1] ),
    .X(_1695_));
 sky130_fd_sc_hd__mux4_1 _4712_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][7] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][7] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][7] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][7] ),
    .S0(net152),
    .S1(net161),
    .X(_1696_));
 sky130_fd_sc_hd__mux2_2 _4713_ (.A0(_1696_),
    .A1(_1695_),
    .S(\z80.tv80s.i_tv80_core.RegAddrC[2] ),
    .X(_1697_));
 sky130_fd_sc_hd__mux2_1 _4714_ (.A0(\z80.tv80s.i_tv80_core.SP[15] ),
    .A1(_1697_),
    .S(net138),
    .X(_1698_));
 sky130_fd_sc_hd__xor2_1 _4715_ (.A(_1577_),
    .B(_1698_),
    .X(_1699_));
 sky130_fd_sc_hd__and3_1 _4716_ (.A(_1684_),
    .B(_1689_),
    .C(_1699_),
    .X(_1700_));
 sky130_fd_sc_hd__a21oi_1 _4717_ (.A1(_1684_),
    .A2(_1689_),
    .B1(_1699_),
    .Y(_1701_));
 sky130_fd_sc_hd__or2_1 _4718_ (.A(_1700_),
    .B(_1701_),
    .X(_1702_));
 sky130_fd_sc_hd__a22o_1 _4719_ (.A1(net675),
    .A2(_1488_),
    .B1(_1702_),
    .B2(_1473_),
    .X(_1703_));
 sky130_fd_sc_hd__a21o_1 _4720_ (.A1(net675),
    .A2(net102),
    .B1(_1610_),
    .X(_1704_));
 sky130_fd_sc_hd__a21o_1 _4721_ (.A1(net100),
    .A2(_1703_),
    .B1(_1704_),
    .X(_1705_));
 sky130_fd_sc_hd__o21a_1 _4722_ (.A1(\z80.tv80s.di_reg[7] ),
    .A2(_1611_),
    .B1(net111),
    .X(_1706_));
 sky130_fd_sc_hd__a22o_1 _4723_ (.A1(net156),
    .A2(net675),
    .B1(_1705_),
    .B2(_1706_),
    .X(_0191_));
 sky130_fd_sc_hd__a22o_1 _4724_ (.A1(net160),
    .A2(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .B1(net53),
    .B2(_1457_),
    .X(_0192_));
 sky130_fd_sc_hd__or2_1 _4725_ (.A(net124),
    .B(net151),
    .X(_1707_));
 sky130_fd_sc_hd__or4_1 _4726_ (.A(_2769_),
    .B(_2794_),
    .C(_2809_),
    .D(_2881_),
    .X(_1708_));
 sky130_fd_sc_hd__or3_1 _4727_ (.A(_2803_),
    .B(_2823_),
    .C(_1708_),
    .X(_1709_));
 sky130_fd_sc_hd__or4_1 _4728_ (.A(_2759_),
    .B(_2765_),
    .C(_2815_),
    .D(_2886_),
    .X(_1710_));
 sky130_fd_sc_hd__or4_1 _4729_ (.A(_2831_),
    .B(_2867_),
    .C(_1709_),
    .D(_1710_),
    .X(_1711_));
 sky130_fd_sc_hd__a211o_1 _4730_ (.A1(net116),
    .A2(_2860_),
    .B1(_1420_),
    .C1(_1711_),
    .X(_1712_));
 sky130_fd_sc_hd__mux2_1 _4731_ (.A0(\z80.tv80s.i_tv80_core.IR[7] ),
    .A1(net124),
    .S(_0480_),
    .X(_1713_));
 sky130_fd_sc_hd__a22o_1 _4732_ (.A1(_1707_),
    .A2(_1712_),
    .B1(_1713_),
    .B2(_2859_),
    .X(_1714_));
 sky130_fd_sc_hd__a31o_1 _4733_ (.A1(net126),
    .A2(_2856_),
    .A3(_0384_),
    .B1(_0434_),
    .X(_1715_));
 sky130_fd_sc_hd__o21a_1 _4734_ (.A1(net125),
    .A2(_1453_),
    .B1(_1715_),
    .X(_1716_));
 sky130_fd_sc_hd__nand2_1 _4735_ (.A(_2702_),
    .B(_0384_),
    .Y(_1717_));
 sky130_fd_sc_hd__a221o_1 _4736_ (.A1(_2844_),
    .A2(_1707_),
    .B1(_1717_),
    .B2(_1452_),
    .C1(_1187_),
    .X(_1718_));
 sky130_fd_sc_hd__nor2_1 _4737_ (.A(net126),
    .B(_0470_),
    .Y(_1719_));
 sky130_fd_sc_hd__or4_1 _4738_ (.A(_1439_),
    .B(_1716_),
    .C(_1718_),
    .D(_1719_),
    .X(_1720_));
 sky130_fd_sc_hd__or2_1 _4739_ (.A(net124),
    .B(_1440_),
    .X(_1721_));
 sky130_fd_sc_hd__a211o_1 _4740_ (.A1(_2920_),
    .A2(_0384_),
    .B1(_1175_),
    .C1(_1436_),
    .X(_1722_));
 sky130_fd_sc_hd__a221o_1 _4741_ (.A1(net135),
    .A2(_2933_),
    .B1(_1722_),
    .B2(net124),
    .C1(_0497_),
    .X(_1723_));
 sky130_fd_sc_hd__a22o_1 _4742_ (.A1(net163),
    .A2(_1714_),
    .B1(_1723_),
    .B2(net166),
    .X(_1724_));
 sky130_fd_sc_hd__a31o_1 _4743_ (.A1(_0377_),
    .A2(_1720_),
    .A3(_1721_),
    .B1(_1724_),
    .X(_1725_));
 sky130_fd_sc_hd__a22o_1 _4744_ (.A1(net160),
    .A2(net154),
    .B1(net53),
    .B2(_1725_),
    .X(_0193_));
 sky130_fd_sc_hd__a22o_1 _4745_ (.A1(net160),
    .A2(net835),
    .B1(net53),
    .B2(_1445_),
    .X(_0194_));
 sky130_fd_sc_hd__o2bb2a_1 _4746_ (.A1_N(net165),
    .A2_N(_1171_),
    .B1(_0470_),
    .B2(net106),
    .X(_1726_));
 sky130_fd_sc_hd__o21ai_1 _4747_ (.A1(_2708_),
    .A2(_1438_),
    .B1(_1726_),
    .Y(_1727_));
 sky130_fd_sc_hd__a22o_1 _4748_ (.A1(net160),
    .A2(net831),
    .B1(net53),
    .B2(_1727_),
    .X(_0195_));
 sky130_fd_sc_hd__or3_1 _4749_ (.A(_1187_),
    .B(_1428_),
    .C(_1453_),
    .X(_1728_));
 sky130_fd_sc_hd__or3_1 _4750_ (.A(_0612_),
    .B(_1172_),
    .C(_1424_),
    .X(_1729_));
 sky130_fd_sc_hd__a221o_1 _4751_ (.A1(net107),
    .A2(_1728_),
    .B1(_1729_),
    .B2(net166),
    .C1(_1423_),
    .X(_1730_));
 sky130_fd_sc_hd__a22o_1 _4752_ (.A1(net159),
    .A2(net845),
    .B1(net53),
    .B2(_1730_),
    .X(_0196_));
 sky130_fd_sc_hd__a2bb2o_1 _4753_ (.A1_N(_2930_),
    .A2_N(_0587_),
    .B1(net144),
    .B2(_2759_),
    .X(_1731_));
 sky130_fd_sc_hd__a31o_1 _4754_ (.A1(_0466_),
    .A2(_0556_),
    .A3(_0616_),
    .B1(_1731_),
    .X(_1732_));
 sky130_fd_sc_hd__a21oi_2 _4755_ (.A1(_2913_),
    .A2(_0454_),
    .B1(_1732_),
    .Y(_1733_));
 sky130_fd_sc_hd__o21ai_4 _4756_ (.A1(net115),
    .A2(_1733_),
    .B1(_0657_),
    .Y(_1734_));
 sky130_fd_sc_hd__nand2_1 _4757_ (.A(net92),
    .B(_1468_),
    .Y(_1735_));
 sky130_fd_sc_hd__a211oi_1 _4758_ (.A1(_2702_),
    .A2(_2812_),
    .B1(_2815_),
    .C1(net115),
    .Y(_1736_));
 sky130_fd_sc_hd__and3_1 _4759_ (.A(_0384_),
    .B(_0466_),
    .C(_0626_),
    .X(_1737_));
 sky130_fd_sc_hd__and4b_1 _4760_ (.A_N(_0631_),
    .B(_1604_),
    .C(_1736_),
    .D(_1737_),
    .X(_1738_));
 sky130_fd_sc_hd__or2_2 _4761_ (.A(_1486_),
    .B(_1738_),
    .X(_1739_));
 sky130_fd_sc_hd__and2_2 _4762_ (.A(\z80.tv80s.i_tv80_core.NMICycle ),
    .B(_0646_),
    .X(_1740_));
 sky130_fd_sc_hd__nor2_2 _4763_ (.A(net63),
    .B(_1740_),
    .Y(_1741_));
 sky130_fd_sc_hd__and3_2 _4764_ (.A(net143),
    .B(\z80.tv80s.i_tv80_core.IntCycle ),
    .C(\z80.tv80s.i_tv80_core.IStatus[1] ),
    .X(_1742_));
 sky130_fd_sc_hd__nand3_2 _4765_ (.A(net143),
    .B(\z80.tv80s.i_tv80_core.IntCycle ),
    .C(\z80.tv80s.i_tv80_core.IStatus[1] ),
    .Y(_1743_));
 sky130_fd_sc_hd__nor2_2 _4766_ (.A(_0406_),
    .B(_0439_),
    .Y(_1744_));
 sky130_fd_sc_hd__or2_2 _4767_ (.A(_0406_),
    .B(_0439_),
    .X(_1745_));
 sky130_fd_sc_hd__nor3b_4 _4768_ (.A(_0440_),
    .B(_0405_),
    .C_N(_0389_),
    .Y(_1746_));
 sky130_fd_sc_hd__nor2_8 _4769_ (.A(_0389_),
    .B(_0440_),
    .Y(_1747_));
 sky130_fd_sc_hd__and3_4 _4770_ (.A(_0389_),
    .B(_0405_),
    .C(_0439_),
    .X(_1748_));
 sky130_fd_sc_hd__and3_4 _4771_ (.A(_0390_),
    .B(_0406_),
    .C(_0440_),
    .X(_1749_));
 sky130_fd_sc_hd__or4_1 _4772_ (.A(net115),
    .B(_2879_),
    .C(_2886_),
    .D(_0625_),
    .X(_1750_));
 sky130_fd_sc_hd__a2111o_1 _4773_ (.A1(_2702_),
    .A2(_2812_),
    .B1(_2815_),
    .C1(_0631_),
    .D1(_1750_),
    .X(_1751_));
 sky130_fd_sc_hd__nor2_1 _4774_ (.A(_1483_),
    .B(_1751_),
    .Y(_1752_));
 sky130_fd_sc_hd__o21a_4 _4775_ (.A1(_0559_),
    .A2(_1752_),
    .B1(_0472_),
    .X(_1753_));
 sky130_fd_sc_hd__inv_2 _4776_ (.A(_1753_),
    .Y(_1754_));
 sky130_fd_sc_hd__xor2_1 _4777_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .B(_1753_),
    .X(_1755_));
 sky130_fd_sc_hd__mux2_1 _4778_ (.A0(\z80.tv80s.i_tv80_core.PC[0] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .S(_0446_),
    .X(_1756_));
 sky130_fd_sc_hd__or2_1 _4779_ (.A(net104),
    .B(_1468_),
    .X(_1757_));
 sky130_fd_sc_hd__o211a_1 _4780_ (.A1(_0443_),
    .A2(_1756_),
    .B1(_1757_),
    .C1(net58),
    .X(_1758_));
 sky130_fd_sc_hd__a221o_1 _4781_ (.A1(\z80.tv80s.i_tv80_core.SP[0] ),
    .A2(_1746_),
    .B1(_1747_),
    .B2(_1468_),
    .C1(net57),
    .X(_1759_));
 sky130_fd_sc_hd__a221o_1 _4782_ (.A1(\z80.tv80s.di_reg[0] ),
    .A2(_1748_),
    .B1(_1749_),
    .B2(_1755_),
    .C1(_1759_),
    .X(_1760_));
 sky130_fd_sc_hd__o22a_1 _4783_ (.A1(\z80.tv80s.i_tv80_core.PC[0] ),
    .A2(_1745_),
    .B1(_1758_),
    .B2(_1760_),
    .X(_1761_));
 sky130_fd_sc_hd__mux2_1 _4784_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .A1(_1761_),
    .S(net98),
    .X(_1762_));
 sky130_fd_sc_hd__a22o_1 _4785_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .A2(net63),
    .B1(net60),
    .B2(_1762_),
    .X(_1763_));
 sky130_fd_sc_hd__a21bo_1 _4786_ (.A1(net86),
    .A2(_1763_),
    .B1_N(_1735_),
    .X(_1764_));
 sky130_fd_sc_hd__mux2_1 _4787_ (.A0(_1764_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .S(net67),
    .X(_1765_));
 sky130_fd_sc_hd__mux2_1 _4788_ (.A0(net599),
    .A1(_1765_),
    .S(net53),
    .X(_0197_));
 sky130_fd_sc_hd__nand2_1 _4789_ (.A(net92),
    .B(_1494_),
    .Y(_1766_));
 sky130_fd_sc_hd__a21o_1 _4790_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .A2(_1742_),
    .B1(_1740_),
    .X(_1767_));
 sky130_fd_sc_hd__a22o_1 _4791_ (.A1(_1494_),
    .A2(_1747_),
    .B1(_1748_),
    .B2(\z80.tv80s.di_reg[1] ),
    .X(_1768_));
 sky130_fd_sc_hd__mux2_1 _4792_ (.A0(\z80.tv80s.i_tv80_core.PC[1] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .S(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(_1769_));
 sky130_fd_sc_hd__mux2_1 _4793_ (.A0(_1494_),
    .A1(_1769_),
    .S(net104),
    .X(_1770_));
 sky130_fd_sc_hd__and3_1 _4794_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .C(_1753_),
    .X(_1771_));
 sky130_fd_sc_hd__a21oi_1 _4795_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .A2(_1753_),
    .B1(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .Y(_1772_));
 sky130_fd_sc_hd__nor2_1 _4796_ (.A(_1771_),
    .B(_1772_),
    .Y(_1773_));
 sky130_fd_sc_hd__a22o_1 _4797_ (.A1(net58),
    .A2(_1770_),
    .B1(_1773_),
    .B2(_1749_),
    .X(_1774_));
 sky130_fd_sc_hd__a211o_1 _4798_ (.A1(\z80.tv80s.i_tv80_core.SP[1] ),
    .A2(_1746_),
    .B1(_1768_),
    .C1(_1774_),
    .X(_1775_));
 sky130_fd_sc_hd__a21o_1 _4799_ (.A1(\z80.tv80s.i_tv80_core.PC[1] ),
    .A2(net57),
    .B1(_1775_),
    .X(_1776_));
 sky130_fd_sc_hd__a21o_1 _4800_ (.A1(net98),
    .A2(_1776_),
    .B1(_1767_),
    .X(_1777_));
 sky130_fd_sc_hd__mux2_1 _4801_ (.A0(_1777_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .S(net63),
    .X(_1778_));
 sky130_fd_sc_hd__a21bo_1 _4802_ (.A1(net86),
    .A2(_1778_),
    .B1_N(_1766_),
    .X(_1779_));
 sky130_fd_sc_hd__mux2_1 _4803_ (.A0(_1779_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .S(net67),
    .X(_1780_));
 sky130_fd_sc_hd__mux2_1 _4804_ (.A0(net558),
    .A1(_1780_),
    .S(net53),
    .X(_0198_));
 sky130_fd_sc_hd__nand2_1 _4805_ (.A(net92),
    .B(_1507_),
    .Y(_1781_));
 sky130_fd_sc_hd__a21o_1 _4806_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .A2(_1742_),
    .B1(_1740_),
    .X(_1782_));
 sky130_fd_sc_hd__and2_1 _4807_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .B(_1771_),
    .X(_1783_));
 sky130_fd_sc_hd__or2_1 _4808_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .B(_1771_),
    .X(_1784_));
 sky130_fd_sc_hd__and3b_1 _4809_ (.A_N(_1783_),
    .B(_1784_),
    .C(_1749_),
    .X(_1785_));
 sky130_fd_sc_hd__mux2_1 _4810_ (.A0(\z80.tv80s.i_tv80_core.PC[2] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .S(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(_1786_));
 sky130_fd_sc_hd__mux2_1 _4811_ (.A0(_1507_),
    .A1(_1786_),
    .S(net104),
    .X(_1787_));
 sky130_fd_sc_hd__a221o_1 _4812_ (.A1(\z80.tv80s.i_tv80_core.SP[2] ),
    .A2(_1746_),
    .B1(_1747_),
    .B2(_1507_),
    .C1(net57),
    .X(_1788_));
 sky130_fd_sc_hd__a22o_1 _4813_ (.A1(\z80.tv80s.di_reg[2] ),
    .A2(_1748_),
    .B1(_1787_),
    .B2(net58),
    .X(_1789_));
 sky130_fd_sc_hd__or3_1 _4814_ (.A(_1785_),
    .B(_1788_),
    .C(_1789_),
    .X(_1790_));
 sky130_fd_sc_hd__nand2_1 _4815_ (.A(_2741_),
    .B(net57),
    .Y(_1791_));
 sky130_fd_sc_hd__a31o_1 _4816_ (.A1(net98),
    .A2(_1790_),
    .A3(_1791_),
    .B1(_1782_),
    .X(_1792_));
 sky130_fd_sc_hd__mux2_1 _4817_ (.A0(_1792_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .S(net63),
    .X(_1793_));
 sky130_fd_sc_hd__a21bo_1 _4818_ (.A1(net86),
    .A2(_1793_),
    .B1_N(_1781_),
    .X(_1794_));
 sky130_fd_sc_hd__mux2_1 _4819_ (.A0(_1794_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .S(net67),
    .X(_1795_));
 sky130_fd_sc_hd__mux2_1 _4820_ (.A0(net526),
    .A1(_1795_),
    .S(net53),
    .X(_0199_));
 sky130_fd_sc_hd__nand2_1 _4821_ (.A(net92),
    .B(_1521_),
    .Y(_1796_));
 sky130_fd_sc_hd__or2_1 _4822_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .B(_1783_),
    .X(_1797_));
 sky130_fd_sc_hd__and3_1 _4823_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .C(_1771_),
    .X(_1798_));
 sky130_fd_sc_hd__and3b_1 _4824_ (.A_N(_1798_),
    .B(_1749_),
    .C(_1797_),
    .X(_1799_));
 sky130_fd_sc_hd__mux2_1 _4825_ (.A0(\z80.tv80s.i_tv80_core.PC[3] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .S(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(_1800_));
 sky130_fd_sc_hd__mux2_1 _4826_ (.A0(_1521_),
    .A1(_1800_),
    .S(net104),
    .X(_1801_));
 sky130_fd_sc_hd__a221o_1 _4827_ (.A1(\z80.tv80s.i_tv80_core.SP[3] ),
    .A2(_1746_),
    .B1(_1747_),
    .B2(_1521_),
    .C1(net57),
    .X(_1802_));
 sky130_fd_sc_hd__a22o_1 _4828_ (.A1(\z80.tv80s.di_reg[3] ),
    .A2(_1748_),
    .B1(_1801_),
    .B2(net58),
    .X(_1803_));
 sky130_fd_sc_hd__or3_1 _4829_ (.A(_1799_),
    .B(_1802_),
    .C(_1803_),
    .X(_1804_));
 sky130_fd_sc_hd__a21oi_1 _4830_ (.A1(_2742_),
    .A2(net57),
    .B1(_1742_),
    .Y(_1805_));
 sky130_fd_sc_hd__a22o_1 _4831_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .A2(_1742_),
    .B1(_1804_),
    .B2(_1805_),
    .X(_1806_));
 sky130_fd_sc_hd__a22o_1 _4832_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .A2(net63),
    .B1(net60),
    .B2(_1806_),
    .X(_1807_));
 sky130_fd_sc_hd__a21bo_1 _4833_ (.A1(net86),
    .A2(_1807_),
    .B1_N(_1796_),
    .X(_1808_));
 sky130_fd_sc_hd__mux2_1 _4834_ (.A0(_1808_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .S(net67),
    .X(_1809_));
 sky130_fd_sc_hd__mux2_1 _4835_ (.A0(net568),
    .A1(_1809_),
    .S(net53),
    .X(_0200_));
 sky130_fd_sc_hd__nand2_1 _4836_ (.A(net92),
    .B(_1536_),
    .Y(_1810_));
 sky130_fd_sc_hd__mux2_1 _4837_ (.A0(\z80.tv80s.i_tv80_core.PC[4] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .S(_0446_),
    .X(_1811_));
 sky130_fd_sc_hd__mux2_1 _4838_ (.A0(_1536_),
    .A1(_1811_),
    .S(net104),
    .X(_1812_));
 sky130_fd_sc_hd__and3_1 _4839_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .C(_1783_),
    .X(_1813_));
 sky130_fd_sc_hd__o21ai_1 _4840_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .A2(_1798_),
    .B1(_1749_),
    .Y(_1814_));
 sky130_fd_sc_hd__nor2_1 _4841_ (.A(_1813_),
    .B(_1814_),
    .Y(_1815_));
 sky130_fd_sc_hd__a221o_1 _4842_ (.A1(\z80.tv80s.i_tv80_core.SP[4] ),
    .A2(_1746_),
    .B1(_1747_),
    .B2(_1536_),
    .C1(net57),
    .X(_1816_));
 sky130_fd_sc_hd__a221o_1 _4843_ (.A1(\z80.tv80s.di_reg[4] ),
    .A2(_1748_),
    .B1(_1812_),
    .B2(net58),
    .C1(_1815_),
    .X(_1817_));
 sky130_fd_sc_hd__o22a_1 _4844_ (.A1(\z80.tv80s.i_tv80_core.PC[4] ),
    .A2(_1745_),
    .B1(_1816_),
    .B2(_1817_),
    .X(_1818_));
 sky130_fd_sc_hd__mux2_1 _4845_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .A1(_1818_),
    .S(net98),
    .X(_1819_));
 sky130_fd_sc_hd__a22o_1 _4846_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .A2(net64),
    .B1(net60),
    .B2(_1819_),
    .X(_1820_));
 sky130_fd_sc_hd__a21bo_1 _4847_ (.A1(net86),
    .A2(_1820_),
    .B1_N(_1810_),
    .X(_1821_));
 sky130_fd_sc_hd__mux2_1 _4848_ (.A0(_1821_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .S(net67),
    .X(_1822_));
 sky130_fd_sc_hd__mux2_1 _4849_ (.A0(net545),
    .A1(_1822_),
    .S(net53),
    .X(_0201_));
 sky130_fd_sc_hd__nand2_1 _4850_ (.A(net92),
    .B(_1551_),
    .Y(_1823_));
 sky130_fd_sc_hd__a21o_1 _4851_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .A2(_1742_),
    .B1(_1740_),
    .X(_1824_));
 sky130_fd_sc_hd__mux2_1 _4852_ (.A0(\z80.tv80s.i_tv80_core.PC[5] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .S(_0446_),
    .X(_1825_));
 sky130_fd_sc_hd__mux2_1 _4853_ (.A0(_1551_),
    .A1(_1825_),
    .S(net104),
    .X(_1826_));
 sky130_fd_sc_hd__and2_1 _4854_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .B(_1813_),
    .X(_1827_));
 sky130_fd_sc_hd__o21ai_1 _4855_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .A2(_1813_),
    .B1(_1749_),
    .Y(_1828_));
 sky130_fd_sc_hd__nor2_1 _4856_ (.A(_1827_),
    .B(_1828_),
    .Y(_1829_));
 sky130_fd_sc_hd__a221o_1 _4857_ (.A1(\z80.tv80s.i_tv80_core.SP[5] ),
    .A2(_1746_),
    .B1(_1747_),
    .B2(_1551_),
    .C1(net57),
    .X(_1830_));
 sky130_fd_sc_hd__a221o_1 _4858_ (.A1(\z80.tv80s.di_reg[5] ),
    .A2(_1748_),
    .B1(_1826_),
    .B2(net58),
    .C1(_1829_),
    .X(_1831_));
 sky130_fd_sc_hd__o22a_1 _4859_ (.A1(\z80.tv80s.i_tv80_core.PC[5] ),
    .A2(_1745_),
    .B1(_1830_),
    .B2(_1831_),
    .X(_1832_));
 sky130_fd_sc_hd__a21o_1 _4860_ (.A1(net98),
    .A2(_1832_),
    .B1(_1824_),
    .X(_1833_));
 sky130_fd_sc_hd__mux2_1 _4861_ (.A0(_1833_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .S(net63),
    .X(_1834_));
 sky130_fd_sc_hd__a21bo_1 _4862_ (.A1(net86),
    .A2(_1834_),
    .B1_N(_1823_),
    .X(_1835_));
 sky130_fd_sc_hd__mux2_1 _4863_ (.A0(_1835_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .S(net67),
    .X(_1836_));
 sky130_fd_sc_hd__mux2_1 _4864_ (.A0(net564),
    .A1(_1836_),
    .S(net53),
    .X(_0202_));
 sky130_fd_sc_hd__nand2_1 _4865_ (.A(net92),
    .B(_1566_),
    .Y(_1837_));
 sky130_fd_sc_hd__a21o_1 _4866_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .A2(_1742_),
    .B1(_1740_),
    .X(_1838_));
 sky130_fd_sc_hd__mux2_1 _4867_ (.A0(\z80.tv80s.i_tv80_core.PC[6] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .S(_0446_),
    .X(_1839_));
 sky130_fd_sc_hd__mux2_1 _4868_ (.A0(_1566_),
    .A1(_1839_),
    .S(_0444_),
    .X(_1840_));
 sky130_fd_sc_hd__o21ai_1 _4869_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .A2(_1827_),
    .B1(_1749_),
    .Y(_1841_));
 sky130_fd_sc_hd__a21oi_1 _4870_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .A2(_1827_),
    .B1(_1841_),
    .Y(_1842_));
 sky130_fd_sc_hd__a221o_1 _4871_ (.A1(\z80.tv80s.i_tv80_core.SP[6] ),
    .A2(net56),
    .B1(_1747_),
    .B2(_1566_),
    .C1(net57),
    .X(_1843_));
 sky130_fd_sc_hd__a22o_1 _4872_ (.A1(\z80.tv80s.di_reg[6] ),
    .A2(_1748_),
    .B1(_1840_),
    .B2(net58),
    .X(_1844_));
 sky130_fd_sc_hd__o32a_1 _4873_ (.A1(_1842_),
    .A2(_1843_),
    .A3(_1844_),
    .B1(_1745_),
    .B2(\z80.tv80s.i_tv80_core.PC[6] ),
    .X(_1845_));
 sky130_fd_sc_hd__a21o_1 _4874_ (.A1(net98),
    .A2(_1845_),
    .B1(_1838_),
    .X(_1846_));
 sky130_fd_sc_hd__mux2_1 _4875_ (.A0(_1846_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .S(net63),
    .X(_1847_));
 sky130_fd_sc_hd__a21bo_1 _4876_ (.A1(net86),
    .A2(_1847_),
    .B1_N(_1837_),
    .X(_1848_));
 sky130_fd_sc_hd__mux2_1 _4877_ (.A0(_1848_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .S(net67),
    .X(_1849_));
 sky130_fd_sc_hd__mux2_1 _4878_ (.A0(net547),
    .A1(_1849_),
    .S(net53),
    .X(_0203_));
 sky130_fd_sc_hd__nand2_1 _4879_ (.A(net92),
    .B(_1580_),
    .Y(_1850_));
 sky130_fd_sc_hd__mux2_1 _4880_ (.A0(\z80.tv80s.i_tv80_core.PC[7] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .S(_0446_),
    .X(_1851_));
 sky130_fd_sc_hd__mux2_1 _4881_ (.A0(_1580_),
    .A1(_1851_),
    .S(net104),
    .X(_1852_));
 sky130_fd_sc_hd__a31o_1 _4882_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .A2(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .A3(_1813_),
    .B1(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .X(_1853_));
 sky130_fd_sc_hd__and4_1 _4883_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .C(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .D(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .X(_1854_));
 sky130_fd_sc_hd__and4_1 _4884_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .C(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .D(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .X(_1855_));
 sky130_fd_sc_hd__nand2_1 _4885_ (.A(_1854_),
    .B(_1855_),
    .Y(_1856_));
 sky130_fd_sc_hd__a221o_1 _4886_ (.A1(\z80.tv80s.i_tv80_core.SP[7] ),
    .A2(net56),
    .B1(_1747_),
    .B2(_1580_),
    .C1(net57),
    .X(_1857_));
 sky130_fd_sc_hd__o211a_1 _4887_ (.A1(_1754_),
    .A2(_1856_),
    .B1(_1853_),
    .C1(_1749_),
    .X(_1858_));
 sky130_fd_sc_hd__a221o_1 _4888_ (.A1(\z80.tv80s.di_reg[7] ),
    .A2(_1748_),
    .B1(_1852_),
    .B2(net58),
    .C1(_1858_),
    .X(_1859_));
 sky130_fd_sc_hd__o22a_1 _4889_ (.A1(\z80.tv80s.i_tv80_core.PC[7] ),
    .A2(_1745_),
    .B1(_1857_),
    .B2(_1859_),
    .X(_1860_));
 sky130_fd_sc_hd__mux2_1 _4890_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .A1(_1860_),
    .S(net98),
    .X(_1861_));
 sky130_fd_sc_hd__a22o_1 _4891_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .A2(net63),
    .B1(net60),
    .B2(_1861_),
    .X(_1862_));
 sky130_fd_sc_hd__a21bo_1 _4892_ (.A1(net86),
    .A2(_1862_),
    .B1_N(_1850_),
    .X(_1863_));
 sky130_fd_sc_hd__mux2_1 _4893_ (.A0(_1863_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .S(_1734_),
    .X(_1864_));
 sky130_fd_sc_hd__mux2_1 _4894_ (.A0(net530),
    .A1(_1864_),
    .S(net53),
    .X(_0204_));
 sky130_fd_sc_hd__nand2_1 _4895_ (.A(net92),
    .B(_1593_),
    .Y(_1865_));
 sky130_fd_sc_hd__and2_1 _4896_ (.A(\z80.tv80s.i_tv80_core.ACC[0] ),
    .B(_1748_),
    .X(_1866_));
 sky130_fd_sc_hd__a221o_1 _4897_ (.A1(\z80.tv80s.i_tv80_core.SP[8] ),
    .A2(net56),
    .B1(_1747_),
    .B2(_1593_),
    .C1(_1866_),
    .X(_1867_));
 sky130_fd_sc_hd__mux2_1 _4898_ (.A0(\z80.tv80s.i_tv80_core.PC[8] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .S(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(_1868_));
 sky130_fd_sc_hd__mux2_1 _4899_ (.A0(_1593_),
    .A1(_1868_),
    .S(net104),
    .X(_1869_));
 sky130_fd_sc_hd__nor2_1 _4900_ (.A(_2746_),
    .B(_1856_),
    .Y(_1870_));
 sky130_fd_sc_hd__and2_1 _4901_ (.A(_2746_),
    .B(_1856_),
    .X(_1871_));
 sky130_fd_sc_hd__nor2_1 _4902_ (.A(_1870_),
    .B(_1871_),
    .Y(_1872_));
 sky130_fd_sc_hd__mux2_1 _4903_ (.A0(\z80.tv80s.di_reg[0] ),
    .A1(_1872_),
    .S(_1753_),
    .X(_1873_));
 sky130_fd_sc_hd__a22o_1 _4904_ (.A1(net58),
    .A2(_1869_),
    .B1(_1873_),
    .B2(_1749_),
    .X(_1874_));
 sky130_fd_sc_hd__a211o_1 _4905_ (.A1(\z80.tv80s.i_tv80_core.PC[8] ),
    .A2(net57),
    .B1(_1867_),
    .C1(_1874_),
    .X(_1875_));
 sky130_fd_sc_hd__mux2_1 _4906_ (.A0(\z80.tv80s.i_tv80_core.I[0] ),
    .A1(_1875_),
    .S(net98),
    .X(_1876_));
 sky130_fd_sc_hd__a22o_1 _4907_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .A2(_1739_),
    .B1(net60),
    .B2(_1876_),
    .X(_1877_));
 sky130_fd_sc_hd__a21bo_1 _4908_ (.A1(net87),
    .A2(_1877_),
    .B1_N(_1865_),
    .X(_1878_));
 sky130_fd_sc_hd__mux2_1 _4909_ (.A0(_1878_),
    .A1(\z80.tv80s.di_reg[0] ),
    .S(_1734_),
    .X(_1879_));
 sky130_fd_sc_hd__mux2_1 _4910_ (.A0(net528),
    .A1(_1879_),
    .S(net53),
    .X(_0205_));
 sky130_fd_sc_hd__nand2_1 _4911_ (.A(net92),
    .B(_1616_),
    .Y(_1880_));
 sky130_fd_sc_hd__and2_1 _4912_ (.A(\z80.tv80s.i_tv80_core.ACC[1] ),
    .B(_1748_),
    .X(_1881_));
 sky130_fd_sc_hd__a221o_1 _4913_ (.A1(\z80.tv80s.i_tv80_core.SP[9] ),
    .A2(net56),
    .B1(_1747_),
    .B2(_1616_),
    .C1(_1881_),
    .X(_1882_));
 sky130_fd_sc_hd__mux2_1 _4914_ (.A0(\z80.tv80s.i_tv80_core.PC[9] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .S(_0446_),
    .X(_1883_));
 sky130_fd_sc_hd__or2_1 _4915_ (.A(net104),
    .B(_1616_),
    .X(_1884_));
 sky130_fd_sc_hd__o211a_1 _4916_ (.A1(_0443_),
    .A2(_1883_),
    .B1(_1884_),
    .C1(net58),
    .X(_1885_));
 sky130_fd_sc_hd__and2_1 _4917_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .B(_1870_),
    .X(_1886_));
 sky130_fd_sc_hd__nor2_1 _4918_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .B(_1870_),
    .Y(_1887_));
 sky130_fd_sc_hd__or2_1 _4919_ (.A(\z80.tv80s.di_reg[1] ),
    .B(_1753_),
    .X(_1888_));
 sky130_fd_sc_hd__o21ai_1 _4920_ (.A1(_1886_),
    .A2(_1887_),
    .B1(_1753_),
    .Y(_1889_));
 sky130_fd_sc_hd__a31o_1 _4921_ (.A1(_1749_),
    .A2(_1888_),
    .A3(_1889_),
    .B1(_1885_),
    .X(_1890_));
 sky130_fd_sc_hd__a211o_1 _4922_ (.A1(\z80.tv80s.i_tv80_core.PC[9] ),
    .A2(net57),
    .B1(_1882_),
    .C1(_1890_),
    .X(_1891_));
 sky130_fd_sc_hd__mux2_1 _4923_ (.A0(\z80.tv80s.i_tv80_core.I[1] ),
    .A1(_1891_),
    .S(net99),
    .X(_1892_));
 sky130_fd_sc_hd__a22o_1 _4924_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .A2(net64),
    .B1(net60),
    .B2(_1892_),
    .X(_1893_));
 sky130_fd_sc_hd__a21bo_1 _4925_ (.A1(net87),
    .A2(_1893_),
    .B1_N(_1880_),
    .X(_1894_));
 sky130_fd_sc_hd__mux2_1 _4926_ (.A0(_1894_),
    .A1(\z80.tv80s.di_reg[1] ),
    .S(_1734_),
    .X(_1895_));
 sky130_fd_sc_hd__mux2_1 _4927_ (.A0(net574),
    .A1(_1895_),
    .S(net53),
    .X(_0206_));
 sky130_fd_sc_hd__nand2_1 _4928_ (.A(net92),
    .B(_1629_),
    .Y(_1896_));
 sky130_fd_sc_hd__and2_1 _4929_ (.A(\z80.tv80s.i_tv80_core.ACC[2] ),
    .B(_1748_),
    .X(_1897_));
 sky130_fd_sc_hd__a221o_1 _4930_ (.A1(\z80.tv80s.i_tv80_core.SP[10] ),
    .A2(net56),
    .B1(_1747_),
    .B2(_1629_),
    .C1(_1897_),
    .X(_1898_));
 sky130_fd_sc_hd__mux2_1 _4931_ (.A0(\z80.tv80s.i_tv80_core.PC[10] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .S(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(_1899_));
 sky130_fd_sc_hd__mux2_1 _4932_ (.A0(_1629_),
    .A1(_1899_),
    .S(net104),
    .X(_1900_));
 sky130_fd_sc_hd__xor2_1 _4933_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .B(_1886_),
    .X(_1901_));
 sky130_fd_sc_hd__mux2_1 _4934_ (.A0(\z80.tv80s.di_reg[2] ),
    .A1(_1901_),
    .S(_1753_),
    .X(_1902_));
 sky130_fd_sc_hd__a22o_1 _4935_ (.A1(net58),
    .A2(_1900_),
    .B1(_1902_),
    .B2(_1749_),
    .X(_1903_));
 sky130_fd_sc_hd__a211o_1 _4936_ (.A1(\z80.tv80s.i_tv80_core.PC[10] ),
    .A2(net57),
    .B1(_1898_),
    .C1(_1903_),
    .X(_1904_));
 sky130_fd_sc_hd__mux2_1 _4937_ (.A0(\z80.tv80s.i_tv80_core.I[2] ),
    .A1(_1904_),
    .S(net99),
    .X(_1905_));
 sky130_fd_sc_hd__a22oi_1 _4938_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .A2(net64),
    .B1(net60),
    .B2(_1905_),
    .Y(_1906_));
 sky130_fd_sc_hd__o21a_1 _4939_ (.A1(net92),
    .A2(_1906_),
    .B1(_1896_),
    .X(_1907_));
 sky130_fd_sc_hd__nand2_1 _4940_ (.A(\z80.tv80s.di_reg[2] ),
    .B(net68),
    .Y(_1908_));
 sky130_fd_sc_hd__o21ai_2 _4941_ (.A1(net68),
    .A2(_1907_),
    .B1(_1908_),
    .Y(_1909_));
 sky130_fd_sc_hd__mux2_1 _4942_ (.A0(net613),
    .A1(_1909_),
    .S(_1389_),
    .X(_0207_));
 sky130_fd_sc_hd__nand2_1 _4943_ (.A(net92),
    .B(_1644_),
    .Y(_1910_));
 sky130_fd_sc_hd__and2_1 _4944_ (.A(\z80.tv80s.i_tv80_core.ACC[3] ),
    .B(_1748_),
    .X(_1911_));
 sky130_fd_sc_hd__a221o_1 _4945_ (.A1(\z80.tv80s.i_tv80_core.SP[11] ),
    .A2(net56),
    .B1(_1747_),
    .B2(_1644_),
    .C1(_1911_),
    .X(_1912_));
 sky130_fd_sc_hd__mux2_1 _4946_ (.A0(\z80.tv80s.i_tv80_core.PC[11] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .S(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(_1913_));
 sky130_fd_sc_hd__mux2_1 _4947_ (.A0(_1644_),
    .A1(_1913_),
    .S(net104),
    .X(_1914_));
 sky130_fd_sc_hd__and3_1 _4948_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .C(_1886_),
    .X(_1915_));
 sky130_fd_sc_hd__a21oi_1 _4949_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .A2(_1886_),
    .B1(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .Y(_1916_));
 sky130_fd_sc_hd__nor2_1 _4950_ (.A(_1915_),
    .B(_1916_),
    .Y(_1917_));
 sky130_fd_sc_hd__mux2_1 _4951_ (.A0(\z80.tv80s.di_reg[3] ),
    .A1(_1917_),
    .S(_1753_),
    .X(_1918_));
 sky130_fd_sc_hd__a22o_1 _4952_ (.A1(net58),
    .A2(_1914_),
    .B1(_1918_),
    .B2(_1749_),
    .X(_1919_));
 sky130_fd_sc_hd__a211o_1 _4953_ (.A1(\z80.tv80s.i_tv80_core.PC[11] ),
    .A2(net57),
    .B1(_1912_),
    .C1(_1919_),
    .X(_1920_));
 sky130_fd_sc_hd__mux2_1 _4954_ (.A0(\z80.tv80s.i_tv80_core.I[3] ),
    .A1(_1920_),
    .S(net99),
    .X(_1921_));
 sky130_fd_sc_hd__a22o_1 _4955_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .A2(net64),
    .B1(net60),
    .B2(_1921_),
    .X(_1922_));
 sky130_fd_sc_hd__a21bo_1 _4956_ (.A1(net87),
    .A2(_1922_),
    .B1_N(_1910_),
    .X(_1923_));
 sky130_fd_sc_hd__mux2_1 _4957_ (.A0(_1923_),
    .A1(\z80.tv80s.di_reg[3] ),
    .S(net68),
    .X(_1924_));
 sky130_fd_sc_hd__mux2_1 _4958_ (.A0(net560),
    .A1(_1924_),
    .S(_1389_),
    .X(_0208_));
 sky130_fd_sc_hd__nand2_1 _4959_ (.A(net92),
    .B(_1657_),
    .Y(_1925_));
 sky130_fd_sc_hd__and2_1 _4960_ (.A(\z80.tv80s.i_tv80_core.ACC[4] ),
    .B(_1748_),
    .X(_1926_));
 sky130_fd_sc_hd__a221o_1 _4961_ (.A1(\z80.tv80s.i_tv80_core.SP[12] ),
    .A2(net56),
    .B1(_1747_),
    .B2(_1657_),
    .C1(_1926_),
    .X(_1927_));
 sky130_fd_sc_hd__mux2_1 _4962_ (.A0(\z80.tv80s.i_tv80_core.PC[12] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .S(_0446_),
    .X(_1928_));
 sky130_fd_sc_hd__or2_1 _4963_ (.A(net104),
    .B(_1657_),
    .X(_1929_));
 sky130_fd_sc_hd__o211a_1 _4964_ (.A1(_0443_),
    .A2(_1928_),
    .B1(_1929_),
    .C1(net58),
    .X(_1930_));
 sky130_fd_sc_hd__and2_1 _4965_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .B(_1915_),
    .X(_1931_));
 sky130_fd_sc_hd__nor2_1 _4966_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .B(_1915_),
    .Y(_1932_));
 sky130_fd_sc_hd__or2_1 _4967_ (.A(\z80.tv80s.di_reg[4] ),
    .B(_1753_),
    .X(_1933_));
 sky130_fd_sc_hd__o21ai_1 _4968_ (.A1(_1931_),
    .A2(_1932_),
    .B1(_1753_),
    .Y(_1934_));
 sky130_fd_sc_hd__a31o_1 _4969_ (.A1(_1749_),
    .A2(_1933_),
    .A3(_1934_),
    .B1(_1930_),
    .X(_1935_));
 sky130_fd_sc_hd__a211o_1 _4970_ (.A1(\z80.tv80s.i_tv80_core.PC[12] ),
    .A2(net57),
    .B1(_1927_),
    .C1(_1935_),
    .X(_1936_));
 sky130_fd_sc_hd__mux2_1 _4971_ (.A0(\z80.tv80s.i_tv80_core.I[4] ),
    .A1(_1936_),
    .S(net99),
    .X(_1937_));
 sky130_fd_sc_hd__a22o_1 _4972_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .A2(net64),
    .B1(net60),
    .B2(_1937_),
    .X(_1938_));
 sky130_fd_sc_hd__a21bo_1 _4973_ (.A1(net87),
    .A2(_1938_),
    .B1_N(_1925_),
    .X(_1939_));
 sky130_fd_sc_hd__mux2_1 _4974_ (.A0(_1939_),
    .A1(\z80.tv80s.di_reg[4] ),
    .S(net68),
    .X(_1940_));
 sky130_fd_sc_hd__mux2_1 _4975_ (.A0(net582),
    .A1(_1940_),
    .S(_1389_),
    .X(_0209_));
 sky130_fd_sc_hd__nand2_1 _4976_ (.A(net92),
    .B(_1671_),
    .Y(_1941_));
 sky130_fd_sc_hd__and2_1 _4977_ (.A(\z80.tv80s.i_tv80_core.ACC[5] ),
    .B(_1748_),
    .X(_1942_));
 sky130_fd_sc_hd__a221o_1 _4978_ (.A1(\z80.tv80s.i_tv80_core.SP[13] ),
    .A2(net56),
    .B1(_1747_),
    .B2(_1671_),
    .C1(_1942_),
    .X(_1943_));
 sky130_fd_sc_hd__mux2_1 _4979_ (.A0(\z80.tv80s.i_tv80_core.PC[13] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .S(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(_1944_));
 sky130_fd_sc_hd__mux2_1 _4980_ (.A0(_1671_),
    .A1(_1944_),
    .S(_0444_),
    .X(_1945_));
 sky130_fd_sc_hd__xor2_1 _4981_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .B(_1931_),
    .X(_1946_));
 sky130_fd_sc_hd__mux2_1 _4982_ (.A0(\z80.tv80s.di_reg[5] ),
    .A1(_1946_),
    .S(_1753_),
    .X(_1947_));
 sky130_fd_sc_hd__a22o_1 _4983_ (.A1(net58),
    .A2(_1945_),
    .B1(_1947_),
    .B2(_1749_),
    .X(_1948_));
 sky130_fd_sc_hd__a211o_1 _4984_ (.A1(\z80.tv80s.i_tv80_core.PC[13] ),
    .A2(net57),
    .B1(_1943_),
    .C1(_1948_),
    .X(_1949_));
 sky130_fd_sc_hd__mux2_1 _4985_ (.A0(\z80.tv80s.i_tv80_core.I[5] ),
    .A1(_1949_),
    .S(net99),
    .X(_1950_));
 sky130_fd_sc_hd__a22o_1 _4986_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .A2(net64),
    .B1(net60),
    .B2(_1950_),
    .X(_1951_));
 sky130_fd_sc_hd__a21bo_1 _4987_ (.A1(net87),
    .A2(_1951_),
    .B1_N(_1941_),
    .X(_1952_));
 sky130_fd_sc_hd__mux2_1 _4988_ (.A0(_1952_),
    .A1(\z80.tv80s.di_reg[5] ),
    .S(net68),
    .X(_1953_));
 sky130_fd_sc_hd__mux2_1 _4989_ (.A0(net556),
    .A1(_1953_),
    .S(_1389_),
    .X(_0210_));
 sky130_fd_sc_hd__nand2_1 _4990_ (.A(net92),
    .B(_1682_),
    .Y(_1954_));
 sky130_fd_sc_hd__and2_1 _4991_ (.A(\z80.tv80s.i_tv80_core.ACC[6] ),
    .B(_1748_),
    .X(_1955_));
 sky130_fd_sc_hd__a221o_1 _4992_ (.A1(\z80.tv80s.i_tv80_core.SP[14] ),
    .A2(net56),
    .B1(_1747_),
    .B2(_1682_),
    .C1(_1955_),
    .X(_1956_));
 sky130_fd_sc_hd__mux2_1 _4993_ (.A0(\z80.tv80s.i_tv80_core.PC[14] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .S(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(_1957_));
 sky130_fd_sc_hd__mux2_1 _4994_ (.A0(_1682_),
    .A1(_1957_),
    .S(_0444_),
    .X(_1958_));
 sky130_fd_sc_hd__and3_1 _4995_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .C(_1931_),
    .X(_1959_));
 sky130_fd_sc_hd__a21oi_1 _4996_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .A2(_1931_),
    .B1(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .Y(_1960_));
 sky130_fd_sc_hd__nor2_1 _4997_ (.A(_1959_),
    .B(_1960_),
    .Y(_1961_));
 sky130_fd_sc_hd__mux2_1 _4998_ (.A0(\z80.tv80s.di_reg[6] ),
    .A1(_1961_),
    .S(_1753_),
    .X(_1962_));
 sky130_fd_sc_hd__a22o_1 _4999_ (.A1(net58),
    .A2(_1958_),
    .B1(_1962_),
    .B2(_1749_),
    .X(_1963_));
 sky130_fd_sc_hd__a211o_1 _5000_ (.A1(\z80.tv80s.i_tv80_core.PC[14] ),
    .A2(_1744_),
    .B1(_1956_),
    .C1(_1963_),
    .X(_1964_));
 sky130_fd_sc_hd__mux2_1 _5001_ (.A0(net549),
    .A1(_1964_),
    .S(net99),
    .X(_1965_));
 sky130_fd_sc_hd__a22oi_1 _5002_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .A2(net64),
    .B1(net60),
    .B2(_1965_),
    .Y(_1966_));
 sky130_fd_sc_hd__o21a_1 _5003_ (.A1(_1238_),
    .A2(_1966_),
    .B1(_1954_),
    .X(_1967_));
 sky130_fd_sc_hd__nand2_1 _5004_ (.A(\z80.tv80s.di_reg[6] ),
    .B(net68),
    .Y(_1968_));
 sky130_fd_sc_hd__o21ai_2 _5005_ (.A1(net68),
    .A2(_1967_),
    .B1(_1968_),
    .Y(_1969_));
 sky130_fd_sc_hd__mux2_1 _5006_ (.A0(net562),
    .A1(_1969_),
    .S(_1389_),
    .X(_0211_));
 sky130_fd_sc_hd__nand2_1 _5007_ (.A(_1238_),
    .B(_1697_),
    .Y(_1970_));
 sky130_fd_sc_hd__and2_1 _5008_ (.A(\z80.tv80s.i_tv80_core.ACC[7] ),
    .B(_1748_),
    .X(_1971_));
 sky130_fd_sc_hd__a221o_1 _5009_ (.A1(\z80.tv80s.i_tv80_core.SP[15] ),
    .A2(net56),
    .B1(_1747_),
    .B2(_1697_),
    .C1(_1971_),
    .X(_1972_));
 sky130_fd_sc_hd__mux2_1 _5010_ (.A0(\z80.tv80s.i_tv80_core.PC[15] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[15] ),
    .S(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(_1973_));
 sky130_fd_sc_hd__mux2_1 _5011_ (.A0(_1697_),
    .A1(_1973_),
    .S(_0444_),
    .X(_1974_));
 sky130_fd_sc_hd__xor2_1 _5012_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[15] ),
    .B(_1959_),
    .X(_1975_));
 sky130_fd_sc_hd__mux2_1 _5013_ (.A0(\z80.tv80s.di_reg[7] ),
    .A1(_1975_),
    .S(_1753_),
    .X(_1976_));
 sky130_fd_sc_hd__a22o_1 _5014_ (.A1(_0441_),
    .A2(_1974_),
    .B1(_1976_),
    .B2(_1749_),
    .X(_1977_));
 sky130_fd_sc_hd__a211o_1 _5015_ (.A1(\z80.tv80s.i_tv80_core.PC[15] ),
    .A2(_1744_),
    .B1(_1972_),
    .C1(_1977_),
    .X(_1978_));
 sky130_fd_sc_hd__mux2_1 _5016_ (.A0(\z80.tv80s.i_tv80_core.I[7] ),
    .A1(_1978_),
    .S(net99),
    .X(_1979_));
 sky130_fd_sc_hd__a22o_1 _5017_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[15] ),
    .A2(net64),
    .B1(net60),
    .B2(_1979_),
    .X(_1980_));
 sky130_fd_sc_hd__a21bo_1 _5018_ (.A1(net87),
    .A2(_1980_),
    .B1_N(_1970_),
    .X(_1981_));
 sky130_fd_sc_hd__mux2_1 _5019_ (.A0(_1981_),
    .A1(\z80.tv80s.di_reg[7] ),
    .S(net68),
    .X(_1982_));
 sky130_fd_sc_hd__mux2_1 _5020_ (.A0(net536),
    .A1(_1982_),
    .S(_1389_),
    .X(_0212_));
 sky130_fd_sc_hd__and3b_2 _5021_ (.A_N(_0692_),
    .B(_0705_),
    .C(_0714_),
    .X(_1983_));
 sky130_fd_sc_hd__o21ba_1 _5022_ (.A1(_2719_),
    .A2(_0642_),
    .B1_N(_1983_),
    .X(_1984_));
 sky130_fd_sc_hd__or2_1 _5023_ (.A(net157),
    .B(_1984_),
    .X(_1985_));
 sky130_fd_sc_hd__or2_1 _5024_ (.A(net108),
    .B(_0764_),
    .X(_1986_));
 sky130_fd_sc_hd__nor2_2 _5025_ (.A(_2722_),
    .B(_1986_),
    .Y(_1987_));
 sky130_fd_sc_hd__inv_2 _5026_ (.A(_1987_),
    .Y(_1988_));
 sky130_fd_sc_hd__a211o_1 _5027_ (.A1(_2711_),
    .A2(\z80.tv80s.i_tv80_core.Z16_r ),
    .B1(_0781_),
    .C1(_0828_),
    .X(_1989_));
 sky130_fd_sc_hd__or3b_1 _5028_ (.A(_1989_),
    .B(_0951_),
    .C_N(_0907_),
    .X(_1990_));
 sky130_fd_sc_hd__or3_1 _5029_ (.A(_0995_),
    .B(_1038_),
    .C(_1990_),
    .X(_1991_));
 sky130_fd_sc_hd__o31a_1 _5030_ (.A1(_1074_),
    .A2(_1136_),
    .A3(_1991_),
    .B1(_2731_),
    .X(_1992_));
 sky130_fd_sc_hd__a211o_1 _5031_ (.A1(_2711_),
    .A2(\z80.tv80s.i_tv80_core.Arith16_r ),
    .B1(_1992_),
    .C1(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .X(_1993_));
 sky130_fd_sc_hd__nand2_1 _5032_ (.A(_0975_),
    .B(_1051_),
    .Y(_1994_));
 sky130_fd_sc_hd__or3b_1 _5033_ (.A(_0790_),
    .B(_0910_),
    .C_N(_0957_),
    .X(_1995_));
 sky130_fd_sc_hd__or4b_1 _5034_ (.A(\z80.tv80s.i_tv80_core.BusA[0] ),
    .B(_1994_),
    .C(_1995_),
    .D_N(_0840_),
    .X(_1996_));
 sky130_fd_sc_hd__or4_1 _5035_ (.A(_0912_),
    .B(_0959_),
    .C(_0979_),
    .D(_1053_),
    .X(_1997_));
 sky130_fd_sc_hd__or3_1 _5036_ (.A(_0793_),
    .B(_0830_),
    .C(_1997_),
    .X(_1998_));
 sky130_fd_sc_hd__o31a_1 _5037_ (.A1(_1084_),
    .A2(_1156_),
    .A3(_1998_),
    .B1(net115),
    .X(_1999_));
 sky130_fd_sc_hd__o21ai_1 _5038_ (.A1(net115),
    .A2(\z80.tv80s.i_tv80_core.F[6] ),
    .B1(_0791_),
    .Y(_2000_));
 sky130_fd_sc_hd__or2_1 _5039_ (.A(_1999_),
    .B(_2000_),
    .X(_2001_));
 sky130_fd_sc_hd__a22o_1 _5040_ (.A1(\z80.tv80s.i_tv80_core.BusB[3] ),
    .A2(_0581_),
    .B1(_0832_),
    .B2(\z80.tv80s.i_tv80_core.BusB[1] ),
    .X(_2002_));
 sky130_fd_sc_hd__a21o_1 _5041_ (.A1(\z80.tv80s.i_tv80_core.BusB[0] ),
    .A2(_0782_),
    .B1(_2002_),
    .X(_2003_));
 sky130_fd_sc_hd__a22o_1 _5042_ (.A1(\z80.tv80s.i_tv80_core.BusB[6] ),
    .A2(_2891_),
    .B1(_0411_),
    .B2(\z80.tv80s.i_tv80_core.BusB[5] ),
    .X(_2004_));
 sky130_fd_sc_hd__a221o_1 _5043_ (.A1(\z80.tv80s.i_tv80_core.BusB[4] ),
    .A2(_0409_),
    .B1(_0914_),
    .B2(\z80.tv80s.i_tv80_core.BusB[2] ),
    .C1(_2004_),
    .X(_2005_));
 sky130_fd_sc_hd__or4b_1 _5044_ (.A(_1149_),
    .B(_2003_),
    .C(_2005_),
    .D_N(_0785_),
    .X(_2006_));
 sky130_fd_sc_hd__or4_1 _5045_ (.A(_0788_),
    .B(_0829_),
    .C(_0911_),
    .D(_0958_),
    .X(_2007_));
 sky130_fd_sc_hd__or4_1 _5046_ (.A(net139),
    .B(\z80.tv80s.i_tv80_core.BusA[4] ),
    .C(\z80.tv80s.i_tv80_core.BusA[5] ),
    .D(\z80.tv80s.i_tv80_core.BusA[6] ),
    .X(_2008_));
 sky130_fd_sc_hd__o311a_1 _5047_ (.A1(_0787_),
    .A2(_2007_),
    .A3(_2008_),
    .B1(_1988_),
    .C1(_2006_),
    .X(_2009_));
 sky130_fd_sc_hd__o31a_1 _5048_ (.A1(_1082_),
    .A2(_1148_),
    .A3(_1996_),
    .B1(_2009_),
    .X(_2010_));
 sky130_fd_sc_hd__a32o_1 _5049_ (.A1(_1993_),
    .A2(_2001_),
    .A3(_2010_),
    .B1(_1987_),
    .B2(_2711_),
    .X(_2011_));
 sky130_fd_sc_hd__and2b_1 _5050_ (.A_N(_1983_),
    .B(_2011_),
    .X(_2012_));
 sky130_fd_sc_hd__or2_1 _5051_ (.A(_1985_),
    .B(_2012_),
    .X(_2013_));
 sky130_fd_sc_hd__and4_1 _5052_ (.A(_0871_),
    .B(_0894_),
    .C(_0938_),
    .D(_1983_),
    .X(_2014_));
 sky130_fd_sc_hd__and4_1 _5053_ (.A(_1011_),
    .B(_1026_),
    .C(_1108_),
    .D(_2014_),
    .X(_2015_));
 sky130_fd_sc_hd__and4_1 _5054_ (.A(_1124_),
    .B(_1266_),
    .C(_1279_),
    .D(_2015_),
    .X(_2016_));
 sky130_fd_sc_hd__and4_1 _5055_ (.A(_1293_),
    .B(_1305_),
    .C(_1322_),
    .D(_2016_),
    .X(_2017_));
 sky130_fd_sc_hd__a41o_1 _5056_ (.A1(_1336_),
    .A2(_1351_),
    .A3(_1363_),
    .A4(_2017_),
    .B1(_2013_),
    .X(_2018_));
 sky130_fd_sc_hd__a21bo_1 _5057_ (.A1(net485),
    .A2(_1985_),
    .B1_N(_2018_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _5058_ (.A0(_2748_),
    .A1(_0760_),
    .S(net109),
    .X(_2019_));
 sky130_fd_sc_hd__inv_2 _5059_ (.A(_2019_),
    .Y(_0214_));
 sky130_fd_sc_hd__mux2_1 _5060_ (.A0(net228),
    .A1(_0867_),
    .S(net109),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _5061_ (.A0(net224),
    .A1(_0892_),
    .S(net109),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _5062_ (.A0(net236),
    .A1(_0933_),
    .S(net111),
    .X(_0217_));
 sky130_fd_sc_hd__mux2_1 _5063_ (.A0(net230),
    .A1(_1008_),
    .S(net111),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _5064_ (.A0(net234),
    .A1(_1022_),
    .S(net111),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _5065_ (.A0(net218),
    .A1(_1102_),
    .S(net109),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _5066_ (.A0(net220),
    .A1(_1121_),
    .S(net109),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _5067_ (.A0(net238),
    .A1(_1262_),
    .S(net111),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _5068_ (.A0(net253),
    .A1(_1275_),
    .S(net111),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_1 _5069_ (.A0(net232),
    .A1(_1288_),
    .S(net111),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _5070_ (.A0(net226),
    .A1(_1302_),
    .S(net111),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _5071_ (.A0(net246),
    .A1(_1318_),
    .S(net114),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _5072_ (.A0(net248),
    .A1(_1331_),
    .S(net114),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _5073_ (.A0(net222),
    .A1(_1346_),
    .S(net111),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _5074_ (.A0(net242),
    .A1(_1361_),
    .S(net114),
    .X(_0229_));
 sky130_fd_sc_hd__o21ai_1 _5075_ (.A1(_0406_),
    .A2(_1240_),
    .B1(_1241_),
    .Y(_2020_));
 sky130_fd_sc_hd__mux2_1 _5076_ (.A0(net153),
    .A1(_2020_),
    .S(net109),
    .X(_0230_));
 sky130_fd_sc_hd__a221o_1 _5077_ (.A1(_2829_),
    .A2(_2936_),
    .B1(_0612_),
    .B2(_2805_),
    .C1(_1208_),
    .X(_2021_));
 sky130_fd_sc_hd__or3_1 _5078_ (.A(_0681_),
    .B(_0683_),
    .C(_2021_),
    .X(_2022_));
 sky130_fd_sc_hd__a21oi_1 _5079_ (.A1(_2925_),
    .A2(_1415_),
    .B1(_2022_),
    .Y(_2023_));
 sky130_fd_sc_hd__nor2_1 _5080_ (.A(net115),
    .B(_2023_),
    .Y(_2024_));
 sky130_fd_sc_hd__a31o_1 _5081_ (.A1(net149),
    .A2(_2890_),
    .A3(_2891_),
    .B1(net105),
    .X(_2025_));
 sky130_fd_sc_hd__a22o_1 _5082_ (.A1(net148),
    .A2(_2844_),
    .B1(_1217_),
    .B2(_2805_),
    .X(_2026_));
 sky130_fd_sc_hd__o221a_4 _5083_ (.A1(net107),
    .A2(_2024_),
    .B1(_2025_),
    .B2(_2026_),
    .C1(_2697_),
    .X(_2027_));
 sky130_fd_sc_hd__inv_2 _5084_ (.A(_2027_),
    .Y(_2028_));
 sky130_fd_sc_hd__nand2_1 _5085_ (.A(_1233_),
    .B(_2027_),
    .Y(_2029_));
 sky130_fd_sc_hd__a31oi_4 _5086_ (.A1(_1221_),
    .A2(_1233_),
    .A3(_2027_),
    .B1(net157),
    .Y(_2030_));
 sky130_fd_sc_hd__or2_2 _5087_ (.A(_1233_),
    .B(_2028_),
    .X(_2031_));
 sky130_fd_sc_hd__inv_2 _5088_ (.A(_2031_),
    .Y(_2032_));
 sky130_fd_sc_hd__a31o_1 _5089_ (.A1(net164),
    .A2(net96),
    .A3(_1215_),
    .B1(_1207_),
    .X(_2033_));
 sky130_fd_sc_hd__o211a_1 _5090_ (.A1(net144),
    .A2(_1402_),
    .B1(_1394_),
    .C1(_0590_),
    .X(_2034_));
 sky130_fd_sc_hd__a32o_1 _5091_ (.A1(net126),
    .A2(net148),
    .A3(_2890_),
    .B1(_1395_),
    .B2(_2856_),
    .X(_2035_));
 sky130_fd_sc_hd__o31a_1 _5092_ (.A1(_1187_),
    .A2(_2034_),
    .A3(_2035_),
    .B1(net107),
    .X(_2036_));
 sky130_fd_sc_hd__nor2_1 _5093_ (.A(_2942_),
    .B(_0415_),
    .Y(_2037_));
 sky130_fd_sc_hd__o31a_1 _5094_ (.A1(_0398_),
    .A2(_0593_),
    .A3(_2037_),
    .B1(_0396_),
    .X(_2038_));
 sky130_fd_sc_hd__o211a_1 _5095_ (.A1(net116),
    .A2(_2805_),
    .B1(_2925_),
    .C1(_2936_),
    .X(_2039_));
 sky130_fd_sc_hd__a221o_1 _5096_ (.A1(_2885_),
    .A2(_0430_),
    .B1(_1395_),
    .B2(_2920_),
    .C1(_2039_),
    .X(_2040_));
 sky130_fd_sc_hd__a221o_1 _5097_ (.A1(net146),
    .A2(_2769_),
    .B1(_2834_),
    .B2(net135),
    .C1(_2040_),
    .X(_2041_));
 sky130_fd_sc_hd__a211o_1 _5098_ (.A1(_2768_),
    .A2(_0423_),
    .B1(_0599_),
    .C1(_2829_),
    .X(_2042_));
 sky130_fd_sc_hd__a211o_1 _5099_ (.A1(net149),
    .A2(_2042_),
    .B1(_2041_),
    .C1(_2038_),
    .X(_2043_));
 sky130_fd_sc_hd__a21oi_1 _5100_ (.A1(net164),
    .A2(_2043_),
    .B1(_2036_),
    .Y(_2044_));
 sky130_fd_sc_hd__o2bb2a_4 _5101_ (.A1_N(net135),
    .A2_N(_2033_),
    .B1(_2044_),
    .B2(net142),
    .X(_2045_));
 sky130_fd_sc_hd__inv_2 _5102_ (.A(_2045_),
    .Y(_2046_));
 sky130_fd_sc_hd__nand2_1 _5103_ (.A(_1221_),
    .B(_2046_),
    .Y(_2047_));
 sky130_fd_sc_hd__nor2_2 _5104_ (.A(_2031_),
    .B(_2047_),
    .Y(_2048_));
 sky130_fd_sc_hd__or2_1 _5105_ (.A(_1221_),
    .B(_2046_),
    .X(_2049_));
 sky130_fd_sc_hd__nor2_2 _5106_ (.A(_2031_),
    .B(_2049_),
    .Y(_2050_));
 sky130_fd_sc_hd__nand2_1 _5107_ (.A(_1233_),
    .B(_2028_),
    .Y(_2051_));
 sky130_fd_sc_hd__nor2_2 _5108_ (.A(_2047_),
    .B(_2051_),
    .Y(_2052_));
 sky130_fd_sc_hd__a21oi_4 _5109_ (.A1(_1221_),
    .A2(_1233_),
    .B1(_2027_),
    .Y(_2053_));
 sky130_fd_sc_hd__a221o_1 _5110_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ),
    .A2(net140),
    .B1(net82),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ),
    .C1(net81),
    .X(_2054_));
 sky130_fd_sc_hd__a221o_1 _5111_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ),
    .A2(net140),
    .B1(net82),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ),
    .C1(net79),
    .X(_2055_));
 sky130_fd_sc_hd__a221o_1 _5112_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ),
    .A2(net141),
    .B1(net83),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ),
    .C1(net80),
    .X(_2056_));
 sky130_fd_sc_hd__a221o_1 _5113_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ),
    .A2(net141),
    .B1(net83),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ),
    .C1(net79),
    .X(_2057_));
 sky130_fd_sc_hd__and3_1 _5114_ (.A(_0808_),
    .B(_2054_),
    .C(_2055_),
    .X(_2058_));
 sky130_fd_sc_hd__a211o_1 _5115_ (.A1(_0734_),
    .A2(_0809_),
    .B1(_2045_),
    .C1(_2058_),
    .X(_2059_));
 sky130_fd_sc_hd__and3_1 _5116_ (.A(_0808_),
    .B(_2056_),
    .C(_2057_),
    .X(_2060_));
 sky130_fd_sc_hd__a211o_1 _5117_ (.A1(_0809_),
    .A2(_1252_),
    .B1(_2046_),
    .C1(_2060_),
    .X(_2061_));
 sky130_fd_sc_hd__or2_1 _5118_ (.A(_1221_),
    .B(_2045_),
    .X(_2062_));
 sky130_fd_sc_hd__nor2_2 _5119_ (.A(_2029_),
    .B(_2062_),
    .Y(_2063_));
 sky130_fd_sc_hd__nand2_1 _5120_ (.A(_1221_),
    .B(_2045_),
    .Y(_2064_));
 sky130_fd_sc_hd__nor2_2 _5121_ (.A(_2051_),
    .B(_2064_),
    .Y(_2065_));
 sky130_fd_sc_hd__nor2_2 _5122_ (.A(_2029_),
    .B(_2049_),
    .Y(_2066_));
 sky130_fd_sc_hd__o21ai_1 _5123_ (.A1(_2747_),
    .A2(_2062_),
    .B1(_2064_),
    .Y(_2067_));
 sky130_fd_sc_hd__a32o_1 _5124_ (.A1(_2053_),
    .A2(_2059_),
    .A3(_2061_),
    .B1(_2050_),
    .B2(\z80.tv80s.i_tv80_core.SP[0] ),
    .X(_2068_));
 sky130_fd_sc_hd__a221o_1 _5125_ (.A1(\z80.tv80s.i_tv80_core.F[0] ),
    .A2(_2048_),
    .B1(_2052_),
    .B2(\z80.tv80s.i_tv80_core.ACC[0] ),
    .C1(_2068_),
    .X(_2069_));
 sky130_fd_sc_hd__a221o_1 _5126_ (.A1(\z80.tv80s.di_reg[0] ),
    .A2(_2065_),
    .B1(_2067_),
    .B2(_2032_),
    .C1(_2069_),
    .X(_2070_));
 sky130_fd_sc_hd__a221o_1 _5127_ (.A1(\z80.tv80s.i_tv80_core.PC[8] ),
    .A2(_2063_),
    .B1(_2066_),
    .B2(\z80.tv80s.i_tv80_core.PC[0] ),
    .C1(_2070_),
    .X(_2071_));
 sky130_fd_sc_hd__a22o_1 _5128_ (.A1(net160),
    .A2(net580),
    .B1(_2030_),
    .B2(_2071_),
    .X(_0231_));
 sky130_fd_sc_hd__nor2_2 _5129_ (.A(_2031_),
    .B(_2062_),
    .Y(_2072_));
 sky130_fd_sc_hd__a22o_1 _5130_ (.A1(\z80.tv80s.i_tv80_core.ACC[1] ),
    .A2(_2052_),
    .B1(_2072_),
    .B2(\z80.tv80s.i_tv80_core.SP[9] ),
    .X(_2073_));
 sky130_fd_sc_hd__a221o_1 _5131_ (.A1(\z80.tv80s.i_tv80_core.SP[1] ),
    .A2(_2050_),
    .B1(_2066_),
    .B2(\z80.tv80s.i_tv80_core.PC[1] ),
    .C1(_2073_),
    .X(_2074_));
 sky130_fd_sc_hd__o221a_1 _5132_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ),
    .A2(net141),
    .B1(net83),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ),
    .C1(net79),
    .X(_2075_));
 sky130_fd_sc_hd__o221a_1 _5133_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ),
    .A2(net141),
    .B1(net83),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ),
    .C1(net80),
    .X(_2076_));
 sky130_fd_sc_hd__or3_1 _5134_ (.A(_0809_),
    .B(_2075_),
    .C(_2076_),
    .X(_2077_));
 sky130_fd_sc_hd__o211a_1 _5135_ (.A1(_0808_),
    .A2(_1282_),
    .B1(_2045_),
    .C1(_2077_),
    .X(_2078_));
 sky130_fd_sc_hd__a21o_1 _5136_ (.A1(_0816_),
    .A2(_2046_),
    .B1(_2078_),
    .X(_2079_));
 sky130_fd_sc_hd__a22o_1 _5137_ (.A1(\z80.tv80s.i_tv80_core.F[1] ),
    .A2(_2048_),
    .B1(_2053_),
    .B2(_2079_),
    .X(_2080_));
 sky130_fd_sc_hd__a221o_1 _5138_ (.A1(\z80.tv80s.i_tv80_core.PC[9] ),
    .A2(_2063_),
    .B1(_2065_),
    .B2(\z80.tv80s.di_reg[1] ),
    .C1(_2080_),
    .X(_2081_));
 sky130_fd_sc_hd__or2_1 _5139_ (.A(_2074_),
    .B(_2081_),
    .X(_2082_));
 sky130_fd_sc_hd__a22o_1 _5140_ (.A1(net160),
    .A2(net701),
    .B1(_2030_),
    .B2(_2082_),
    .X(_0232_));
 sky130_fd_sc_hd__a22o_1 _5141_ (.A1(\z80.tv80s.i_tv80_core.SP[2] ),
    .A2(_2050_),
    .B1(_2066_),
    .B2(net609),
    .X(_2083_));
 sky130_fd_sc_hd__o221a_1 _5142_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ),
    .A2(net141),
    .B1(net83),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ),
    .C1(net79),
    .X(_2084_));
 sky130_fd_sc_hd__o221a_1 _5143_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ),
    .A2(net141),
    .B1(net83),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ),
    .C1(net80),
    .X(_2085_));
 sky130_fd_sc_hd__or3_1 _5144_ (.A(_0809_),
    .B(_2084_),
    .C(_2085_),
    .X(_2086_));
 sky130_fd_sc_hd__o211a_1 _5145_ (.A1(_0808_),
    .A2(_1296_),
    .B1(_2045_),
    .C1(_2086_),
    .X(_2087_));
 sky130_fd_sc_hd__a21o_1 _5146_ (.A1(_0882_),
    .A2(_2046_),
    .B1(_2087_),
    .X(_2088_));
 sky130_fd_sc_hd__a22o_1 _5147_ (.A1(\z80.tv80s.i_tv80_core.F[2] ),
    .A2(_2048_),
    .B1(_2065_),
    .B2(\z80.tv80s.di_reg[2] ),
    .X(_2089_));
 sky130_fd_sc_hd__a22o_1 _5148_ (.A1(\z80.tv80s.i_tv80_core.PC[10] ),
    .A2(_2063_),
    .B1(_2088_),
    .B2(_2053_),
    .X(_2090_));
 sky130_fd_sc_hd__a221o_1 _5149_ (.A1(\z80.tv80s.i_tv80_core.ACC[2] ),
    .A2(_2052_),
    .B1(_2072_),
    .B2(\z80.tv80s.i_tv80_core.SP[10] ),
    .C1(_2090_),
    .X(_2091_));
 sky130_fd_sc_hd__or3_1 _5150_ (.A(_2083_),
    .B(_2089_),
    .C(_2091_),
    .X(_2092_));
 sky130_fd_sc_hd__a22o_1 _5151_ (.A1(net157),
    .A2(net652),
    .B1(_2030_),
    .B2(_2092_),
    .X(_0233_));
 sky130_fd_sc_hd__a22o_1 _5152_ (.A1(\z80.tv80s.di_reg[3] ),
    .A2(_2065_),
    .B1(_2066_),
    .B2(\z80.tv80s.i_tv80_core.PC[3] ),
    .X(_2093_));
 sky130_fd_sc_hd__a22o_1 _5153_ (.A1(\z80.tv80s.i_tv80_core.SP[3] ),
    .A2(_2050_),
    .B1(_2072_),
    .B2(\z80.tv80s.i_tv80_core.SP[11] ),
    .X(_2094_));
 sky130_fd_sc_hd__a22o_1 _5154_ (.A1(net621),
    .A2(_2048_),
    .B1(_2063_),
    .B2(\z80.tv80s.i_tv80_core.PC[11] ),
    .X(_2095_));
 sky130_fd_sc_hd__o221a_1 _5155_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ),
    .A2(net140),
    .B1(net82),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ),
    .C1(net79),
    .X(_2096_));
 sky130_fd_sc_hd__o221a_1 _5156_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ),
    .A2(net140),
    .B1(net85),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][3] ),
    .C1(net81),
    .X(_2097_));
 sky130_fd_sc_hd__or2_1 _5157_ (.A(_2096_),
    .B(_2097_),
    .X(_2098_));
 sky130_fd_sc_hd__o221a_1 _5158_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ),
    .A2(net141),
    .B1(net83),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ),
    .C1(net79),
    .X(_2099_));
 sky130_fd_sc_hd__o221a_1 _5159_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ),
    .A2(net141),
    .B1(net83),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][3] ),
    .C1(net80),
    .X(_2100_));
 sky130_fd_sc_hd__or2_1 _5160_ (.A(_2099_),
    .B(_2100_),
    .X(_2101_));
 sky130_fd_sc_hd__mux4_2 _5161_ (.A0(_0971_),
    .A1(_1308_),
    .A2(_2098_),
    .A3(_2101_),
    .S0(_2045_),
    .S1(_0808_),
    .X(_2102_));
 sky130_fd_sc_hd__a22o_1 _5162_ (.A1(\z80.tv80s.i_tv80_core.ACC[3] ),
    .A2(_2052_),
    .B1(_2053_),
    .B2(_2102_),
    .X(_2103_));
 sky130_fd_sc_hd__or4_1 _5163_ (.A(_2093_),
    .B(_2094_),
    .C(_2095_),
    .D(_2103_),
    .X(_2104_));
 sky130_fd_sc_hd__a22o_1 _5164_ (.A1(net160),
    .A2(net627),
    .B1(_2030_),
    .B2(_2104_),
    .X(_0234_));
 sky130_fd_sc_hd__a22o_1 _5165_ (.A1(\z80.tv80s.i_tv80_core.SP[4] ),
    .A2(_2050_),
    .B1(_2052_),
    .B2(\z80.tv80s.i_tv80_core.ACC[4] ),
    .X(_2105_));
 sky130_fd_sc_hd__a22o_1 _5166_ (.A1(\z80.tv80s.di_reg[4] ),
    .A2(_2065_),
    .B1(_2066_),
    .B2(\z80.tv80s.i_tv80_core.PC[4] ),
    .X(_2106_));
 sky130_fd_sc_hd__o221a_1 _5167_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ),
    .A2(net141),
    .B1(net83),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ),
    .C1(_0733_),
    .X(_2107_));
 sky130_fd_sc_hd__o221a_1 _5168_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ),
    .A2(net140),
    .B1(net85),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ),
    .C1(net81),
    .X(_2108_));
 sky130_fd_sc_hd__or2_1 _5169_ (.A(_2107_),
    .B(_2108_),
    .X(_2109_));
 sky130_fd_sc_hd__o221a_1 _5170_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ),
    .A2(net141),
    .B1(net84),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][4] ),
    .C1(net79),
    .X(_2110_));
 sky130_fd_sc_hd__o221a_1 _5171_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ),
    .A2(net141),
    .B1(net84),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][4] ),
    .C1(net80),
    .X(_2111_));
 sky130_fd_sc_hd__or2_1 _5172_ (.A(_2110_),
    .B(_2111_),
    .X(_2112_));
 sky130_fd_sc_hd__mux4_2 _5173_ (.A0(_1014_),
    .A1(_1325_),
    .A2(_2109_),
    .A3(_2112_),
    .S0(_2045_),
    .S1(_0808_),
    .X(_2113_));
 sky130_fd_sc_hd__a22o_1 _5174_ (.A1(\z80.tv80s.i_tv80_core.PC[12] ),
    .A2(_2063_),
    .B1(_2113_),
    .B2(_2053_),
    .X(_2114_));
 sky130_fd_sc_hd__a221o_1 _5175_ (.A1(\z80.tv80s.i_tv80_core.F[4] ),
    .A2(_2048_),
    .B1(_2072_),
    .B2(\z80.tv80s.i_tv80_core.SP[12] ),
    .C1(_2114_),
    .X(_2115_));
 sky130_fd_sc_hd__or3_1 _5176_ (.A(_2105_),
    .B(_2106_),
    .C(_2115_),
    .X(_2116_));
 sky130_fd_sc_hd__a22o_1 _5177_ (.A1(net157),
    .A2(net590),
    .B1(_2030_),
    .B2(_2116_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_1 _5178_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ),
    .S(net81),
    .X(_2117_));
 sky130_fd_sc_hd__mux2_1 _5179_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][5] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ),
    .S(net81),
    .X(_2118_));
 sky130_fd_sc_hd__o22a_1 _5180_ (.A1(net85),
    .A2(_2117_),
    .B1(_2118_),
    .B2(net140),
    .X(_2119_));
 sky130_fd_sc_hd__mux2_1 _5181_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ),
    .S(net80),
    .X(_2120_));
 sky130_fd_sc_hd__mux2_1 _5182_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ),
    .S(net80),
    .X(_2121_));
 sky130_fd_sc_hd__o22a_1 _5183_ (.A1(net84),
    .A2(_2120_),
    .B1(_2121_),
    .B2(net141),
    .X(_2122_));
 sky130_fd_sc_hd__mux2_1 _5184_ (.A0(_2119_),
    .A1(_2122_),
    .S(_2045_),
    .X(_2123_));
 sky130_fd_sc_hd__mux2_1 _5185_ (.A0(_1063_),
    .A1(_1339_),
    .S(_2045_),
    .X(_2124_));
 sky130_fd_sc_hd__mux2_1 _5186_ (.A0(_2123_),
    .A1(_2124_),
    .S(_0809_),
    .X(_2125_));
 sky130_fd_sc_hd__a22o_1 _5187_ (.A1(\z80.tv80s.i_tv80_core.F[5] ),
    .A2(_2048_),
    .B1(_2050_),
    .B2(\z80.tv80s.i_tv80_core.SP[5] ),
    .X(_2126_));
 sky130_fd_sc_hd__a22o_1 _5188_ (.A1(\z80.tv80s.i_tv80_core.ACC[5] ),
    .A2(_2052_),
    .B1(_2063_),
    .B2(\z80.tv80s.i_tv80_core.PC[13] ),
    .X(_2127_));
 sky130_fd_sc_hd__a22o_1 _5189_ (.A1(\z80.tv80s.i_tv80_core.PC[5] ),
    .A2(_2066_),
    .B1(_2125_),
    .B2(_2053_),
    .X(_2128_));
 sky130_fd_sc_hd__a211o_1 _5190_ (.A1(\z80.tv80s.di_reg[5] ),
    .A2(_2065_),
    .B1(_2126_),
    .C1(_2128_),
    .X(_2129_));
 sky130_fd_sc_hd__a211o_1 _5191_ (.A1(\z80.tv80s.i_tv80_core.SP[13] ),
    .A2(_2072_),
    .B1(_2127_),
    .C1(_2129_),
    .X(_2130_));
 sky130_fd_sc_hd__a22o_1 _5192_ (.A1(net157),
    .A2(net605),
    .B1(_2030_),
    .B2(_2130_),
    .X(_0236_));
 sky130_fd_sc_hd__a22o_1 _5193_ (.A1(\z80.tv80s.i_tv80_core.F[6] ),
    .A2(_2048_),
    .B1(_2050_),
    .B2(\z80.tv80s.i_tv80_core.SP[6] ),
    .X(_2131_));
 sky130_fd_sc_hd__a22o_1 _5194_ (.A1(\z80.tv80s.i_tv80_core.ACC[6] ),
    .A2(_2052_),
    .B1(_2072_),
    .B2(net473),
    .X(_2132_));
 sky130_fd_sc_hd__a22o_1 _5195_ (.A1(\z80.tv80s.i_tv80_core.PC[14] ),
    .A2(_2063_),
    .B1(_2065_),
    .B2(\z80.tv80s.di_reg[6] ),
    .X(_2133_));
 sky130_fd_sc_hd__o221a_1 _5196_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ),
    .A2(net140),
    .B1(net82),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ),
    .C1(net79),
    .X(_2134_));
 sky130_fd_sc_hd__o221a_1 _5197_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][6] ),
    .A2(net140),
    .B1(net82),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ),
    .C1(net81),
    .X(_2135_));
 sky130_fd_sc_hd__or2_1 _5198_ (.A(_2134_),
    .B(_2135_),
    .X(_2136_));
 sky130_fd_sc_hd__o221a_1 _5199_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ),
    .A2(net141),
    .B1(net83),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ),
    .C1(net79),
    .X(_2137_));
 sky130_fd_sc_hd__o221a_1 _5200_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ),
    .A2(net141),
    .B1(net83),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ),
    .C1(net80),
    .X(_2138_));
 sky130_fd_sc_hd__or2_1 _5201_ (.A(_2137_),
    .B(_2138_),
    .X(_2139_));
 sky130_fd_sc_hd__mux4_2 _5202_ (.A0(_1111_),
    .A1(_1354_),
    .A2(_2136_),
    .A3(_2139_),
    .S0(_2045_),
    .S1(_0808_),
    .X(_2140_));
 sky130_fd_sc_hd__a22o_1 _5203_ (.A1(\z80.tv80s.i_tv80_core.PC[6] ),
    .A2(_2066_),
    .B1(_2140_),
    .B2(_2053_),
    .X(_2141_));
 sky130_fd_sc_hd__or4_1 _5204_ (.A(_2131_),
    .B(_2132_),
    .C(_2133_),
    .D(_2141_),
    .X(_2142_));
 sky130_fd_sc_hd__a22o_1 _5205_ (.A1(net156),
    .A2(net601),
    .B1(_2030_),
    .B2(_2142_),
    .X(_0237_));
 sky130_fd_sc_hd__a22o_1 _5206_ (.A1(\z80.tv80s.i_tv80_core.F[7] ),
    .A2(_2048_),
    .B1(_2066_),
    .B2(\z80.tv80s.i_tv80_core.PC[7] ),
    .X(_2143_));
 sky130_fd_sc_hd__o221a_1 _5207_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ),
    .A2(net140),
    .B1(net82),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][7] ),
    .C1(net79),
    .X(_2144_));
 sky130_fd_sc_hd__o221a_1 _5208_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][7] ),
    .A2(net140),
    .B1(net85),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][7] ),
    .C1(net81),
    .X(_2145_));
 sky130_fd_sc_hd__or3_1 _5209_ (.A(_0809_),
    .B(_2144_),
    .C(_2145_),
    .X(_2146_));
 sky130_fd_sc_hd__o211a_1 _5210_ (.A1(_0808_),
    .A2(_1165_),
    .B1(_2046_),
    .C1(_2146_),
    .X(_2147_));
 sky130_fd_sc_hd__a21o_1 _5211_ (.A1(_1372_),
    .A2(_2045_),
    .B1(_2147_),
    .X(_2148_));
 sky130_fd_sc_hd__a221o_1 _5212_ (.A1(\z80.tv80s.di_reg[7] ),
    .A2(_2065_),
    .B1(_2072_),
    .B2(\z80.tv80s.i_tv80_core.SP[15] ),
    .C1(_2143_),
    .X(_2149_));
 sky130_fd_sc_hd__a221o_1 _5213_ (.A1(\z80.tv80s.i_tv80_core.PC[15] ),
    .A2(_2063_),
    .B1(_2148_),
    .B2(_2053_),
    .C1(_2149_),
    .X(_2150_));
 sky130_fd_sc_hd__a221o_1 _5214_ (.A1(\z80.tv80s.i_tv80_core.SP[7] ),
    .A2(_2050_),
    .B1(_2052_),
    .B2(\z80.tv80s.i_tv80_core.ACC[7] ),
    .C1(_2150_),
    .X(_2151_));
 sky130_fd_sc_hd__a22o_1 _5215_ (.A1(net157),
    .A2(net625),
    .B1(_2030_),
    .B2(_2151_),
    .X(_0238_));
 sky130_fd_sc_hd__and2_2 _5216_ (.A(_0446_),
    .B(_0522_),
    .X(_2152_));
 sky130_fd_sc_hd__inv_2 _5217_ (.A(_2152_),
    .Y(_2153_));
 sky130_fd_sc_hd__and2_2 _5218_ (.A(_2697_),
    .B(_0648_),
    .X(_2154_));
 sky130_fd_sc_hd__nor2_1 _5219_ (.A(_0033_),
    .B(_0034_),
    .Y(_2155_));
 sky130_fd_sc_hd__nor2_1 _5220_ (.A(_2697_),
    .B(net713),
    .Y(_2156_));
 sky130_fd_sc_hd__or3_1 _5221_ (.A(net733),
    .B(net802),
    .C(net713),
    .X(_2157_));
 sky130_fd_sc_hd__nand3_1 _5222_ (.A(net733),
    .B(net802),
    .C(net713),
    .Y(_2158_));
 sky130_fd_sc_hd__a31o_1 _5223_ (.A1(net142),
    .A2(_2157_),
    .A3(_2158_),
    .B1(_2154_),
    .X(_2159_));
 sky130_fd_sc_hd__a2bb2o_1 _5224_ (.A1_N(_2153_),
    .A2_N(_2159_),
    .B1(net147),
    .B2(_0521_),
    .X(_0239_));
 sky130_fd_sc_hd__and2b_1 _5225_ (.A_N(_0034_),
    .B(net733),
    .X(_2160_));
 sky130_fd_sc_hd__a22o_1 _5226_ (.A1(net147),
    .A2(_2154_),
    .B1(_2156_),
    .B2(net734),
    .X(_2161_));
 sky130_fd_sc_hd__a22o_1 _5227_ (.A1(net145),
    .A2(_0521_),
    .B1(_2152_),
    .B2(_2161_),
    .X(_0240_));
 sky130_fd_sc_hd__and2b_1 _5228_ (.A_N(net733),
    .B(net802),
    .X(_2162_));
 sky130_fd_sc_hd__a22o_1 _5229_ (.A1(net145),
    .A2(_2154_),
    .B1(_2156_),
    .B2(_2162_),
    .X(_2163_));
 sky130_fd_sc_hd__a22o_1 _5230_ (.A1(net143),
    .A2(_0521_),
    .B1(_2152_),
    .B2(_2163_),
    .X(_0241_));
 sky130_fd_sc_hd__a32o_1 _5231_ (.A1(net733),
    .A2(net802),
    .A3(_2156_),
    .B1(_2154_),
    .B2(net143),
    .X(_2164_));
 sky130_fd_sc_hd__a22o_1 _5232_ (.A1(net821),
    .A2(_0521_),
    .B1(_2152_),
    .B2(_2164_),
    .X(_0242_));
 sky130_fd_sc_hd__a32o_1 _5233_ (.A1(net142),
    .A2(net713),
    .A3(_2155_),
    .B1(_2154_),
    .B2(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .X(_2165_));
 sky130_fd_sc_hd__a22o_1 _5234_ (.A1(net267),
    .A2(_0521_),
    .B1(_2152_),
    .B2(net714),
    .X(_0243_));
 sky130_fd_sc_hd__a32o_1 _5235_ (.A1(net142),
    .A2(net713),
    .A3(net734),
    .B1(_2154_),
    .B2(net267),
    .X(_2166_));
 sky130_fd_sc_hd__o22a_1 _5236_ (.A1(net555),
    .A2(_0522_),
    .B1(_2153_),
    .B2(net735),
    .X(_0244_));
 sky130_fd_sc_hd__a32o_1 _5237_ (.A1(net142),
    .A2(net713),
    .A3(_2162_),
    .B1(_2154_),
    .B2(net555),
    .X(_2167_));
 sky130_fd_sc_hd__a22o_1 _5238_ (.A1(net142),
    .A2(_0521_),
    .B1(_2152_),
    .B2(net803),
    .X(_0245_));
 sky130_fd_sc_hd__a21o_1 _5239_ (.A1(_0445_),
    .A2(_1233_),
    .B1(_1221_),
    .X(_2168_));
 sky130_fd_sc_hd__mux2_1 _5240_ (.A0(net140),
    .A1(_2168_),
    .S(net109),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _5241_ (.A0(net524),
    .A1(_1233_),
    .S(net110),
    .X(_0247_));
 sky130_fd_sc_hd__and2b_1 _5242_ (.A_N(net10),
    .B(\z80.tv80s.i_tv80_core.Oldnmi_n ),
    .X(_2169_));
 sky130_fd_sc_hd__o21ba_1 _5243_ (.A1(net504),
    .A2(_2169_),
    .B1_N(net519),
    .X(_0248_));
 sky130_fd_sc_hd__o21a_1 _5244_ (.A1(_1191_),
    .A2(_1204_),
    .B1(_1418_),
    .X(_2170_));
 sky130_fd_sc_hd__nor2_2 _5245_ (.A(net159),
    .B(_2170_),
    .Y(_2171_));
 sky130_fd_sc_hd__nand2_1 _5246_ (.A(_1261_),
    .B(_1406_),
    .Y(_2172_));
 sky130_fd_sc_hd__nand2_1 _5247_ (.A(_1191_),
    .B(_1204_),
    .Y(_2173_));
 sky130_fd_sc_hd__a21oi_4 _5248_ (.A1(_1191_),
    .A2(_1204_),
    .B1(_1418_),
    .Y(_2174_));
 sky130_fd_sc_hd__nand2_1 _5249_ (.A(_0760_),
    .B(_1407_),
    .Y(_2175_));
 sky130_fd_sc_hd__or3b_1 _5250_ (.A(_1191_),
    .B(_1204_),
    .C_N(_1418_),
    .X(_2176_));
 sky130_fd_sc_hd__nor2_2 _5251_ (.A(_1407_),
    .B(_2176_),
    .Y(_2177_));
 sky130_fd_sc_hd__nor2_2 _5252_ (.A(_1406_),
    .B(_2176_),
    .Y(_2178_));
 sky130_fd_sc_hd__nor2_2 _5253_ (.A(_1407_),
    .B(_2173_),
    .Y(_2179_));
 sky130_fd_sc_hd__nor2_2 _5254_ (.A(_1406_),
    .B(_2173_),
    .Y(_2180_));
 sky130_fd_sc_hd__a22o_1 _5255_ (.A1(\z80.tv80s.di_reg[0] ),
    .A2(_2179_),
    .B1(_2180_),
    .B2(\z80.tv80s.i_tv80_core.ACC[0] ),
    .X(_2181_));
 sky130_fd_sc_hd__a221o_1 _5256_ (.A1(\z80.tv80s.i_tv80_core.SP[0] ),
    .A2(_2177_),
    .B1(_2178_),
    .B2(net703),
    .C1(_2181_),
    .X(_2182_));
 sky130_fd_sc_hd__a31o_1 _5257_ (.A1(_2172_),
    .A2(_2174_),
    .A3(_2175_),
    .B1(_2182_),
    .X(_2183_));
 sky130_fd_sc_hd__a22o_1 _5258_ (.A1(net159),
    .A2(net725),
    .B1(_2171_),
    .B2(_2183_),
    .X(_0249_));
 sky130_fd_sc_hd__nand2_1 _5259_ (.A(_0866_),
    .B(_1407_),
    .Y(_2184_));
 sky130_fd_sc_hd__o211a_1 _5260_ (.A1(_1275_),
    .A2(_1407_),
    .B1(_2174_),
    .C1(_2184_),
    .X(_2185_));
 sky130_fd_sc_hd__a221o_1 _5261_ (.A1(\z80.tv80s.di_reg[1] ),
    .A2(_2179_),
    .B1(_2180_),
    .B2(\z80.tv80s.i_tv80_core.ACC[1] ),
    .C1(_2185_),
    .X(_2186_));
 sky130_fd_sc_hd__a221o_1 _5262_ (.A1(net723),
    .A2(_2177_),
    .B1(_2178_),
    .B2(\z80.tv80s.i_tv80_core.SP[9] ),
    .C1(_2186_),
    .X(_2187_));
 sky130_fd_sc_hd__a22o_1 _5263_ (.A1(net158),
    .A2(net739),
    .B1(_2171_),
    .B2(_2187_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _5264_ (.A0(_0892_),
    .A1(_1288_),
    .S(_1406_),
    .X(_2188_));
 sky130_fd_sc_hd__a22o_1 _5265_ (.A1(\z80.tv80s.di_reg[2] ),
    .A2(_2179_),
    .B1(_2180_),
    .B2(\z80.tv80s.i_tv80_core.ACC[2] ),
    .X(_2189_));
 sky130_fd_sc_hd__a221o_1 _5266_ (.A1(\z80.tv80s.i_tv80_core.SP[2] ),
    .A2(_2177_),
    .B1(_2178_),
    .B2(\z80.tv80s.i_tv80_core.SP[10] ),
    .C1(_2189_),
    .X(_2190_));
 sky130_fd_sc_hd__a21o_1 _5267_ (.A1(_2174_),
    .A2(_2188_),
    .B1(_2190_),
    .X(_2191_));
 sky130_fd_sc_hd__a22o_1 _5268_ (.A1(net158),
    .A2(net636),
    .B1(_2171_),
    .B2(_2191_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _5269_ (.A0(_0933_),
    .A1(_1302_),
    .S(_1406_),
    .X(_2192_));
 sky130_fd_sc_hd__a22o_1 _5270_ (.A1(\z80.tv80s.di_reg[3] ),
    .A2(_2179_),
    .B1(_2180_),
    .B2(\z80.tv80s.i_tv80_core.ACC[3] ),
    .X(_2193_));
 sky130_fd_sc_hd__a221o_1 _5271_ (.A1(\z80.tv80s.i_tv80_core.SP[3] ),
    .A2(_2177_),
    .B1(_2178_),
    .B2(\z80.tv80s.i_tv80_core.SP[11] ),
    .C1(_2193_),
    .X(_2194_));
 sky130_fd_sc_hd__a21o_1 _5272_ (.A1(_2174_),
    .A2(_2192_),
    .B1(_2194_),
    .X(_2195_));
 sky130_fd_sc_hd__a22o_1 _5273_ (.A1(net158),
    .A2(net617),
    .B1(_2171_),
    .B2(_2195_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _5274_ (.A0(_1008_),
    .A1(_1318_),
    .S(_1406_),
    .X(_2196_));
 sky130_fd_sc_hd__a22o_1 _5275_ (.A1(\z80.tv80s.di_reg[4] ),
    .A2(_2179_),
    .B1(_2180_),
    .B2(\z80.tv80s.i_tv80_core.ACC[4] ),
    .X(_2197_));
 sky130_fd_sc_hd__a221o_1 _5276_ (.A1(\z80.tv80s.i_tv80_core.SP[4] ),
    .A2(_2177_),
    .B1(_2178_),
    .B2(\z80.tv80s.i_tv80_core.SP[12] ),
    .C1(_2197_),
    .X(_2198_));
 sky130_fd_sc_hd__a21o_1 _5277_ (.A1(_2174_),
    .A2(_2196_),
    .B1(_2198_),
    .X(_2199_));
 sky130_fd_sc_hd__a22o_1 _5278_ (.A1(net159),
    .A2(net633),
    .B1(_2171_),
    .B2(_2199_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _5279_ (.A0(_1022_),
    .A1(_1331_),
    .S(_1406_),
    .X(_2200_));
 sky130_fd_sc_hd__a22o_1 _5280_ (.A1(\z80.tv80s.di_reg[5] ),
    .A2(_2179_),
    .B1(_2180_),
    .B2(\z80.tv80s.i_tv80_core.ACC[5] ),
    .X(_2201_));
 sky130_fd_sc_hd__a221o_1 _5281_ (.A1(\z80.tv80s.i_tv80_core.SP[5] ),
    .A2(_2177_),
    .B1(_2178_),
    .B2(\z80.tv80s.i_tv80_core.SP[13] ),
    .C1(_2201_),
    .X(_2202_));
 sky130_fd_sc_hd__a21o_1 _5282_ (.A1(_2174_),
    .A2(_2200_),
    .B1(_2202_),
    .X(_2203_));
 sky130_fd_sc_hd__a22o_1 _5283_ (.A1(net158),
    .A2(net623),
    .B1(_2171_),
    .B2(_2203_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _5284_ (.A0(_1102_),
    .A1(_1346_),
    .S(_1406_),
    .X(_2204_));
 sky130_fd_sc_hd__a22o_1 _5285_ (.A1(\z80.tv80s.di_reg[6] ),
    .A2(_2179_),
    .B1(_2180_),
    .B2(\z80.tv80s.i_tv80_core.ACC[6] ),
    .X(_2205_));
 sky130_fd_sc_hd__a221o_1 _5286_ (.A1(\z80.tv80s.i_tv80_core.SP[6] ),
    .A2(_2177_),
    .B1(_2178_),
    .B2(net473),
    .C1(_2205_),
    .X(_2206_));
 sky130_fd_sc_hd__a21o_1 _5287_ (.A1(_2174_),
    .A2(_2204_),
    .B1(_2206_),
    .X(_2207_));
 sky130_fd_sc_hd__a22o_1 _5288_ (.A1(net159),
    .A2(net699),
    .B1(_2171_),
    .B2(_2207_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _5289_ (.A0(_1121_),
    .A1(_1361_),
    .S(_1406_),
    .X(_2208_));
 sky130_fd_sc_hd__a22o_1 _5290_ (.A1(net853),
    .A2(_2179_),
    .B1(_2180_),
    .B2(net808),
    .X(_2209_));
 sky130_fd_sc_hd__a221o_1 _5291_ (.A1(net800),
    .A2(_2177_),
    .B1(_2178_),
    .B2(net771),
    .C1(_2209_),
    .X(_2210_));
 sky130_fd_sc_hd__a21o_1 _5292_ (.A1(_2174_),
    .A2(_2208_),
    .B1(_2210_),
    .X(_2211_));
 sky130_fd_sc_hd__a22o_1 _5293_ (.A1(net159),
    .A2(net139),
    .B1(_2171_),
    .B2(_2211_),
    .X(_0256_));
 sky130_fd_sc_hd__a21o_1 _5294_ (.A1(_0445_),
    .A2(_1204_),
    .B1(_1191_),
    .X(_2212_));
 sky130_fd_sc_hd__mux2_1 _5295_ (.A0(net265),
    .A1(_2212_),
    .S(net110),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _5296_ (.A0(net240),
    .A1(_1204_),
    .S(net109),
    .X(_0258_));
 sky130_fd_sc_hd__nor2_4 _5297_ (.A(_0709_),
    .B(_0751_),
    .Y(_2213_));
 sky130_fd_sc_hd__mux2_1 _5298_ (.A0(net301),
    .A1(_0807_),
    .S(_2213_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _5299_ (.A0(net349),
    .A1(_0875_),
    .S(_2213_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _5300_ (.A0(net291),
    .A1(_0926_),
    .S(_2213_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _5301_ (.A0(net329),
    .A1(_0972_),
    .S(_2213_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _5302_ (.A0(net277),
    .A1(_1015_),
    .S(_2213_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _5303_ (.A0(net433),
    .A1(_1064_),
    .S(_2213_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _5304_ (.A0(net396),
    .A1(_1112_),
    .S(_2213_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _5305_ (.A0(net293),
    .A1(_1166_),
    .S(_2213_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _5306_ (.A0(net1),
    .A1(net854),
    .S(_0546_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _5307_ (.A0(net2),
    .A1(net849),
    .S(_0546_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _5308_ (.A0(net3),
    .A1(net848),
    .S(_0546_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _5309_ (.A0(net4),
    .A1(net840),
    .S(_0546_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _5310_ (.A0(net5),
    .A1(net846),
    .S(_0546_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _5311_ (.A0(net6),
    .A1(net852),
    .S(_0546_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _5312_ (.A0(net7),
    .A1(net847),
    .S(_0546_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _5313_ (.A0(net8),
    .A1(net853),
    .S(_0546_),
    .X(_0274_));
 sky130_fd_sc_hd__nor2_1 _5314_ (.A(net749),
    .B(net54),
    .Y(_2214_));
 sky130_fd_sc_hd__o221a_1 _5315_ (.A1(net515),
    .A2(_0500_),
    .B1(_0637_),
    .B2(net450),
    .C1(net54),
    .X(_2215_));
 sky130_fd_sc_hd__o21ai_4 _5316_ (.A1(_2214_),
    .A2(_2215_),
    .B1(_0663_),
    .Y(_2216_));
 sky130_fd_sc_hd__nor2_2 _5317_ (.A(_0518_),
    .B(_2216_),
    .Y(_2217_));
 sky130_fd_sc_hd__a22o_1 _5318_ (.A1(\z80.tv80s.i_tv80_core.ts[0] ),
    .A2(_2216_),
    .B1(_2217_),
    .B2(net497),
    .X(_0275_));
 sky130_fd_sc_hd__or2_1 _5319_ (.A(net716),
    .B(_0516_),
    .X(_2218_));
 sky130_fd_sc_hd__mux2_1 _5320_ (.A0(_2218_),
    .A1(net656),
    .S(_2216_),
    .X(_0276_));
 sky130_fd_sc_hd__a22o_1 _5321_ (.A1(\z80.tv80s.i_tv80_core.ts[2] ),
    .A2(_2216_),
    .B1(_2217_),
    .B2(net656),
    .X(_0277_));
 sky130_fd_sc_hd__a22o_1 _5322_ (.A1(net136),
    .A2(_2216_),
    .B1(_2217_),
    .B2(net844),
    .X(_0278_));
 sky130_fd_sc_hd__a22o_1 _5323_ (.A1(net398),
    .A2(_2216_),
    .B1(_2217_),
    .B2(net136),
    .X(_0279_));
 sky130_fd_sc_hd__a22o_1 _5324_ (.A1(net255),
    .A2(_2216_),
    .B1(_2217_),
    .B2(net398),
    .X(_0280_));
 sky130_fd_sc_hd__a22o_1 _5325_ (.A1(net874),
    .A2(_2216_),
    .B1(_2217_),
    .B2(net255),
    .X(_0281_));
 sky130_fd_sc_hd__and4b_2 _5326_ (.A_N(net542),
    .B(net635),
    .C(_0673_),
    .D(net679),
    .X(_2219_));
 sky130_fd_sc_hd__nand4b_4 _5327_ (.A_N(net542),
    .B(net635),
    .C(_0673_),
    .D(net679),
    .Y(_2220_));
 sky130_fd_sc_hd__a21oi_4 _5328_ (.A1(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .A2(_0642_),
    .B1(_0785_),
    .Y(_2221_));
 sky130_fd_sc_hd__a21o_2 _5329_ (.A1(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .A2(_0642_),
    .B1(_0785_),
    .X(_2222_));
 sky130_fd_sc_hd__or2_1 _5330_ (.A(net543),
    .B(_2221_),
    .X(_2223_));
 sky130_fd_sc_hd__a21bo_1 _5331_ (.A1(\z80.tv80s.i_tv80_core.BusA[7] ),
    .A2(_1126_),
    .B1_N(_1130_),
    .X(_2224_));
 sky130_fd_sc_hd__nor2_1 _5332_ (.A(_1986_),
    .B(_2224_),
    .Y(_2225_));
 sky130_fd_sc_hd__nor2_1 _5333_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(net154),
    .Y(_2226_));
 sky130_fd_sc_hd__a21o_1 _5334_ (.A1(_2224_),
    .A2(_2226_),
    .B1(_2225_),
    .X(_2227_));
 sky130_fd_sc_hd__a21o_1 _5335_ (.A1(net119),
    .A2(net139),
    .B1(_1154_),
    .X(_2228_));
 sky130_fd_sc_hd__a32o_1 _5336_ (.A1(\z80.tv80s.i_tv80_core.F[0] ),
    .A2(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .A3(_0771_),
    .B1(_0791_),
    .B2(_2228_),
    .X(_2229_));
 sky130_fd_sc_hd__a221o_1 _5337_ (.A1(_0789_),
    .A2(_1043_),
    .B1(_2227_),
    .B2(_2722_),
    .C1(_2229_),
    .X(_2230_));
 sky130_fd_sc_hd__nor4_1 _5338_ (.A(_0629_),
    .B(_1431_),
    .C(_1435_),
    .D(_1483_),
    .Y(_2231_));
 sky130_fd_sc_hd__and2_4 _5339_ (.A(net168),
    .B(net93),
    .X(_2232_));
 sky130_fd_sc_hd__nand2_1 _5340_ (.A(net168),
    .B(net93),
    .Y(_2233_));
 sky130_fd_sc_hd__nand2_4 _5341_ (.A(net101),
    .B(_2232_),
    .Y(_2234_));
 sky130_fd_sc_hd__nand2_1 _5342_ (.A(_1387_),
    .B(_2234_),
    .Y(_2235_));
 sky130_fd_sc_hd__o311a_2 _5343_ (.A1(_2779_),
    .A2(_2790_),
    .A3(_2811_),
    .B1(_1736_),
    .C1(_2231_),
    .X(_2236_));
 sky130_fd_sc_hd__a32o_1 _5344_ (.A1(net168),
    .A2(_2789_),
    .A3(_2812_),
    .B1(_2236_),
    .B2(_2710_),
    .X(_2237_));
 sky130_fd_sc_hd__o21ai_1 _5345_ (.A1(_2710_),
    .A2(_2236_),
    .B1(_2233_),
    .Y(_2238_));
 sky130_fd_sc_hd__o32a_1 _5346_ (.A1(net55),
    .A2(_2237_),
    .A3(_2238_),
    .B1(_2233_),
    .B2(net673),
    .X(_2239_));
 sky130_fd_sc_hd__o22a_1 _5347_ (.A1(\z80.tv80s.i_tv80_core.F[0] ),
    .A2(_2235_),
    .B1(_2239_),
    .B2(_0540_),
    .X(_2240_));
 sky130_fd_sc_hd__mux2_1 _5348_ (.A0(_2230_),
    .A1(_2240_),
    .S(_2223_),
    .X(_2241_));
 sky130_fd_sc_hd__mux2_1 _5349_ (.A0(_0803_),
    .A1(_2241_),
    .S(_2220_),
    .X(_2242_));
 sky130_fd_sc_hd__mux2_1 _5350_ (.A0(net866),
    .A1(_2242_),
    .S(net112),
    .X(_0282_));
 sky130_fd_sc_hd__or4bb_4 _5351_ (.A(net115),
    .B(net54),
    .C_N(_2231_),
    .D_N(_0411_),
    .X(_2243_));
 sky130_fd_sc_hd__inv_2 _5352_ (.A(_2243_),
    .Y(_2244_));
 sky130_fd_sc_hd__a31oi_2 _5353_ (.A1(net168),
    .A2(_2789_),
    .A3(_2812_),
    .B1(_2236_),
    .Y(_2245_));
 sky130_fd_sc_hd__nor2_1 _5354_ (.A(net55),
    .B(_2245_),
    .Y(_2246_));
 sky130_fd_sc_hd__o2bb2a_1 _5355_ (.A1_N(net101),
    .A2_N(_2246_),
    .B1(_2244_),
    .B2(\z80.tv80s.i_tv80_core.F[1] ),
    .X(_2247_));
 sky130_fd_sc_hd__and4_4 _5356_ (.A(net123),
    .B(\z80.tv80s.i_tv80_core.ts[3] ),
    .C(_2854_),
    .D(_0377_),
    .X(_2248_));
 sky130_fd_sc_hd__clkinv_4 _5357_ (.A(_2248_),
    .Y(_2249_));
 sky130_fd_sc_hd__o22a_1 _5358_ (.A1(net695),
    .A2(_2234_),
    .B1(_2247_),
    .B2(_2232_),
    .X(_2250_));
 sky130_fd_sc_hd__o211a_1 _5359_ (.A1(\z80.tv80s.i_tv80_core.F[1] ),
    .A2(net101),
    .B1(_2249_),
    .C1(_2250_),
    .X(_2251_));
 sky130_fd_sc_hd__or4_4 _5360_ (.A(_2705_),
    .B(net106),
    .C(net54),
    .D(_1182_),
    .X(_2252_));
 sky130_fd_sc_hd__inv_2 _5361_ (.A(_2252_),
    .Y(_2253_));
 sky130_fd_sc_hd__or4_4 _5362_ (.A(_2713_),
    .B(_2838_),
    .C(net106),
    .D(_0587_),
    .X(_2254_));
 sky130_fd_sc_hd__and3_1 _5363_ (.A(_2220_),
    .B(_2252_),
    .C(_2254_),
    .X(_2255_));
 sky130_fd_sc_hd__o2bb2a_1 _5364_ (.A1_N(_0790_),
    .A2_N(_1986_),
    .B1(_2722_),
    .B2(\z80.tv80s.i_tv80_core.F[1] ),
    .X(_2256_));
 sky130_fd_sc_hd__mux2_1 _5365_ (.A0(_2251_),
    .A1(_2256_),
    .S(_2222_),
    .X(_2257_));
 sky130_fd_sc_hd__a22o_1 _5366_ (.A1(_0845_),
    .A2(_2219_),
    .B1(_2255_),
    .B2(_2257_),
    .X(_2258_));
 sky130_fd_sc_hd__mux2_1 _5367_ (.A0(net868),
    .A1(_2258_),
    .S(net112),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _5368_ (.A0(\z80.tv80s.i_tv80_core.Fp[2] ),
    .A1(\z80.tv80s.i_tv80_core.F[2] ),
    .S(_2234_),
    .X(_2259_));
 sky130_fd_sc_hd__mux2_1 _5369_ (.A0(_2259_),
    .A1(\z80.tv80s.i_tv80_core.IntE_FF2 ),
    .S(_2248_),
    .X(_2260_));
 sky130_fd_sc_hd__or3b_1 _5370_ (.A(\z80.tv80s.i_tv80_core.BusA[7] ),
    .B(_1128_),
    .C_N(_1126_),
    .X(_2261_));
 sky130_fd_sc_hd__o21ai_1 _5371_ (.A1(_1126_),
    .A2(_1130_),
    .B1(_2261_),
    .Y(_2262_));
 sky130_fd_sc_hd__xnor2_1 _5372_ (.A(_1074_),
    .B(_1136_),
    .Y(_2263_));
 sky130_fd_sc_hd__xnor2_1 _5373_ (.A(_0995_),
    .B(_1038_),
    .Y(_2264_));
 sky130_fd_sc_hd__xor2_1 _5374_ (.A(_0781_),
    .B(_0828_),
    .X(_2265_));
 sky130_fd_sc_hd__xnor2_1 _5375_ (.A(_0907_),
    .B(_0951_),
    .Y(_2266_));
 sky130_fd_sc_hd__xnor2_1 _5376_ (.A(_2265_),
    .B(_2266_),
    .Y(_2267_));
 sky130_fd_sc_hd__xnor2_1 _5377_ (.A(_2264_),
    .B(_2267_),
    .Y(_2268_));
 sky130_fd_sc_hd__nor2_1 _5378_ (.A(_2263_),
    .B(_2268_),
    .Y(_2269_));
 sky130_fd_sc_hd__a21o_1 _5379_ (.A1(_2263_),
    .A2(_2268_),
    .B1(_0777_),
    .X(_2270_));
 sky130_fd_sc_hd__o22a_1 _5380_ (.A1(_0776_),
    .A2(_2262_),
    .B1(_2269_),
    .B2(_2270_),
    .X(_2271_));
 sky130_fd_sc_hd__a21oi_1 _5381_ (.A1(_2709_),
    .A2(\z80.tv80s.i_tv80_core.Arith16_r ),
    .B1(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .Y(_2272_));
 sky130_fd_sc_hd__o21a_1 _5382_ (.A1(\z80.tv80s.i_tv80_core.Arith16_r ),
    .A2(_2271_),
    .B1(_2272_),
    .X(_2273_));
 sky130_fd_sc_hd__xnor2_1 _5383_ (.A(\z80.tv80s.i_tv80_core.BusA[0] ),
    .B(_0840_),
    .Y(_2274_));
 sky130_fd_sc_hd__xor2_1 _5384_ (.A(_1082_),
    .B(_1148_),
    .X(_2275_));
 sky130_fd_sc_hd__xnor2_1 _5385_ (.A(_2274_),
    .B(_2275_),
    .Y(_2276_));
 sky130_fd_sc_hd__xnor2_1 _5386_ (.A(_0975_),
    .B(_1050_),
    .Y(_2277_));
 sky130_fd_sc_hd__xnor2_1 _5387_ (.A(_0910_),
    .B(_0957_),
    .Y(_2278_));
 sky130_fd_sc_hd__xnor2_1 _5388_ (.A(_2277_),
    .B(_2278_),
    .Y(_2279_));
 sky130_fd_sc_hd__xnor2_1 _5389_ (.A(_2276_),
    .B(_2279_),
    .Y(_2280_));
 sky130_fd_sc_hd__nand2_1 _5390_ (.A(\z80.tv80s.i_tv80_core.F[1] ),
    .B(_1145_),
    .Y(_2281_));
 sky130_fd_sc_hd__o211a_1 _5391_ (.A1(\z80.tv80s.i_tv80_core.F[1] ),
    .A2(_1041_),
    .B1(_1043_),
    .C1(_2281_),
    .X(_2282_));
 sky130_fd_sc_hd__nor2_1 _5392_ (.A(_2280_),
    .B(_2282_),
    .Y(_2283_));
 sky130_fd_sc_hd__a21o_1 _5393_ (.A1(_2280_),
    .A2(_2282_),
    .B1(_0790_),
    .X(_2284_));
 sky130_fd_sc_hd__xor2_1 _5394_ (.A(_1084_),
    .B(_1156_),
    .X(_2285_));
 sky130_fd_sc_hd__xor2_1 _5395_ (.A(_0793_),
    .B(_0830_),
    .X(_2286_));
 sky130_fd_sc_hd__xor2_1 _5396_ (.A(_0912_),
    .B(_0959_),
    .X(_2287_));
 sky130_fd_sc_hd__xor2_1 _5397_ (.A(_0979_),
    .B(_1053_),
    .X(_2288_));
 sky130_fd_sc_hd__xnor2_1 _5398_ (.A(_2287_),
    .B(_2288_),
    .Y(_2289_));
 sky130_fd_sc_hd__xnor2_1 _5399_ (.A(_2286_),
    .B(_2289_),
    .Y(_2290_));
 sky130_fd_sc_hd__nor2_1 _5400_ (.A(_2285_),
    .B(_2290_),
    .Y(_2291_));
 sky130_fd_sc_hd__a21o_1 _5401_ (.A1(_2285_),
    .A2(_2290_),
    .B1(net168),
    .X(_2292_));
 sky130_fd_sc_hd__o22a_1 _5402_ (.A1(_2707_),
    .A2(\z80.tv80s.i_tv80_core.F[2] ),
    .B1(_2291_),
    .B2(_2292_),
    .X(_2293_));
 sky130_fd_sc_hd__xor2_1 _5403_ (.A(_0911_),
    .B(_0958_),
    .X(_2294_));
 sky130_fd_sc_hd__xor2_1 _5404_ (.A(_0788_),
    .B(_0829_),
    .X(_2295_));
 sky130_fd_sc_hd__xnor2_1 _5405_ (.A(_2294_),
    .B(_2295_),
    .Y(_2296_));
 sky130_fd_sc_hd__xnor2_1 _5406_ (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .B(\z80.tv80s.i_tv80_core.BusA[5] ),
    .Y(_2297_));
 sky130_fd_sc_hd__xnor2_1 _5407_ (.A(_1138_),
    .B(_2297_),
    .Y(_2298_));
 sky130_fd_sc_hd__nor2_1 _5408_ (.A(_2296_),
    .B(_2298_),
    .Y(_2299_));
 sky130_fd_sc_hd__a211o_1 _5409_ (.A1(_2296_),
    .A2(_2298_),
    .B1(_2299_),
    .C1(_0787_),
    .X(_2300_));
 sky130_fd_sc_hd__o2111ai_1 _5410_ (.A1(_2709_),
    .A2(_1988_),
    .B1(_2006_),
    .C1(_2222_),
    .D1(_2300_),
    .Y(_2301_));
 sky130_fd_sc_hd__a21oi_1 _5411_ (.A1(_0791_),
    .A2(_2293_),
    .B1(_2301_),
    .Y(_2302_));
 sky130_fd_sc_hd__o21ai_1 _5412_ (.A1(_2283_),
    .A2(_2284_),
    .B1(_2302_),
    .Y(_2303_));
 sky130_fd_sc_hd__o22a_1 _5413_ (.A1(_2222_),
    .A2(_2260_),
    .B1(_2273_),
    .B2(_2303_),
    .X(_2304_));
 sky130_fd_sc_hd__nor2_1 _5414_ (.A(_2253_),
    .B(_2304_),
    .Y(_2305_));
 sky130_fd_sc_hd__xnor2_1 _5415_ (.A(\z80.tv80s.di_reg[3] ),
    .B(\z80.tv80s.di_reg[2] ),
    .Y(_2306_));
 sky130_fd_sc_hd__xor2_1 _5416_ (.A(\z80.tv80s.di_reg[7] ),
    .B(\z80.tv80s.di_reg[6] ),
    .X(_2307_));
 sky130_fd_sc_hd__xnor2_1 _5417_ (.A(_2306_),
    .B(_2307_),
    .Y(_2308_));
 sky130_fd_sc_hd__or2_1 _5418_ (.A(\z80.tv80s.di_reg[5] ),
    .B(\z80.tv80s.di_reg[4] ),
    .X(_2309_));
 sky130_fd_sc_hd__nand2_1 _5419_ (.A(\z80.tv80s.di_reg[5] ),
    .B(\z80.tv80s.di_reg[4] ),
    .Y(_2310_));
 sky130_fd_sc_hd__nand2_1 _5420_ (.A(_2309_),
    .B(_2310_),
    .Y(_2311_));
 sky130_fd_sc_hd__xnor2_1 _5421_ (.A(\z80.tv80s.di_reg[1] ),
    .B(\z80.tv80s.di_reg[0] ),
    .Y(_2312_));
 sky130_fd_sc_hd__xnor2_1 _5422_ (.A(_2311_),
    .B(_2312_),
    .Y(_2313_));
 sky130_fd_sc_hd__xnor2_1 _5423_ (.A(_2308_),
    .B(_2313_),
    .Y(_2314_));
 sky130_fd_sc_hd__nor3_2 _5424_ (.A(_2840_),
    .B(net106),
    .C(_0587_),
    .Y(_2315_));
 sky130_fd_sc_hd__a211o_1 _5425_ (.A1(_2253_),
    .A2(_2314_),
    .B1(_2315_),
    .C1(_2305_),
    .X(_2316_));
 sky130_fd_sc_hd__nand2_1 _5426_ (.A(net485),
    .B(_2315_),
    .Y(_2317_));
 sky130_fd_sc_hd__a21oi_1 _5427_ (.A1(_2316_),
    .A2(_2317_),
    .B1(_2219_),
    .Y(_2318_));
 sky130_fd_sc_hd__o21ai_1 _5428_ (.A1(_0921_),
    .A2(_2220_),
    .B1(net112),
    .Y(_2319_));
 sky130_fd_sc_hd__o22a_1 _5429_ (.A1(net784),
    .A2(net112),
    .B1(_2318_),
    .B2(_2319_),
    .X(_0284_));
 sky130_fd_sc_hd__a21oi_1 _5430_ (.A1(\z80.tv80s.i_tv80_core.F[3] ),
    .A2(_2243_),
    .B1(_2246_),
    .Y(_2320_));
 sky130_fd_sc_hd__a21oi_1 _5431_ (.A1(_2738_),
    .A2(_0518_),
    .B1(_2320_),
    .Y(_2321_));
 sky130_fd_sc_hd__o211a_1 _5432_ (.A1(\z80.tv80s.i_tv80_core.F[3] ),
    .A2(_2244_),
    .B1(_2245_),
    .C1(_2738_),
    .X(_2322_));
 sky130_fd_sc_hd__or3_1 _5433_ (.A(_2232_),
    .B(_2321_),
    .C(_2322_),
    .X(_2323_));
 sky130_fd_sc_hd__o211a_1 _5434_ (.A1(\z80.tv80s.i_tv80_core.Fp[3] ),
    .A2(_2233_),
    .B1(_2323_),
    .C1(net101),
    .X(_2324_));
 sky130_fd_sc_hd__a211o_1 _5435_ (.A1(net621),
    .A2(net103),
    .B1(_2222_),
    .C1(_2324_),
    .X(_2325_));
 sky130_fd_sc_hd__mux2_1 _5436_ (.A0(net790),
    .A1(_0951_),
    .S(_0669_),
    .X(_2326_));
 sky130_fd_sc_hd__a311o_1 _5437_ (.A1(net627),
    .A2(_2860_),
    .A3(_0785_),
    .B1(_0960_),
    .C1(_0961_),
    .X(_2327_));
 sky130_fd_sc_hd__a221o_1 _5438_ (.A1(\z80.tv80s.i_tv80_core.F[3] ),
    .A2(_1987_),
    .B1(_2326_),
    .B2(_2722_),
    .C1(_2221_),
    .X(_2328_));
 sky130_fd_sc_hd__o211ai_1 _5439_ (.A1(_2327_),
    .A2(_2328_),
    .B1(_2254_),
    .C1(_2325_),
    .Y(_2329_));
 sky130_fd_sc_hd__o211a_1 _5440_ (.A1(_0965_),
    .A2(_2254_),
    .B1(_2329_),
    .C1(_2220_),
    .X(_2330_));
 sky130_fd_sc_hd__a21o_1 _5441_ (.A1(_0967_),
    .A2(_2219_),
    .B1(net158),
    .X(_2331_));
 sky130_fd_sc_hd__a2bb2o_1 _5442_ (.A1_N(_2330_),
    .A2_N(_2331_),
    .B1(net158),
    .B2(net621),
    .X(_0285_));
 sky130_fd_sc_hd__a211o_1 _5443_ (.A1(_0518_),
    .A2(_2236_),
    .B1(_2244_),
    .C1(\z80.tv80s.i_tv80_core.F[4] ),
    .X(_2332_));
 sky130_fd_sc_hd__a21boi_1 _5444_ (.A1(_1388_),
    .A2(_2237_),
    .B1_N(_2332_),
    .Y(_2333_));
 sky130_fd_sc_hd__nand2_1 _5445_ (.A(_2730_),
    .B(net103),
    .Y(_2334_));
 sky130_fd_sc_hd__o22a_1 _5446_ (.A1(net731),
    .A2(_2234_),
    .B1(_2333_),
    .B2(_2232_),
    .X(_2335_));
 sky130_fd_sc_hd__a31o_1 _5447_ (.A1(_2249_),
    .A2(_2334_),
    .A3(_2335_),
    .B1(_2222_),
    .X(_2336_));
 sky130_fd_sc_hd__nor2_1 _5448_ (.A(_0988_),
    .B(_1986_),
    .Y(_2337_));
 sky130_fd_sc_hd__a221o_1 _5449_ (.A1(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .A2(_0770_),
    .B1(_0988_),
    .B2(_2226_),
    .C1(_2337_),
    .X(_2338_));
 sky130_fd_sc_hd__a2bb2o_1 _5450_ (.A1_N(_0790_),
    .A2_N(_0974_),
    .B1(_1987_),
    .B2(\z80.tv80s.i_tv80_core.F[4] ),
    .X(_2339_));
 sky130_fd_sc_hd__a2111o_1 _5451_ (.A1(_2722_),
    .A2(_2338_),
    .B1(_2339_),
    .C1(_0785_),
    .D1(_2221_),
    .X(_2340_));
 sky130_fd_sc_hd__a32o_1 _5452_ (.A1(_2255_),
    .A2(_2336_),
    .A3(_2340_),
    .B1(_2219_),
    .B2(_0999_),
    .X(_2341_));
 sky130_fd_sc_hd__mux2_1 _5453_ (.A0(net833),
    .A1(_2341_),
    .S(net112),
    .X(_0286_));
 sky130_fd_sc_hd__a21oi_1 _5454_ (.A1(\z80.tv80s.i_tv80_core.F[5] ),
    .A2(_2243_),
    .B1(_2246_),
    .Y(_2342_));
 sky130_fd_sc_hd__a21oi_1 _5455_ (.A1(_2739_),
    .A2(_0518_),
    .B1(_2342_),
    .Y(_2343_));
 sky130_fd_sc_hd__o211a_1 _5456_ (.A1(\z80.tv80s.i_tv80_core.F[5] ),
    .A2(_2244_),
    .B1(_2245_),
    .C1(_2739_),
    .X(_2344_));
 sky130_fd_sc_hd__or3_1 _5457_ (.A(_2232_),
    .B(_2343_),
    .C(_2344_),
    .X(_2345_));
 sky130_fd_sc_hd__o211a_1 _5458_ (.A1(\z80.tv80s.i_tv80_core.Fp[5] ),
    .A2(_2233_),
    .B1(_2345_),
    .C1(net101),
    .X(_2346_));
 sky130_fd_sc_hd__a211o_1 _5459_ (.A1(net793),
    .A2(_0540_),
    .B1(_2222_),
    .C1(_2346_),
    .X(_2347_));
 sky130_fd_sc_hd__mux2_1 _5460_ (.A0(\z80.tv80s.i_tv80_core.BusB[5] ),
    .A1(_1038_),
    .S(_0669_),
    .X(_2348_));
 sky130_fd_sc_hd__a311o_1 _5461_ (.A1(\z80.tv80s.i_tv80_core.BusB[5] ),
    .A2(_2860_),
    .A3(_0785_),
    .B1(_1052_),
    .C1(_1054_),
    .X(_2349_));
 sky130_fd_sc_hd__a221o_1 _5462_ (.A1(\z80.tv80s.i_tv80_core.F[5] ),
    .A2(_1987_),
    .B1(_2348_),
    .B2(_2722_),
    .C1(_2349_),
    .X(_2350_));
 sky130_fd_sc_hd__o21a_1 _5463_ (.A1(_2221_),
    .A2(_2350_),
    .B1(_2254_),
    .X(_2351_));
 sky130_fd_sc_hd__a2bb2o_1 _5464_ (.A1_N(_0842_),
    .A2_N(_2254_),
    .B1(_2347_),
    .B2(_2351_),
    .X(_2352_));
 sky130_fd_sc_hd__mux2_1 _5465_ (.A0(_1060_),
    .A1(_2352_),
    .S(_2220_),
    .X(_2353_));
 sky130_fd_sc_hd__mux2_1 _5466_ (.A0(net793),
    .A1(_2353_),
    .S(net112),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _5467_ (.A0(\z80.tv80s.i_tv80_core.Fp[6] ),
    .A1(\z80.tv80s.i_tv80_core.F[6] ),
    .S(_2234_),
    .X(_2354_));
 sky130_fd_sc_hd__or4_1 _5468_ (.A(\z80.tv80s.i_tv80_core.I[5] ),
    .B(\z80.tv80s.i_tv80_core.I[4] ),
    .C(\z80.tv80s.i_tv80_core.I[7] ),
    .D(\z80.tv80s.i_tv80_core.I[6] ),
    .X(_2355_));
 sky130_fd_sc_hd__or4_1 _5469_ (.A(\z80.tv80s.i_tv80_core.I[1] ),
    .B(\z80.tv80s.i_tv80_core.I[0] ),
    .C(\z80.tv80s.i_tv80_core.I[3] ),
    .D(\z80.tv80s.i_tv80_core.I[2] ),
    .X(_2356_));
 sky130_fd_sc_hd__o21ai_1 _5470_ (.A1(_2355_),
    .A2(_2356_),
    .B1(_2248_),
    .Y(_2357_));
 sky130_fd_sc_hd__o211a_1 _5471_ (.A1(_2248_),
    .A2(_2354_),
    .B1(_2357_),
    .C1(_2221_),
    .X(_2358_));
 sky130_fd_sc_hd__o21ba_1 _5472_ (.A1(_2011_),
    .A2(_2221_),
    .B1_N(_2358_),
    .X(_2359_));
 sky130_fd_sc_hd__or4_1 _5473_ (.A(\z80.tv80s.di_reg[3] ),
    .B(\z80.tv80s.di_reg[2] ),
    .C(\z80.tv80s.di_reg[7] ),
    .D(\z80.tv80s.di_reg[6] ),
    .X(_2360_));
 sky130_fd_sc_hd__or4_1 _5474_ (.A(\z80.tv80s.di_reg[1] ),
    .B(\z80.tv80s.di_reg[0] ),
    .C(_2309_),
    .D(_2360_),
    .X(_2361_));
 sky130_fd_sc_hd__mux2_1 _5475_ (.A0(_2359_),
    .A1(_2361_),
    .S(_2253_),
    .X(_2362_));
 sky130_fd_sc_hd__mux2_1 _5476_ (.A0(_1091_),
    .A1(_2362_),
    .S(_2220_),
    .X(_2363_));
 sky130_fd_sc_hd__inv_2 _5477_ (.A(_2363_),
    .Y(_2364_));
 sky130_fd_sc_hd__mux2_1 _5478_ (.A0(net823),
    .A1(_2364_),
    .S(net112),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _5479_ (.A0(\z80.tv80s.i_tv80_core.F[7] ),
    .A1(_1136_),
    .S(_2731_),
    .X(_2365_));
 sky130_fd_sc_hd__mux2_1 _5480_ (.A0(\z80.tv80s.i_tv80_core.F[7] ),
    .A1(_1156_),
    .S(_2707_),
    .X(_2366_));
 sky130_fd_sc_hd__a221o_1 _5481_ (.A1(\z80.tv80s.i_tv80_core.F[7] ),
    .A2(_1987_),
    .B1(_2366_),
    .B2(_0791_),
    .C1(_2221_),
    .X(_2367_));
 sky130_fd_sc_hd__a211o_1 _5482_ (.A1(_2722_),
    .A2(_2365_),
    .B1(_2367_),
    .C1(_1151_),
    .X(_2368_));
 sky130_fd_sc_hd__mux2_1 _5483_ (.A0(\z80.tv80s.i_tv80_core.Fp[7] ),
    .A1(\z80.tv80s.i_tv80_core.F[7] ),
    .S(_2234_),
    .X(_2369_));
 sky130_fd_sc_hd__mux2_1 _5484_ (.A0(_2369_),
    .A1(net578),
    .S(_2248_),
    .X(_2370_));
 sky130_fd_sc_hd__o21a_1 _5485_ (.A1(_2222_),
    .A2(_2370_),
    .B1(_2252_),
    .X(_2371_));
 sky130_fd_sc_hd__a22o_1 _5486_ (.A1(\z80.tv80s.di_reg[7] ),
    .A2(_2253_),
    .B1(_2368_),
    .B2(_2371_),
    .X(_2372_));
 sky130_fd_sc_hd__mux2_1 _5487_ (.A0(_1162_),
    .A1(_2372_),
    .S(_2220_),
    .X(_2373_));
 sky130_fd_sc_hd__mux2_1 _5488_ (.A0(net818),
    .A1(_2373_),
    .S(net112),
    .X(_0289_));
 sky130_fd_sc_hd__nand4_4 _5489_ (.A(\z80.tv80s.i_tv80_core.ts[3] ),
    .B(_2786_),
    .C(_2854_),
    .D(_0561_),
    .Y(_2374_));
 sky130_fd_sc_hd__mux2_1 _5490_ (.A0(\z80.tv80s.i_tv80_core.ACC[0] ),
    .A1(net588),
    .S(_2374_),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _5491_ (.A0(\z80.tv80s.i_tv80_core.ACC[1] ),
    .A1(net629),
    .S(_2374_),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_1 _5492_ (.A0(\z80.tv80s.i_tv80_core.ACC[2] ),
    .A1(net566),
    .S(_2374_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _5493_ (.A0(\z80.tv80s.i_tv80_core.ACC[3] ),
    .A1(net615),
    .S(_2374_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _5494_ (.A0(\z80.tv80s.i_tv80_core.ACC[4] ),
    .A1(net644),
    .S(_2374_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _5495_ (.A0(\z80.tv80s.i_tv80_core.ACC[5] ),
    .A1(net597),
    .S(_2374_),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _5496_ (.A0(\z80.tv80s.i_tv80_core.ACC[6] ),
    .A1(net549),
    .S(_2374_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _5497_ (.A0(\z80.tv80s.i_tv80_core.ACC[7] ),
    .A1(net578),
    .S(_2374_),
    .X(_0297_));
 sky130_fd_sc_hd__or3_2 _5498_ (.A(net619),
    .B(_0423_),
    .C(_0664_),
    .X(_2375_));
 sky130_fd_sc_hd__o31a_1 _5499_ (.A1(net67),
    .A2(_1738_),
    .A3(_2375_),
    .B1(net103),
    .X(_2376_));
 sky130_fd_sc_hd__a211oi_4 _5500_ (.A1(net103),
    .A2(_0546_),
    .B1(_2376_),
    .C1(net155),
    .Y(_2377_));
 sky130_fd_sc_hd__a31o_1 _5501_ (.A1(_2708_),
    .A2(_2896_),
    .A3(_0385_),
    .B1(net164),
    .X(_2378_));
 sky130_fd_sc_hd__or4_1 _5502_ (.A(net115),
    .B(_2773_),
    .C(_2781_),
    .D(_2878_),
    .X(_2379_));
 sky130_fd_sc_hd__o31a_1 _5503_ (.A1(_2914_),
    .A2(_2943_),
    .A3(_2379_),
    .B1(_0385_),
    .X(_2380_));
 sky130_fd_sc_hd__o31a_1 _5504_ (.A1(_2763_),
    .A2(_0495_),
    .A3(_1446_),
    .B1(net146),
    .X(_2381_));
 sky130_fd_sc_hd__a32o_1 _5505_ (.A1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .A2(_0556_),
    .A3(_0616_),
    .B1(_0430_),
    .B2(_0497_),
    .X(_2382_));
 sky130_fd_sc_hd__o31a_1 _5506_ (.A1(_2380_),
    .A2(_2381_),
    .A3(_2382_),
    .B1(_2378_),
    .X(_2383_));
 sky130_fd_sc_hd__nand2_4 _5507_ (.A(net168),
    .B(_0613_),
    .Y(_2384_));
 sky130_fd_sc_hd__a21o_2 _5508_ (.A1(net168),
    .A2(_0613_),
    .B1(net269),
    .X(_2385_));
 sky130_fd_sc_hd__a21oi_1 _5509_ (.A1(_2708_),
    .A2(_0374_),
    .B1(_2697_),
    .Y(_2386_));
 sky130_fd_sc_hd__o41a_2 _5510_ (.A1(net555),
    .A2(_2383_),
    .A3(_2385_),
    .A4(_2386_),
    .B1(_0545_),
    .X(_2387_));
 sky130_fd_sc_hd__or2_2 _5511_ (.A(net102),
    .B(_2387_),
    .X(_2388_));
 sky130_fd_sc_hd__o21ai_2 _5512_ (.A1(_2733_),
    .A2(_2384_),
    .B1(_2385_),
    .Y(_2389_));
 sky130_fd_sc_hd__nand2_1 _5513_ (.A(\z80.tv80s.i_tv80_core.PC[0] ),
    .B(_2389_),
    .Y(_2390_));
 sky130_fd_sc_hd__xor2_1 _5514_ (.A(net748),
    .B(_2389_),
    .X(_2391_));
 sky130_fd_sc_hd__mux2_1 _5515_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .A1(\z80.tv80s.i_tv80_core.PC[0] ),
    .S(net98),
    .X(_2392_));
 sky130_fd_sc_hd__a22o_1 _5516_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .A2(net63),
    .B1(net60),
    .B2(_2392_),
    .X(_2393_));
 sky130_fd_sc_hd__a21bo_1 _5517_ (.A1(net86),
    .A2(_2393_),
    .B1_N(_1735_),
    .X(_2394_));
 sky130_fd_sc_hd__mux2_1 _5518_ (.A0(_2394_),
    .A1(net744),
    .S(net67),
    .X(_2395_));
 sky130_fd_sc_hd__mux2_1 _5519_ (.A0(_2395_),
    .A1(net748),
    .S(net54),
    .X(_2396_));
 sky130_fd_sc_hd__mux2_1 _5520_ (.A0(_2396_),
    .A1(_2391_),
    .S(net62),
    .X(_2397_));
 sky130_fd_sc_hd__mux2_1 _5521_ (.A0(net748),
    .A1(_2397_),
    .S(net59),
    .X(_0298_));
 sky130_fd_sc_hd__o21ai_1 _5522_ (.A1(\z80.tv80s.di_reg[1] ),
    .A2(_2384_),
    .B1(_2385_),
    .Y(_2398_));
 sky130_fd_sc_hd__nor2_1 _5523_ (.A(_2740_),
    .B(_2398_),
    .Y(_2399_));
 sky130_fd_sc_hd__xnor2_1 _5524_ (.A(_2740_),
    .B(_2398_),
    .Y(_2400_));
 sky130_fd_sc_hd__nor2_1 _5525_ (.A(_2390_),
    .B(_2400_),
    .Y(_2401_));
 sky130_fd_sc_hd__and2_1 _5526_ (.A(_2390_),
    .B(_2400_),
    .X(_2402_));
 sky130_fd_sc_hd__nor2_1 _5527_ (.A(_2401_),
    .B(_2402_),
    .Y(_2403_));
 sky130_fd_sc_hd__a21o_1 _5528_ (.A1(\z80.tv80s.i_tv80_core.PC[1] ),
    .A2(net98),
    .B1(_1767_),
    .X(_2404_));
 sky130_fd_sc_hd__mux2_1 _5529_ (.A0(_2404_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .S(net63),
    .X(_2405_));
 sky130_fd_sc_hd__a21bo_1 _5530_ (.A1(net86),
    .A2(_2405_),
    .B1_N(_1766_),
    .X(_2406_));
 sky130_fd_sc_hd__mux2_1 _5531_ (.A0(_2406_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .S(net67),
    .X(_2407_));
 sky130_fd_sc_hd__mux2_1 _5532_ (.A0(_2407_),
    .A1(net729),
    .S(net54),
    .X(_2408_));
 sky130_fd_sc_hd__mux2_1 _5533_ (.A0(_2408_),
    .A1(_2403_),
    .S(net62),
    .X(_2409_));
 sky130_fd_sc_hd__mux2_1 _5534_ (.A0(net729),
    .A1(_2409_),
    .S(net59),
    .X(_0299_));
 sky130_fd_sc_hd__o21ai_1 _5535_ (.A1(\z80.tv80s.di_reg[2] ),
    .A2(_2384_),
    .B1(_2385_),
    .Y(_2410_));
 sky130_fd_sc_hd__nor2_1 _5536_ (.A(_2741_),
    .B(_2410_),
    .Y(_2411_));
 sky130_fd_sc_hd__inv_2 _5537_ (.A(_2411_),
    .Y(_2412_));
 sky130_fd_sc_hd__xnor2_1 _5538_ (.A(_2741_),
    .B(_2410_),
    .Y(_2413_));
 sky130_fd_sc_hd__o21bai_1 _5539_ (.A1(_2399_),
    .A2(_2401_),
    .B1_N(_2413_),
    .Y(_2414_));
 sky130_fd_sc_hd__or3b_1 _5540_ (.A(_2399_),
    .B(_2401_),
    .C_N(_2413_),
    .X(_2415_));
 sky130_fd_sc_hd__a21o_1 _5541_ (.A1(\z80.tv80s.i_tv80_core.PC[2] ),
    .A2(net98),
    .B1(_1782_),
    .X(_2416_));
 sky130_fd_sc_hd__mux2_1 _5542_ (.A0(_2416_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .S(net63),
    .X(_2417_));
 sky130_fd_sc_hd__a21bo_1 _5543_ (.A1(net86),
    .A2(_2417_),
    .B1_N(_1781_),
    .X(_2418_));
 sky130_fd_sc_hd__mux2_1 _5544_ (.A0(_2418_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .S(net67),
    .X(_2419_));
 sky130_fd_sc_hd__a21oi_1 _5545_ (.A1(_2741_),
    .A2(net54),
    .B1(net62),
    .Y(_2420_));
 sky130_fd_sc_hd__o21a_1 _5546_ (.A1(net54),
    .A2(_2419_),
    .B1(_2420_),
    .X(_2421_));
 sky130_fd_sc_hd__a31o_1 _5547_ (.A1(net62),
    .A2(_2414_),
    .A3(_2415_),
    .B1(_2421_),
    .X(_2422_));
 sky130_fd_sc_hd__mux2_1 _5548_ (.A0(net609),
    .A1(_2422_),
    .S(net59),
    .X(_0300_));
 sky130_fd_sc_hd__o21ai_1 _5549_ (.A1(\z80.tv80s.di_reg[3] ),
    .A2(_2384_),
    .B1(_2385_),
    .Y(_2423_));
 sky130_fd_sc_hd__nor2_1 _5550_ (.A(_2742_),
    .B(_2423_),
    .Y(_2424_));
 sky130_fd_sc_hd__xnor2_1 _5551_ (.A(_2742_),
    .B(_2423_),
    .Y(_2425_));
 sky130_fd_sc_hd__and3_1 _5552_ (.A(_2412_),
    .B(_2414_),
    .C(_2425_),
    .X(_2426_));
 sky130_fd_sc_hd__a21oi_1 _5553_ (.A1(_2412_),
    .A2(_2414_),
    .B1(_2425_),
    .Y(_2427_));
 sky130_fd_sc_hd__mux2_1 _5554_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .A1(\z80.tv80s.i_tv80_core.PC[3] ),
    .S(net98),
    .X(_2428_));
 sky130_fd_sc_hd__a22o_1 _5555_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .A2(net63),
    .B1(net60),
    .B2(_2428_),
    .X(_2429_));
 sky130_fd_sc_hd__a21bo_1 _5556_ (.A1(net86),
    .A2(_2429_),
    .B1_N(_1796_),
    .X(_2430_));
 sky130_fd_sc_hd__mux2_1 _5557_ (.A0(_2430_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .S(net67),
    .X(_2431_));
 sky130_fd_sc_hd__mux2_1 _5558_ (.A0(_2431_),
    .A1(net642),
    .S(net55),
    .X(_2432_));
 sky130_fd_sc_hd__nor2_1 _5559_ (.A(_2426_),
    .B(_2427_),
    .Y(_2433_));
 sky130_fd_sc_hd__mux2_1 _5560_ (.A0(_2432_),
    .A1(_2433_),
    .S(net62),
    .X(_2434_));
 sky130_fd_sc_hd__mux2_1 _5561_ (.A0(net642),
    .A1(_2434_),
    .S(net59),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _5562_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .A1(\z80.tv80s.i_tv80_core.PC[4] ),
    .S(net98),
    .X(_2435_));
 sky130_fd_sc_hd__a22o_1 _5563_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .A2(net63),
    .B1(net60),
    .B2(_2435_),
    .X(_2436_));
 sky130_fd_sc_hd__a21bo_1 _5564_ (.A1(net86),
    .A2(_2436_),
    .B1_N(_1810_),
    .X(_2437_));
 sky130_fd_sc_hd__mux2_1 _5565_ (.A0(_2437_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .S(net67),
    .X(_2438_));
 sky130_fd_sc_hd__mux2_1 _5566_ (.A0(_2438_),
    .A1(net648),
    .S(net54),
    .X(_2439_));
 sky130_fd_sc_hd__o21ai_1 _5567_ (.A1(\z80.tv80s.di_reg[4] ),
    .A2(_2384_),
    .B1(_2385_),
    .Y(_2440_));
 sky130_fd_sc_hd__nor2_1 _5568_ (.A(_2743_),
    .B(_2440_),
    .Y(_2441_));
 sky130_fd_sc_hd__xnor2_1 _5569_ (.A(_2743_),
    .B(_2440_),
    .Y(_2442_));
 sky130_fd_sc_hd__o21ba_1 _5570_ (.A1(_2424_),
    .A2(_2427_),
    .B1_N(_2442_),
    .X(_2443_));
 sky130_fd_sc_hd__or3b_1 _5571_ (.A(_2424_),
    .B(_2427_),
    .C_N(_2442_),
    .X(_2444_));
 sky130_fd_sc_hd__and2b_1 _5572_ (.A_N(_2443_),
    .B(_2444_),
    .X(_2445_));
 sky130_fd_sc_hd__mux2_1 _5573_ (.A0(_2439_),
    .A1(_2445_),
    .S(net62),
    .X(_2446_));
 sky130_fd_sc_hd__mux2_1 _5574_ (.A0(net648),
    .A1(_2446_),
    .S(net59),
    .X(_0302_));
 sky130_fd_sc_hd__a21o_1 _5575_ (.A1(\z80.tv80s.i_tv80_core.PC[5] ),
    .A2(net98),
    .B1(_1824_),
    .X(_2447_));
 sky130_fd_sc_hd__mux2_1 _5576_ (.A0(_2447_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .S(net63),
    .X(_2448_));
 sky130_fd_sc_hd__a21bo_1 _5577_ (.A1(net86),
    .A2(_2448_),
    .B1_N(_1823_),
    .X(_2449_));
 sky130_fd_sc_hd__mux2_1 _5578_ (.A0(_2449_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .S(net67),
    .X(_2450_));
 sky130_fd_sc_hd__mux2_1 _5579_ (.A0(_2450_),
    .A1(net638),
    .S(net55),
    .X(_2451_));
 sky130_fd_sc_hd__o21ai_1 _5580_ (.A1(\z80.tv80s.di_reg[5] ),
    .A2(_2384_),
    .B1(_2385_),
    .Y(_2452_));
 sky130_fd_sc_hd__nor2_1 _5581_ (.A(_2744_),
    .B(_2452_),
    .Y(_2453_));
 sky130_fd_sc_hd__xnor2_1 _5582_ (.A(_2744_),
    .B(_2452_),
    .Y(_2454_));
 sky130_fd_sc_hd__o21ba_1 _5583_ (.A1(_2441_),
    .A2(_2443_),
    .B1_N(_2454_),
    .X(_2455_));
 sky130_fd_sc_hd__or3b_1 _5584_ (.A(_2441_),
    .B(_2443_),
    .C_N(_2454_),
    .X(_2456_));
 sky130_fd_sc_hd__and2b_1 _5585_ (.A_N(_2455_),
    .B(_2456_),
    .X(_2457_));
 sky130_fd_sc_hd__mux2_1 _5586_ (.A0(_2451_),
    .A1(_2457_),
    .S(net62),
    .X(_2458_));
 sky130_fd_sc_hd__mux2_1 _5587_ (.A0(net638),
    .A1(_2458_),
    .S(net59),
    .X(_0303_));
 sky130_fd_sc_hd__o21ai_1 _5588_ (.A1(\z80.tv80s.di_reg[6] ),
    .A2(_2384_),
    .B1(_2385_),
    .Y(_2459_));
 sky130_fd_sc_hd__nor2_1 _5589_ (.A(_2745_),
    .B(_2459_),
    .Y(_2460_));
 sky130_fd_sc_hd__xnor2_1 _5590_ (.A(_2745_),
    .B(_2459_),
    .Y(_2461_));
 sky130_fd_sc_hd__o21ba_1 _5591_ (.A1(_2453_),
    .A2(_2455_),
    .B1_N(_2461_),
    .X(_2462_));
 sky130_fd_sc_hd__or3b_1 _5592_ (.A(_2453_),
    .B(_2455_),
    .C_N(_2461_),
    .X(_2463_));
 sky130_fd_sc_hd__and2b_1 _5593_ (.A_N(_2462_),
    .B(_2463_),
    .X(_2464_));
 sky130_fd_sc_hd__a21o_1 _5594_ (.A1(\z80.tv80s.i_tv80_core.PC[6] ),
    .A2(net98),
    .B1(_1838_),
    .X(_2465_));
 sky130_fd_sc_hd__mux2_1 _5595_ (.A0(_2465_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .S(net63),
    .X(_2466_));
 sky130_fd_sc_hd__a21bo_1 _5596_ (.A1(net86),
    .A2(_2466_),
    .B1_N(_1837_),
    .X(_2467_));
 sky130_fd_sc_hd__mux2_1 _5597_ (.A0(_2467_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .S(net67),
    .X(_2468_));
 sky130_fd_sc_hd__mux2_1 _5598_ (.A0(_2468_),
    .A1(net631),
    .S(net55),
    .X(_2469_));
 sky130_fd_sc_hd__mux2_1 _5599_ (.A0(_2469_),
    .A1(_2464_),
    .S(net62),
    .X(_2470_));
 sky130_fd_sc_hd__mux2_1 _5600_ (.A0(net631),
    .A1(_2470_),
    .S(net59),
    .X(_0304_));
 sky130_fd_sc_hd__o21a_2 _5601_ (.A1(\z80.tv80s.di_reg[7] ),
    .A2(_2384_),
    .B1(_2385_),
    .X(_2471_));
 sky130_fd_sc_hd__xnor2_1 _5602_ (.A(net677),
    .B(net76),
    .Y(_2472_));
 sky130_fd_sc_hd__o21ba_1 _5603_ (.A1(_2460_),
    .A2(_2462_),
    .B1_N(_2472_),
    .X(_2473_));
 sky130_fd_sc_hd__or3b_1 _5604_ (.A(_2460_),
    .B(_2462_),
    .C_N(_2472_),
    .X(_2474_));
 sky130_fd_sc_hd__and2b_1 _5605_ (.A_N(_2473_),
    .B(_2474_),
    .X(_2475_));
 sky130_fd_sc_hd__mux2_1 _5606_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .A1(\z80.tv80s.i_tv80_core.PC[7] ),
    .S(net98),
    .X(_2476_));
 sky130_fd_sc_hd__a22o_1 _5607_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .A2(net63),
    .B1(net60),
    .B2(_2476_),
    .X(_2477_));
 sky130_fd_sc_hd__a21bo_1 _5608_ (.A1(net87),
    .A2(_2477_),
    .B1_N(_1850_),
    .X(_2478_));
 sky130_fd_sc_hd__mux2_1 _5609_ (.A0(_2478_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .S(net67),
    .X(_2479_));
 sky130_fd_sc_hd__mux2_1 _5610_ (.A0(_2479_),
    .A1(net677),
    .S(net55),
    .X(_2480_));
 sky130_fd_sc_hd__mux2_1 _5611_ (.A0(_2480_),
    .A1(_2475_),
    .S(net62),
    .X(_2481_));
 sky130_fd_sc_hd__mux2_1 _5612_ (.A0(net677),
    .A1(_2481_),
    .S(net59),
    .X(_0305_));
 sky130_fd_sc_hd__xnor2_1 _5613_ (.A(net778),
    .B(net76),
    .Y(_2482_));
 sky130_fd_sc_hd__a21o_1 _5614_ (.A1(net677),
    .A2(net76),
    .B1(_2473_),
    .X(_2483_));
 sky130_fd_sc_hd__and2b_1 _5615_ (.A_N(_2482_),
    .B(_2483_),
    .X(_2484_));
 sky130_fd_sc_hd__xnor2_1 _5616_ (.A(_2482_),
    .B(_2483_),
    .Y(_2485_));
 sky130_fd_sc_hd__mux2_1 _5617_ (.A0(\z80.tv80s.i_tv80_core.I[0] ),
    .A1(\z80.tv80s.i_tv80_core.PC[8] ),
    .S(net99),
    .X(_2486_));
 sky130_fd_sc_hd__a22o_1 _5618_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .A2(net64),
    .B1(net61),
    .B2(_2486_),
    .X(_2487_));
 sky130_fd_sc_hd__a21bo_1 _5619_ (.A1(net87),
    .A2(_2487_),
    .B1_N(_1865_),
    .X(_2488_));
 sky130_fd_sc_hd__mux2_1 _5620_ (.A0(_2488_),
    .A1(\z80.tv80s.di_reg[0] ),
    .S(net68),
    .X(_2489_));
 sky130_fd_sc_hd__mux2_1 _5621_ (.A0(_2489_),
    .A1(net778),
    .S(net55),
    .X(_2490_));
 sky130_fd_sc_hd__mux2_1 _5622_ (.A0(_2490_),
    .A1(_2485_),
    .S(net62),
    .X(_2491_));
 sky130_fd_sc_hd__mux2_1 _5623_ (.A0(net778),
    .A1(_2491_),
    .S(net59),
    .X(_0306_));
 sky130_fd_sc_hd__o21a_1 _5624_ (.A1(_0518_),
    .A2(_2388_),
    .B1(net59),
    .X(_2492_));
 sky130_fd_sc_hd__o21ai_1 _5625_ (.A1(_0518_),
    .A2(net62),
    .B1(net59),
    .Y(_2493_));
 sky130_fd_sc_hd__xor2_2 _5626_ (.A(net761),
    .B(net76),
    .X(_2494_));
 sky130_fd_sc_hd__a21oi_1 _5627_ (.A1(\z80.tv80s.i_tv80_core.PC[8] ),
    .A2(net76),
    .B1(_2484_),
    .Y(_2495_));
 sky130_fd_sc_hd__xnor2_1 _5628_ (.A(_2494_),
    .B(_2495_),
    .Y(_2496_));
 sky130_fd_sc_hd__nor2_2 _5629_ (.A(_1387_),
    .B(_2387_),
    .Y(_2497_));
 sky130_fd_sc_hd__mux2_1 _5630_ (.A0(\z80.tv80s.i_tv80_core.I[1] ),
    .A1(\z80.tv80s.i_tv80_core.PC[9] ),
    .S(net99),
    .X(_2498_));
 sky130_fd_sc_hd__a22o_1 _5631_ (.A1(net671),
    .A2(net64),
    .B1(net61),
    .B2(_2498_),
    .X(_2499_));
 sky130_fd_sc_hd__a21bo_1 _5632_ (.A1(net87),
    .A2(_2499_),
    .B1_N(_1880_),
    .X(_2500_));
 sky130_fd_sc_hd__mux2_1 _5633_ (.A0(_2500_),
    .A1(\z80.tv80s.di_reg[1] ),
    .S(net68),
    .X(_2501_));
 sky130_fd_sc_hd__a22o_1 _5634_ (.A1(net62),
    .A2(_2496_),
    .B1(_2497_),
    .B2(_2501_),
    .X(_2502_));
 sky130_fd_sc_hd__a22o_1 _5635_ (.A1(net761),
    .A2(_2493_),
    .B1(_2502_),
    .B2(net59),
    .X(_0307_));
 sky130_fd_sc_hd__xnor2_1 _5636_ (.A(net753),
    .B(net76),
    .Y(_2503_));
 sky130_fd_sc_hd__o21a_1 _5637_ (.A1(\z80.tv80s.i_tv80_core.PC[8] ),
    .A2(\z80.tv80s.i_tv80_core.PC[9] ),
    .B1(net76),
    .X(_2504_));
 sky130_fd_sc_hd__a21o_1 _5638_ (.A1(_2484_),
    .A2(_2494_),
    .B1(_2504_),
    .X(_2505_));
 sky130_fd_sc_hd__and2b_1 _5639_ (.A_N(_2503_),
    .B(_2505_),
    .X(_2506_));
 sky130_fd_sc_hd__xor2_1 _5640_ (.A(_2503_),
    .B(_2505_),
    .X(_2507_));
 sky130_fd_sc_hd__mux2_1 _5641_ (.A0(\z80.tv80s.i_tv80_core.I[2] ),
    .A1(\z80.tv80s.i_tv80_core.PC[10] ),
    .S(net99),
    .X(_2508_));
 sky130_fd_sc_hd__a22o_1 _5642_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .A2(net64),
    .B1(net61),
    .B2(_2508_),
    .X(_2509_));
 sky130_fd_sc_hd__nand2_1 _5643_ (.A(net87),
    .B(_2509_),
    .Y(_2510_));
 sky130_fd_sc_hd__a21o_1 _5644_ (.A1(_1896_),
    .A2(_2510_),
    .B1(net68),
    .X(_2511_));
 sky130_fd_sc_hd__a32o_1 _5645_ (.A1(_1908_),
    .A2(_2497_),
    .A3(_2511_),
    .B1(_2507_),
    .B2(_2388_),
    .X(_2512_));
 sky130_fd_sc_hd__o2bb2a_1 _5646_ (.A1_N(net59),
    .A2_N(_2512_),
    .B1(_2492_),
    .B2(net753),
    .X(_0308_));
 sky130_fd_sc_hd__xnor2_1 _5647_ (.A(net742),
    .B(net76),
    .Y(_2513_));
 sky130_fd_sc_hd__a21o_1 _5648_ (.A1(\z80.tv80s.i_tv80_core.PC[10] ),
    .A2(net76),
    .B1(_2506_),
    .X(_2514_));
 sky130_fd_sc_hd__xnor2_1 _5649_ (.A(_2513_),
    .B(_2514_),
    .Y(_2515_));
 sky130_fd_sc_hd__mux2_1 _5650_ (.A0(\z80.tv80s.i_tv80_core.I[3] ),
    .A1(\z80.tv80s.i_tv80_core.PC[11] ),
    .S(net99),
    .X(_2516_));
 sky130_fd_sc_hd__a22o_1 _5651_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .A2(net64),
    .B1(net61),
    .B2(_2516_),
    .X(_2517_));
 sky130_fd_sc_hd__a21bo_1 _5652_ (.A1(net87),
    .A2(_2517_),
    .B1_N(_1910_),
    .X(_2518_));
 sky130_fd_sc_hd__mux2_1 _5653_ (.A0(_2518_),
    .A1(\z80.tv80s.di_reg[3] ),
    .S(net68),
    .X(_2519_));
 sky130_fd_sc_hd__mux2_1 _5654_ (.A0(_2519_),
    .A1(net742),
    .S(net55),
    .X(_2520_));
 sky130_fd_sc_hd__mux2_1 _5655_ (.A0(_2520_),
    .A1(_2515_),
    .S(net62),
    .X(_2521_));
 sky130_fd_sc_hd__mux2_1 _5656_ (.A0(net742),
    .A1(_2521_),
    .S(net59),
    .X(_0309_));
 sky130_fd_sc_hd__nand2_1 _5657_ (.A(net683),
    .B(net76),
    .Y(_2522_));
 sky130_fd_sc_hd__or2_1 _5658_ (.A(net683),
    .B(net76),
    .X(_2523_));
 sky130_fd_sc_hd__nand2_1 _5659_ (.A(_2522_),
    .B(_2523_),
    .Y(_2524_));
 sky130_fd_sc_hd__nor2_1 _5660_ (.A(_2503_),
    .B(_2513_),
    .Y(_2525_));
 sky130_fd_sc_hd__and2_1 _5661_ (.A(_2494_),
    .B(_2525_),
    .X(_2526_));
 sky130_fd_sc_hd__o41a_1 _5662_ (.A1(\z80.tv80s.i_tv80_core.PC[8] ),
    .A2(\z80.tv80s.i_tv80_core.PC[9] ),
    .A3(\z80.tv80s.i_tv80_core.PC[10] ),
    .A4(\z80.tv80s.i_tv80_core.PC[11] ),
    .B1(net76),
    .X(_2527_));
 sky130_fd_sc_hd__a21oi_1 _5663_ (.A1(_2484_),
    .A2(_2526_),
    .B1(_2527_),
    .Y(_2528_));
 sky130_fd_sc_hd__xnor2_1 _5664_ (.A(_2524_),
    .B(_2528_),
    .Y(_2529_));
 sky130_fd_sc_hd__mux2_1 _5665_ (.A0(\z80.tv80s.i_tv80_core.I[4] ),
    .A1(\z80.tv80s.i_tv80_core.PC[12] ),
    .S(net99),
    .X(_2530_));
 sky130_fd_sc_hd__a22o_1 _5666_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .A2(net64),
    .B1(net61),
    .B2(_2530_),
    .X(_2531_));
 sky130_fd_sc_hd__a21bo_1 _5667_ (.A1(net87),
    .A2(_2531_),
    .B1_N(_1925_),
    .X(_2532_));
 sky130_fd_sc_hd__mux2_1 _5668_ (.A0(_2532_),
    .A1(\z80.tv80s.di_reg[4] ),
    .S(net68),
    .X(_2533_));
 sky130_fd_sc_hd__mux2_1 _5669_ (.A0(_2533_),
    .A1(net683),
    .S(net55),
    .X(_2534_));
 sky130_fd_sc_hd__nor2_1 _5670_ (.A(net62),
    .B(_2534_),
    .Y(_2535_));
 sky130_fd_sc_hd__a21oi_1 _5671_ (.A1(net62),
    .A2(_2529_),
    .B1(_2535_),
    .Y(_2536_));
 sky130_fd_sc_hd__mux2_1 _5672_ (.A0(net683),
    .A1(_2536_),
    .S(net59),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _5673_ (.A0(net597),
    .A1(\z80.tv80s.i_tv80_core.PC[13] ),
    .S(net99),
    .X(_2537_));
 sky130_fd_sc_hd__a22o_1 _5674_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .A2(net64),
    .B1(net61),
    .B2(_2537_),
    .X(_2538_));
 sky130_fd_sc_hd__a21bo_1 _5675_ (.A1(net87),
    .A2(_2538_),
    .B1_N(_1941_),
    .X(_2539_));
 sky130_fd_sc_hd__mux2_1 _5676_ (.A0(_2539_),
    .A1(\z80.tv80s.di_reg[5] ),
    .S(net68),
    .X(_2540_));
 sky130_fd_sc_hd__and2_1 _5677_ (.A(net707),
    .B(net76),
    .X(_2541_));
 sky130_fd_sc_hd__nand2_1 _5678_ (.A(\z80.tv80s.i_tv80_core.PC[13] ),
    .B(net76),
    .Y(_2542_));
 sky130_fd_sc_hd__nor2_1 _5679_ (.A(net707),
    .B(net76),
    .Y(_2543_));
 sky130_fd_sc_hd__o21a_1 _5680_ (.A1(_2524_),
    .A2(_2528_),
    .B1(_2522_),
    .X(_2544_));
 sky130_fd_sc_hd__o21ai_1 _5681_ (.A1(_2541_),
    .A2(_2543_),
    .B1(_2544_),
    .Y(_2545_));
 sky130_fd_sc_hd__or3_1 _5682_ (.A(_2541_),
    .B(_2543_),
    .C(_2544_),
    .X(_2546_));
 sky130_fd_sc_hd__a32o_1 _5683_ (.A1(net62),
    .A2(_2545_),
    .A3(_2546_),
    .B1(_2497_),
    .B2(_2540_),
    .X(_2547_));
 sky130_fd_sc_hd__a22o_1 _5684_ (.A1(net707),
    .A2(_2493_),
    .B1(_2547_),
    .B2(net59),
    .X(_0311_));
 sky130_fd_sc_hd__and2_1 _5685_ (.A(net611),
    .B(net76),
    .X(_2548_));
 sky130_fd_sc_hd__nor2_1 _5686_ (.A(\z80.tv80s.i_tv80_core.PC[14] ),
    .B(_2471_),
    .Y(_2549_));
 sky130_fd_sc_hd__or2_1 _5687_ (.A(_2548_),
    .B(_2549_),
    .X(_2550_));
 sky130_fd_sc_hd__o21a_1 _5688_ (.A1(_2543_),
    .A2(_2544_),
    .B1(_2542_),
    .X(_2551_));
 sky130_fd_sc_hd__nor2_1 _5689_ (.A(_2550_),
    .B(_2551_),
    .Y(_2552_));
 sky130_fd_sc_hd__and2_1 _5690_ (.A(_2550_),
    .B(_2551_),
    .X(_2553_));
 sky130_fd_sc_hd__or2_1 _5691_ (.A(_2552_),
    .B(_2553_),
    .X(_2554_));
 sky130_fd_sc_hd__mux2_1 _5692_ (.A0(\z80.tv80s.i_tv80_core.I[6] ),
    .A1(\z80.tv80s.i_tv80_core.PC[14] ),
    .S(net99),
    .X(_2555_));
 sky130_fd_sc_hd__a22o_1 _5693_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .A2(_1739_),
    .B1(net61),
    .B2(_2555_),
    .X(_2556_));
 sky130_fd_sc_hd__nand2_1 _5694_ (.A(net87),
    .B(_2556_),
    .Y(_2557_));
 sky130_fd_sc_hd__a21o_1 _5695_ (.A1(_1954_),
    .A2(_2557_),
    .B1(net68),
    .X(_2558_));
 sky130_fd_sc_hd__a32o_1 _5696_ (.A1(_1968_),
    .A2(_2497_),
    .A3(_2558_),
    .B1(_2554_),
    .B2(_2388_),
    .X(_2559_));
 sky130_fd_sc_hd__o2bb2a_1 _5697_ (.A1_N(_2377_),
    .A2_N(_2559_),
    .B1(_2492_),
    .B2(net611),
    .X(_0312_));
 sky130_fd_sc_hd__xnor2_1 _5698_ (.A(net667),
    .B(_2471_),
    .Y(_2560_));
 sky130_fd_sc_hd__o21ai_1 _5699_ (.A1(_2548_),
    .A2(_2552_),
    .B1(_2560_),
    .Y(_2561_));
 sky130_fd_sc_hd__o31a_1 _5700_ (.A1(_2548_),
    .A2(_2552_),
    .A3(_2560_),
    .B1(_2388_),
    .X(_2562_));
 sky130_fd_sc_hd__mux2_1 _5701_ (.A0(\z80.tv80s.i_tv80_core.I[7] ),
    .A1(\z80.tv80s.i_tv80_core.PC[15] ),
    .S(net99),
    .X(_2563_));
 sky130_fd_sc_hd__a22o_1 _5702_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[15] ),
    .A2(net64),
    .B1(net61),
    .B2(_2563_),
    .X(_2564_));
 sky130_fd_sc_hd__a21bo_1 _5703_ (.A1(net87),
    .A2(_2564_),
    .B1_N(_1970_),
    .X(_2565_));
 sky130_fd_sc_hd__mux2_1 _5704_ (.A0(_2565_),
    .A1(\z80.tv80s.di_reg[7] ),
    .S(net68),
    .X(_2566_));
 sky130_fd_sc_hd__mux2_1 _5705_ (.A0(_2566_),
    .A1(net667),
    .S(net55),
    .X(_2567_));
 sky130_fd_sc_hd__o2bb2a_1 _5706_ (.A1_N(_2561_),
    .A2_N(_2562_),
    .B1(_2567_),
    .B2(_2388_),
    .X(_2568_));
 sky130_fd_sc_hd__mux2_1 _5707_ (.A0(net667),
    .A1(_2568_),
    .S(_2377_),
    .X(_0313_));
 sky130_fd_sc_hd__or4b_1 _5708_ (.A(net679),
    .B(net542),
    .C(_0672_),
    .D_N(net635),
    .X(_2569_));
 sky130_fd_sc_hd__or2_4 _5709_ (.A(_1248_),
    .B(_2569_),
    .X(_2570_));
 sky130_fd_sc_hd__a21oi_1 _5710_ (.A1(net148),
    .A2(\z80.tv80s.i_tv80_core.ts[4] ),
    .B1(_0545_),
    .Y(_2571_));
 sky130_fd_sc_hd__or2_2 _5711_ (.A(_0698_),
    .B(_2571_),
    .X(_2572_));
 sky130_fd_sc_hd__a21o_2 _5712_ (.A1(_1237_),
    .A2(_2572_),
    .B1(net102),
    .X(_2573_));
 sky130_fd_sc_hd__inv_2 _5713_ (.A(_2573_),
    .Y(_2574_));
 sky130_fd_sc_hd__a21oi_4 _5714_ (.A1(_2570_),
    .A2(_2573_),
    .B1(net156),
    .Y(_2575_));
 sky130_fd_sc_hd__nand2_2 _5715_ (.A(net100),
    .B(_2570_),
    .Y(_2576_));
 sky130_fd_sc_hd__o22a_1 _5716_ (.A1(net88),
    .A2(_1468_),
    .B1(_1472_),
    .B2(net66),
    .X(_2577_));
 sky130_fd_sc_hd__o22a_1 _5717_ (.A1(_0803_),
    .A2(_2570_),
    .B1(_2576_),
    .B2(_2577_),
    .X(_2578_));
 sky130_fd_sc_hd__o22a_1 _5718_ (.A1(net795),
    .A2(_2575_),
    .B1(_2578_),
    .B2(net157),
    .X(_0314_));
 sky130_fd_sc_hd__o22a_1 _5719_ (.A1(net88),
    .A2(_1494_),
    .B1(_1499_),
    .B2(net66),
    .X(_2579_));
 sky130_fd_sc_hd__o22a_1 _5720_ (.A1(_0845_),
    .A2(_2570_),
    .B1(_2576_),
    .B2(_2579_),
    .X(_2580_));
 sky130_fd_sc_hd__o22a_1 _5721_ (.A1(net723),
    .A2(_2575_),
    .B1(_2580_),
    .B2(net157),
    .X(_0315_));
 sky130_fd_sc_hd__o22a_1 _5722_ (.A1(net88),
    .A2(_1507_),
    .B1(_1513_),
    .B2(net66),
    .X(_2581_));
 sky130_fd_sc_hd__o22a_1 _5723_ (.A1(_0922_),
    .A2(_2570_),
    .B1(_2576_),
    .B2(_2581_),
    .X(_2582_));
 sky130_fd_sc_hd__o22a_1 _5724_ (.A1(net687),
    .A2(_2575_),
    .B1(_2582_),
    .B2(net156),
    .X(_0316_));
 sky130_fd_sc_hd__o22a_1 _5725_ (.A1(net88),
    .A2(_1521_),
    .B1(_1527_),
    .B2(net66),
    .X(_2583_));
 sky130_fd_sc_hd__o22a_1 _5726_ (.A1(_0968_),
    .A2(_2570_),
    .B1(_2576_),
    .B2(_2583_),
    .X(_2584_));
 sky130_fd_sc_hd__o22a_1 _5727_ (.A1(net669),
    .A2(_2575_),
    .B1(_2584_),
    .B2(net156),
    .X(_0317_));
 sky130_fd_sc_hd__o22a_1 _5728_ (.A1(net88),
    .A2(_1536_),
    .B1(_1542_),
    .B2(net66),
    .X(_2585_));
 sky130_fd_sc_hd__o22a_1 _5729_ (.A1(_0999_),
    .A2(_2570_),
    .B1(_2576_),
    .B2(_2585_),
    .X(_2586_));
 sky130_fd_sc_hd__o22a_1 _5730_ (.A1(net780),
    .A2(_2575_),
    .B1(_2586_),
    .B2(net157),
    .X(_0318_));
 sky130_fd_sc_hd__o22a_1 _5731_ (.A1(net88),
    .A2(_1551_),
    .B1(_1557_),
    .B2(net66),
    .X(_2587_));
 sky130_fd_sc_hd__o22a_1 _5732_ (.A1(_1060_),
    .A2(_2570_),
    .B1(_2576_),
    .B2(_2587_),
    .X(_2588_));
 sky130_fd_sc_hd__o22a_1 _5733_ (.A1(net786),
    .A2(_2575_),
    .B1(_2588_),
    .B2(net157),
    .X(_0319_));
 sky130_fd_sc_hd__o22a_1 _5734_ (.A1(_1237_),
    .A2(_1566_),
    .B1(_1572_),
    .B2(net66),
    .X(_2589_));
 sky130_fd_sc_hd__o22a_1 _5735_ (.A1(_1092_),
    .A2(_2570_),
    .B1(_2576_),
    .B2(_2589_),
    .X(_2590_));
 sky130_fd_sc_hd__o22a_1 _5736_ (.A1(net767),
    .A2(_2575_),
    .B1(_2590_),
    .B2(net157),
    .X(_0320_));
 sky130_fd_sc_hd__o22a_1 _5737_ (.A1(_1237_),
    .A2(_1580_),
    .B1(_1586_),
    .B2(net66),
    .X(_2591_));
 sky130_fd_sc_hd__o22a_1 _5738_ (.A1(_1162_),
    .A2(_2570_),
    .B1(_2576_),
    .B2(_2591_),
    .X(_2592_));
 sky130_fd_sc_hd__o22a_1 _5739_ (.A1(net800),
    .A2(_2575_),
    .B1(_2592_),
    .B2(net157),
    .X(_0321_));
 sky130_fd_sc_hd__or2_4 _5740_ (.A(_0666_),
    .B(_2569_),
    .X(_2593_));
 sky130_fd_sc_hd__a21oi_4 _5741_ (.A1(_2573_),
    .A2(_2593_),
    .B1(net156),
    .Y(_2594_));
 sky130_fd_sc_hd__nand2_2 _5742_ (.A(net100),
    .B(_2593_),
    .Y(_2595_));
 sky130_fd_sc_hd__o22a_1 _5743_ (.A1(net88),
    .A2(_1593_),
    .B1(_1601_),
    .B2(net66),
    .X(_2596_));
 sky130_fd_sc_hd__o22a_1 _5744_ (.A1(_0803_),
    .A2(_2593_),
    .B1(_2595_),
    .B2(_2596_),
    .X(_2597_));
 sky130_fd_sc_hd__o22a_1 _5745_ (.A1(net703),
    .A2(_2594_),
    .B1(_2597_),
    .B2(net156),
    .X(_0322_));
 sky130_fd_sc_hd__o22a_1 _5746_ (.A1(net88),
    .A2(_1616_),
    .B1(_1622_),
    .B2(net66),
    .X(_2598_));
 sky130_fd_sc_hd__o22a_1 _5747_ (.A1(_0845_),
    .A2(_2593_),
    .B1(_2595_),
    .B2(_2598_),
    .X(_2599_));
 sky130_fd_sc_hd__o22a_1 _5748_ (.A1(net755),
    .A2(_2594_),
    .B1(_2599_),
    .B2(net156),
    .X(_0323_));
 sky130_fd_sc_hd__o22a_1 _5749_ (.A1(net88),
    .A2(_1629_),
    .B1(_1637_),
    .B2(net66),
    .X(_2600_));
 sky130_fd_sc_hd__o22a_1 _5750_ (.A1(_0922_),
    .A2(_2593_),
    .B1(_2595_),
    .B2(_2600_),
    .X(_2601_));
 sky130_fd_sc_hd__o22a_1 _5751_ (.A1(net774),
    .A2(_2594_),
    .B1(_2601_),
    .B2(net156),
    .X(_0324_));
 sky130_fd_sc_hd__o22a_1 _5752_ (.A1(net88),
    .A2(_1644_),
    .B1(_1650_),
    .B2(net66),
    .X(_2602_));
 sky130_fd_sc_hd__o22a_1 _5753_ (.A1(_0968_),
    .A2(_2593_),
    .B1(_2595_),
    .B2(_2602_),
    .X(_2603_));
 sky130_fd_sc_hd__o22a_1 _5754_ (.A1(net788),
    .A2(_2594_),
    .B1(_2603_),
    .B2(net156),
    .X(_0325_));
 sky130_fd_sc_hd__o22a_1 _5755_ (.A1(net88),
    .A2(_1657_),
    .B1(_1664_),
    .B2(net66),
    .X(_2604_));
 sky130_fd_sc_hd__o22a_1 _5756_ (.A1(_0999_),
    .A2(_2593_),
    .B1(_2595_),
    .B2(_2604_),
    .X(_2605_));
 sky130_fd_sc_hd__o22a_1 _5757_ (.A1(net782),
    .A2(_2594_),
    .B1(_2605_),
    .B2(net156),
    .X(_0326_));
 sky130_fd_sc_hd__o22a_1 _5758_ (.A1(net88),
    .A2(_1671_),
    .B1(_1677_),
    .B2(net66),
    .X(_2606_));
 sky130_fd_sc_hd__o22a_1 _5759_ (.A1(_1060_),
    .A2(_2593_),
    .B1(_2595_),
    .B2(_2606_),
    .X(_2607_));
 sky130_fd_sc_hd__o22a_1 _5760_ (.A1(net681),
    .A2(_2594_),
    .B1(_2607_),
    .B2(net156),
    .X(_0327_));
 sky130_fd_sc_hd__nand2b_1 _5761_ (.A_N(net473),
    .B(net66),
    .Y(_2608_));
 sky130_fd_sc_hd__or3_1 _5762_ (.A(net102),
    .B(_1690_),
    .C(net66),
    .X(_2609_));
 sky130_fd_sc_hd__a21bo_1 _5763_ (.A1(_2608_),
    .A2(_2609_),
    .B1_N(net88),
    .X(_2610_));
 sky130_fd_sc_hd__or2_1 _5764_ (.A(net473),
    .B(net100),
    .X(_2611_));
 sky130_fd_sc_hd__o311a_1 _5765_ (.A1(net102),
    .A2(net88),
    .A3(_1682_),
    .B1(_2593_),
    .C1(_2611_),
    .X(_2612_));
 sky130_fd_sc_hd__o2bb2a_1 _5766_ (.A1_N(_2612_),
    .A2_N(_2610_),
    .B1(_2593_),
    .B2(_1091_),
    .X(_2613_));
 sky130_fd_sc_hd__nand2_1 _5767_ (.A(net156),
    .B(net473),
    .Y(_2614_));
 sky130_fd_sc_hd__o21ai_1 _5768_ (.A1(net156),
    .A2(_2613_),
    .B1(net474),
    .Y(_0328_));
 sky130_fd_sc_hd__o32a_1 _5769_ (.A1(_1700_),
    .A2(_1701_),
    .A3(_2572_),
    .B1(_1697_),
    .B2(net88),
    .X(_2615_));
 sky130_fd_sc_hd__o22a_1 _5770_ (.A1(net771),
    .A2(_2574_),
    .B1(_2615_),
    .B2(net102),
    .X(_2616_));
 sky130_fd_sc_hd__mux2_1 _5771_ (.A0(_1162_),
    .A1(_2616_),
    .S(_2593_),
    .X(_2617_));
 sky130_fd_sc_hd__mux2_1 _5772_ (.A0(net771),
    .A1(_2617_),
    .S(net114),
    .X(_0329_));
 sky130_fd_sc_hd__or2_4 _5773_ (.A(net158),
    .B(_2234_),
    .X(_2618_));
 sky130_fd_sc_hd__mux2_1 _5774_ (.A0(\z80.tv80s.i_tv80_core.ACC[0] ),
    .A1(net658),
    .S(_2618_),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _5775_ (.A0(\z80.tv80s.i_tv80_core.ACC[1] ),
    .A1(net709),
    .S(_2618_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _5776_ (.A0(\z80.tv80s.i_tv80_core.ACC[2] ),
    .A1(net654),
    .S(_2618_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _5777_ (.A0(\z80.tv80s.i_tv80_core.ACC[3] ),
    .A1(net705),
    .S(_2618_),
    .X(_0333_));
 sky130_fd_sc_hd__mux2_1 _5778_ (.A0(\z80.tv80s.i_tv80_core.ACC[4] ),
    .A1(net665),
    .S(_2618_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _5779_ (.A0(\z80.tv80s.i_tv80_core.ACC[5] ),
    .A1(net693),
    .S(_2618_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _5780_ (.A0(\z80.tv80s.i_tv80_core.ACC[6] ),
    .A1(net689),
    .S(_2618_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _5781_ (.A0(\z80.tv80s.i_tv80_core.ACC[7] ),
    .A1(net685),
    .S(_2618_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _5782_ (.A0(\z80.tv80s.i_tv80_core.F[0] ),
    .A1(net673),
    .S(_2618_),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _5783_ (.A0(\z80.tv80s.i_tv80_core.F[1] ),
    .A1(net695),
    .S(_2618_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _5784_ (.A0(\z80.tv80s.i_tv80_core.F[2] ),
    .A1(net646),
    .S(_2618_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _5785_ (.A0(net621),
    .A1(\z80.tv80s.i_tv80_core.Fp[3] ),
    .S(_2618_),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _5786_ (.A0(\z80.tv80s.i_tv80_core.F[4] ),
    .A1(net731),
    .S(_2618_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _5787_ (.A0(\z80.tv80s.i_tv80_core.F[5] ),
    .A1(net660),
    .S(_2618_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _5788_ (.A0(\z80.tv80s.i_tv80_core.F[6] ),
    .A1(net650),
    .S(_2618_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _5789_ (.A0(\z80.tv80s.i_tv80_core.F[7] ),
    .A1(net691),
    .S(_2618_),
    .X(_0345_));
 sky130_fd_sc_hd__and4b_4 _5790_ (.A_N(net635),
    .B(_0673_),
    .C(net679),
    .D(net542),
    .X(_2619_));
 sky130_fd_sc_hd__o21a_2 _5791_ (.A1(net102),
    .A2(_2243_),
    .B1(_2234_),
    .X(_2620_));
 sky130_fd_sc_hd__a2bb2o_1 _5792_ (.A1_N(\z80.tv80s.i_tv80_core.ACC[0] ),
    .A2_N(_2243_),
    .B1(_2232_),
    .B2(net658),
    .X(_2621_));
 sky130_fd_sc_hd__a22o_1 _5793_ (.A1(\z80.tv80s.i_tv80_core.ACC[0] ),
    .A2(_2620_),
    .B1(_2621_),
    .B2(net100),
    .X(_2622_));
 sky130_fd_sc_hd__nor2_2 _5794_ (.A(net129),
    .B(_2249_),
    .Y(_2623_));
 sky130_fd_sc_hd__a22o_1 _5795_ (.A1(_2249_),
    .A2(_2622_),
    .B1(_2623_),
    .B2(net588),
    .X(_2624_));
 sky130_fd_sc_hd__mux2_1 _5796_ (.A0(_2624_),
    .A1(_0803_),
    .S(_2619_),
    .X(_2625_));
 sky130_fd_sc_hd__mux2_1 _5797_ (.A0(net815),
    .A1(_2625_),
    .S(net113),
    .X(_0346_));
 sky130_fd_sc_hd__a2bb2o_1 _5798_ (.A1_N(\z80.tv80s.i_tv80_core.ACC[1] ),
    .A2_N(_2243_),
    .B1(_2232_),
    .B2(net709),
    .X(_2626_));
 sky130_fd_sc_hd__a22o_1 _5799_ (.A1(\z80.tv80s.i_tv80_core.ACC[1] ),
    .A2(_2620_),
    .B1(_2626_),
    .B2(net100),
    .X(_2627_));
 sky130_fd_sc_hd__a22o_1 _5800_ (.A1(net629),
    .A2(_2623_),
    .B1(_2627_),
    .B2(_2249_),
    .X(_2628_));
 sky130_fd_sc_hd__mux2_1 _5801_ (.A0(_2628_),
    .A1(_0845_),
    .S(_2619_),
    .X(_2629_));
 sky130_fd_sc_hd__mux2_1 _5802_ (.A0(net820),
    .A1(_2629_),
    .S(net113),
    .X(_0347_));
 sky130_fd_sc_hd__a2bb2o_1 _5803_ (.A1_N(\z80.tv80s.i_tv80_core.ACC[2] ),
    .A2_N(_2243_),
    .B1(_2232_),
    .B2(net654),
    .X(_2630_));
 sky130_fd_sc_hd__a22o_1 _5804_ (.A1(\z80.tv80s.i_tv80_core.ACC[2] ),
    .A2(_2620_),
    .B1(_2630_),
    .B2(net100),
    .X(_2631_));
 sky130_fd_sc_hd__a22o_1 _5805_ (.A1(net566),
    .A2(_2623_),
    .B1(_2631_),
    .B2(_2249_),
    .X(_2632_));
 sky130_fd_sc_hd__mux2_1 _5806_ (.A0(_2632_),
    .A1(_0922_),
    .S(_2619_),
    .X(_2633_));
 sky130_fd_sc_hd__mux2_1 _5807_ (.A0(net810),
    .A1(_2633_),
    .S(net113),
    .X(_0348_));
 sky130_fd_sc_hd__a22o_1 _5808_ (.A1(net705),
    .A2(_2232_),
    .B1(_2244_),
    .B2(_2738_),
    .X(_2634_));
 sky130_fd_sc_hd__a22o_1 _5809_ (.A1(\z80.tv80s.i_tv80_core.ACC[3] ),
    .A2(_2620_),
    .B1(_2634_),
    .B2(net100),
    .X(_2635_));
 sky130_fd_sc_hd__a22o_1 _5810_ (.A1(net615),
    .A2(_2623_),
    .B1(_2635_),
    .B2(_2249_),
    .X(_2636_));
 sky130_fd_sc_hd__mux2_1 _5811_ (.A0(_2636_),
    .A1(_0968_),
    .S(_2619_),
    .X(_2637_));
 sky130_fd_sc_hd__mux2_1 _5812_ (.A0(net816),
    .A1(_2637_),
    .S(net113),
    .X(_0349_));
 sky130_fd_sc_hd__a2bb2o_1 _5813_ (.A1_N(\z80.tv80s.i_tv80_core.ACC[4] ),
    .A2_N(_2243_),
    .B1(_2232_),
    .B2(net665),
    .X(_2638_));
 sky130_fd_sc_hd__a22o_1 _5814_ (.A1(net811),
    .A2(_2620_),
    .B1(_2638_),
    .B2(net100),
    .X(_2639_));
 sky130_fd_sc_hd__a22o_1 _5815_ (.A1(net644),
    .A2(_2623_),
    .B1(_2639_),
    .B2(_2249_),
    .X(_2640_));
 sky130_fd_sc_hd__mux2_1 _5816_ (.A0(_2640_),
    .A1(_0999_),
    .S(_2619_),
    .X(_2641_));
 sky130_fd_sc_hd__mux2_1 _5817_ (.A0(net811),
    .A1(_2641_),
    .S(net113),
    .X(_0350_));
 sky130_fd_sc_hd__a22o_1 _5818_ (.A1(net693),
    .A2(_2232_),
    .B1(_2244_),
    .B2(_2739_),
    .X(_2642_));
 sky130_fd_sc_hd__a22o_1 _5819_ (.A1(\z80.tv80s.i_tv80_core.ACC[5] ),
    .A2(_2620_),
    .B1(_2642_),
    .B2(net100),
    .X(_2643_));
 sky130_fd_sc_hd__a22o_1 _5820_ (.A1(net597),
    .A2(_2623_),
    .B1(_2643_),
    .B2(_2249_),
    .X(_2644_));
 sky130_fd_sc_hd__mux2_1 _5821_ (.A0(_2644_),
    .A1(_1060_),
    .S(_2619_),
    .X(_2645_));
 sky130_fd_sc_hd__mux2_1 _5822_ (.A0(net813),
    .A1(_2645_),
    .S(net113),
    .X(_0351_));
 sky130_fd_sc_hd__a2bb2o_1 _5823_ (.A1_N(\z80.tv80s.i_tv80_core.ACC[6] ),
    .A2_N(_2243_),
    .B1(_2232_),
    .B2(net689),
    .X(_2646_));
 sky130_fd_sc_hd__a22o_1 _5824_ (.A1(\z80.tv80s.i_tv80_core.ACC[6] ),
    .A2(_2620_),
    .B1(_2646_),
    .B2(net100),
    .X(_2647_));
 sky130_fd_sc_hd__a22o_1 _5825_ (.A1(net549),
    .A2(_2623_),
    .B1(_2647_),
    .B2(_2249_),
    .X(_2648_));
 sky130_fd_sc_hd__mux2_1 _5826_ (.A0(_2648_),
    .A1(_1092_),
    .S(_2619_),
    .X(_2649_));
 sky130_fd_sc_hd__mux2_1 _5827_ (.A0(net812),
    .A1(_2649_),
    .S(net113),
    .X(_0352_));
 sky130_fd_sc_hd__a2bb2o_1 _5828_ (.A1_N(\z80.tv80s.i_tv80_core.ACC[7] ),
    .A2_N(_2243_),
    .B1(_2232_),
    .B2(net685),
    .X(_2650_));
 sky130_fd_sc_hd__a22o_1 _5829_ (.A1(net808),
    .A2(_2620_),
    .B1(_2650_),
    .B2(net101),
    .X(_2651_));
 sky130_fd_sc_hd__a22o_1 _5830_ (.A1(net578),
    .A2(_2623_),
    .B1(_2651_),
    .B2(_2249_),
    .X(_2652_));
 sky130_fd_sc_hd__mux2_1 _5831_ (.A0(_2652_),
    .A1(_1162_),
    .S(_2619_),
    .X(_2653_));
 sky130_fd_sc_hd__mux2_1 _5832_ (.A0(net808),
    .A1(_2653_),
    .S(net113),
    .X(_0353_));
 sky130_fd_sc_hd__nor4_1 _5833_ (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ),
    .B(_0667_),
    .C(_0672_),
    .D(_1248_),
    .Y(_2654_));
 sky130_fd_sc_hd__or4_4 _5834_ (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ),
    .B(_0667_),
    .C(_0672_),
    .D(_1248_),
    .X(_2655_));
 sky130_fd_sc_hd__a21oi_4 _5835_ (.A1(_0671_),
    .A2(_2655_),
    .B1(net158),
    .Y(_2656_));
 sky130_fd_sc_hd__inv_2 _5836_ (.A(_2656_),
    .Y(_2657_));
 sky130_fd_sc_hd__or2_2 _5837_ (.A(_0671_),
    .B(_2654_),
    .X(_2658_));
 sky130_fd_sc_hd__and3_4 _5838_ (.A(_0377_),
    .B(_0379_),
    .C(_0472_),
    .X(_2659_));
 sky130_fd_sc_hd__a21o_1 _5839_ (.A1(net119),
    .A2(\z80.tv80s.i_tv80_core.BusB[4] ),
    .B1(_1154_),
    .X(_2660_));
 sky130_fd_sc_hd__mux2_1 _5840_ (.A0(\z80.tv80s.i_tv80_core.BusB[0] ),
    .A1(_2660_),
    .S(_2659_),
    .X(_2661_));
 sky130_fd_sc_hd__o22a_1 _5841_ (.A1(_0803_),
    .A2(_2655_),
    .B1(_2658_),
    .B2(_2661_),
    .X(_2662_));
 sky130_fd_sc_hd__o22a_1 _5842_ (.A1(net553),
    .A2(_2656_),
    .B1(_2662_),
    .B2(net158),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _5843_ (.A0(\z80.tv80s.i_tv80_core.BusB[5] ),
    .A1(\z80.tv80s.i_tv80_core.BusA[1] ),
    .S(net129),
    .X(_2663_));
 sky130_fd_sc_hd__mux2_1 _5844_ (.A0(\z80.tv80s.i_tv80_core.BusB[1] ),
    .A1(_2663_),
    .S(_2659_),
    .X(_2664_));
 sky130_fd_sc_hd__inv_2 _5845_ (.A(_2664_),
    .Y(_2665_));
 sky130_fd_sc_hd__o2bb2a_1 _5846_ (.A1_N(_0845_),
    .A2_N(_2654_),
    .B1(_2658_),
    .B2(_2665_),
    .X(_2666_));
 sky130_fd_sc_hd__a2bb2o_1 _5847_ (.A1_N(net158),
    .A2_N(_2666_),
    .B1(_2657_),
    .B2(net532),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _5848_ (.A0(\z80.tv80s.i_tv80_core.BusB[6] ),
    .A1(\z80.tv80s.i_tv80_core.BusA[2] ),
    .S(net129),
    .X(_2667_));
 sky130_fd_sc_hd__mux2_1 _5849_ (.A0(\z80.tv80s.i_tv80_core.BusB[2] ),
    .A1(_2667_),
    .S(_2659_),
    .X(_2668_));
 sky130_fd_sc_hd__o22a_1 _5850_ (.A1(_0922_),
    .A2(_2655_),
    .B1(_2658_),
    .B2(_2668_),
    .X(_2669_));
 sky130_fd_sc_hd__o22a_1 _5851_ (.A1(net534),
    .A2(_2656_),
    .B1(_2669_),
    .B2(net158),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _5852_ (.A0(\z80.tv80s.i_tv80_core.BusB[7] ),
    .A1(\z80.tv80s.i_tv80_core.BusA[3] ),
    .S(net129),
    .X(_2670_));
 sky130_fd_sc_hd__mux2_1 _5853_ (.A0(\z80.tv80s.i_tv80_core.BusB[3] ),
    .A1(_2670_),
    .S(_2659_),
    .X(_2671_));
 sky130_fd_sc_hd__o22a_1 _5854_ (.A1(_0968_),
    .A2(_2655_),
    .B1(_2658_),
    .B2(_2671_),
    .X(_2672_));
 sky130_fd_sc_hd__o22a_1 _5855_ (.A1(net572),
    .A2(_2656_),
    .B1(_2672_),
    .B2(net158),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _5856_ (.A0(\z80.tv80s.i_tv80_core.BusA[0] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[0] ),
    .S(net129),
    .X(_2673_));
 sky130_fd_sc_hd__mux2_1 _5857_ (.A0(\z80.tv80s.i_tv80_core.BusB[4] ),
    .A1(_2673_),
    .S(_2659_),
    .X(_2674_));
 sky130_fd_sc_hd__o22a_1 _5858_ (.A1(_0999_),
    .A2(_2655_),
    .B1(_2658_),
    .B2(_2674_),
    .X(_2675_));
 sky130_fd_sc_hd__o22a_1 _5859_ (.A1(net551),
    .A2(_2656_),
    .B1(_2675_),
    .B2(net159),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _5860_ (.A0(\z80.tv80s.i_tv80_core.BusA[1] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[1] ),
    .S(net129),
    .X(_2676_));
 sky130_fd_sc_hd__mux2_1 _5861_ (.A0(\z80.tv80s.i_tv80_core.BusB[5] ),
    .A1(_2676_),
    .S(_2659_),
    .X(_2677_));
 sky130_fd_sc_hd__o22a_1 _5862_ (.A1(_1060_),
    .A2(_2655_),
    .B1(_2658_),
    .B2(_2677_),
    .X(_2678_));
 sky130_fd_sc_hd__o22a_1 _5863_ (.A1(net540),
    .A2(_2656_),
    .B1(_2678_),
    .B2(net159),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _5864_ (.A0(\z80.tv80s.i_tv80_core.BusA[2] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[2] ),
    .S(net129),
    .X(_2679_));
 sky130_fd_sc_hd__mux2_1 _5865_ (.A0(\z80.tv80s.i_tv80_core.BusB[6] ),
    .A1(_2679_),
    .S(_2659_),
    .X(_2680_));
 sky130_fd_sc_hd__o22a_1 _5866_ (.A1(_1092_),
    .A2(_2655_),
    .B1(_2658_),
    .B2(_2680_),
    .X(_2681_));
 sky130_fd_sc_hd__o22a_1 _5867_ (.A1(net592),
    .A2(_2656_),
    .B1(_2681_),
    .B2(net159),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _5868_ (.A0(\z80.tv80s.i_tv80_core.BusA[3] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[3] ),
    .S(net129),
    .X(_2682_));
 sky130_fd_sc_hd__mux2_1 _5869_ (.A0(\z80.tv80s.i_tv80_core.BusB[7] ),
    .A1(_2682_),
    .S(_2659_),
    .X(_2683_));
 sky130_fd_sc_hd__o22a_1 _5870_ (.A1(_1162_),
    .A2(_2655_),
    .B1(_2658_),
    .B2(_2683_),
    .X(_2684_));
 sky130_fd_sc_hd__o22a_1 _5871_ (.A1(net603),
    .A2(_2656_),
    .B1(_2684_),
    .B2(net158),
    .X(_0361_));
 sky130_fd_sc_hd__nand2_2 _5872_ (.A(net103),
    .B(_1476_),
    .Y(_2685_));
 sky130_fd_sc_hd__and2_1 _5873_ (.A(net1),
    .B(_2685_),
    .X(_2686_));
 sky130_fd_sc_hd__a21o_1 _5874_ (.A1(net869),
    .A2(net163),
    .B1(net103),
    .X(_2687_));
 sky130_fd_sc_hd__and3_4 _5875_ (.A(net110),
    .B(_0545_),
    .C(_2687_),
    .X(_2688_));
 sky130_fd_sc_hd__o21ai_4 _5876_ (.A1(net101),
    .A2(_1477_),
    .B1(_2688_),
    .Y(_2689_));
 sky130_fd_sc_hd__o22a_1 _5877_ (.A1(net570),
    .A2(_2688_),
    .B1(_2689_),
    .B2(_2686_),
    .X(_0362_));
 sky130_fd_sc_hd__and2_1 _5878_ (.A(net2),
    .B(_2685_),
    .X(_2690_));
 sky130_fd_sc_hd__o22a_1 _5879_ (.A1(net134),
    .A2(_2688_),
    .B1(_2689_),
    .B2(_2690_),
    .X(_0363_));
 sky130_fd_sc_hd__and2_1 _5880_ (.A(net3),
    .B(_2685_),
    .X(_2691_));
 sky130_fd_sc_hd__o22a_1 _5881_ (.A1(net132),
    .A2(_2688_),
    .B1(_2689_),
    .B2(_2691_),
    .X(_0364_));
 sky130_fd_sc_hd__and2_1 _5882_ (.A(net4),
    .B(_2685_),
    .X(_2692_));
 sky130_fd_sc_hd__o22a_1 _5883_ (.A1(net130),
    .A2(_2688_),
    .B1(_2689_),
    .B2(_2692_),
    .X(_0365_));
 sky130_fd_sc_hd__and2_1 _5884_ (.A(net5),
    .B(_2685_),
    .X(_2693_));
 sky130_fd_sc_hd__o22a_1 _5885_ (.A1(net123),
    .A2(_2688_),
    .B1(_2689_),
    .B2(_2693_),
    .X(_0366_));
 sky130_fd_sc_hd__and2_1 _5886_ (.A(net6),
    .B(_2685_),
    .X(_2694_));
 sky130_fd_sc_hd__o22a_1 _5887_ (.A1(net120),
    .A2(_2688_),
    .B1(_2689_),
    .B2(_2694_),
    .X(_0367_));
 sky130_fd_sc_hd__and2_1 _5888_ (.A(net7),
    .B(_2685_),
    .X(_2695_));
 sky130_fd_sc_hd__o22a_1 _5889_ (.A1(net850),
    .A2(_2688_),
    .B1(_2689_),
    .B2(_2695_),
    .X(_0368_));
 sky130_fd_sc_hd__and2_1 _5890_ (.A(net8),
    .B(_2685_),
    .X(_2696_));
 sky130_fd_sc_hd__o22a_1 _5891_ (.A1(net838),
    .A2(_2688_),
    .B1(_2689_),
    .B2(_2696_),
    .X(_0369_));
 sky130_fd_sc_hd__dfxtp_1 _5892_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net334),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5893_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0037_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5894_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0038_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5895_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net440),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5896_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net373),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5897_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0041_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5898_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net489),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5899_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net336),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5900_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net453),
    .RESET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.mcycles[1] ));
 sky130_fd_sc_hd__dfrtp_1 _5901_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net596),
    .RESET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.mcycles[2] ));
 sky130_fd_sc_hd__dfrtp_1 _5902_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net421),
    .RESET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.mcycles[4] ));
 sky130_fd_sc_hd__dfrtp_1 _5903_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net344),
    .RESET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.mcycles[5] ));
 sky130_fd_sc_hd__dfxtp_1 _5904_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(net245),
    .Q(\z80.tv80s.i_tv80_core.RegAddrA_r[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5905_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(net585),
    .Q(\z80.tv80s.i_tv80_core.RegAddrB_r[2] ));
 sky130_fd_sc_hd__dfxtp_1 _5906_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net304),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5907_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0047_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5908_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net312),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5909_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net381),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5910_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net338),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5911_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net316),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5912_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0052_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5913_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net276),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5914_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0054_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrC[2] ));
 sky130_fd_sc_hd__dfrtp_1 _5915_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net544),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.PreserveC_r ));
 sky130_fd_sc_hd__dfstp_1 _5916_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(net799),
    .SET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.ISet[0] ));
 sky130_fd_sc_hd__dfrtp_1 _5917_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net587),
    .RESET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.ISet[1] ));
 sky130_fd_sc_hd__dfrtp_4 _5918_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_0002_),
    .RESET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.ISet[2] ));
 sky130_fd_sc_hd__dfrtp_1 _5919_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net310),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.ISet[3] ));
 sky130_fd_sc_hd__dfxtp_1 _5920_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net395),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5921_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net427),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5922_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net361),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5923_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net342),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5924_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net359),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5925_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net355),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5926_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net375),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5927_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net429),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5928_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0064_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5929_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net296),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5930_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net272),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5931_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net377),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5932_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net286),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5933_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net393),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5934_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net298),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5935_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net371),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][7] ));
 sky130_fd_sc_hd__dfxtp_2 _5936_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0072_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrC[1] ));
 sky130_fd_sc_hd__dfxtp_1 _5937_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net387),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5938_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net280),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5939_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net284),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5940_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net300),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5941_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net288),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5942_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net290),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5943_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net282),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5944_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net328),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5945_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0081_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5946_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0082_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5947_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0083_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5948_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net493),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5949_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0085_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5950_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net384),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5951_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0087_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5952_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net496),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][7] ));
 sky130_fd_sc_hd__dfstp_1 _5953_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_0020_),
    .SET_B(net173),
    .Q(net50));
 sky130_fd_sc_hd__dfstp_1 _5954_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_0018_),
    .SET_B(net173),
    .Q(net47));
 sky130_fd_sc_hd__dfstp_1 _5955_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_0017_),
    .SET_B(net173),
    .Q(net48));
 sky130_fd_sc_hd__dfstp_1 _5956_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net806),
    .SET_B(net173),
    .Q(net49));
 sky130_fd_sc_hd__dfxtp_1 _5957_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net514),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5958_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net539),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5959_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0091_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5960_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net357),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5961_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0093_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5962_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net405),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5963_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net438),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5964_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0096_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5965_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net363),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5966_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0098_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5967_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net318),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5968_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net466),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5969_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0101_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5970_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0102_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5971_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0103_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5972_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net468),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][7] ));
 sky130_fd_sc_hd__dfrtp_1 _5973_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net258),
    .RESET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[1] ));
 sky130_fd_sc_hd__dfrtp_1 _5974_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net260),
    .RESET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[2] ));
 sky130_fd_sc_hd__dfrtp_1 _5975_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net274),
    .RESET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[3] ));
 sky130_fd_sc_hd__dfrtp_1 _5976_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net262),
    .RESET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[4] ));
 sky130_fd_sc_hd__dfrtp_1 _5977_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net462),
    .RESET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[5] ));
 sky130_fd_sc_hd__dfrtp_1 _5978_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(_0011_),
    .RESET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[6] ));
 sky130_fd_sc_hd__dfrtp_1 _5979_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net491),
    .RESET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[7] ));
 sky130_fd_sc_hd__dfxtp_1 _5980_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net435),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5981_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(net367),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5982_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net346),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5983_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0108_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5984_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0109_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5985_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net322),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5986_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net379),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5987_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net324),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5988_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net407),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5989_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0114_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5990_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net306),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5991_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net415),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _5992_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net314),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _5993_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net365),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _5994_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net478),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _5995_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0120_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _5996_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net510),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _5997_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net523),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _5998_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0123_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _5999_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net412),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6000_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0125_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6001_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net320),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6002_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net332),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6003_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0128_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6004_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net348),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6005_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0130_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6006_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0131_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6007_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net326),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6008_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net417),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6009_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net353),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6010_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0135_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6011_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0136_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6012_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0137_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6013_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0138_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6014_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0139_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6015_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0140_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6016_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0141_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6017_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net448),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6018_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net464),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6019_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net512),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6020_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net369),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6021_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net419),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6022_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0147_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6023_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0148_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6024_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net389),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6025_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net446),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6026_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net351),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6027_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net432),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6028_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net340),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6029_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0154_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6030_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0155_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6031_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net391),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6032_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net424),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6033_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net401),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6034_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net443),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6035_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net460),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][7] ));
 sky130_fd_sc_hd__dfrtp_1 _6036_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net518),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.IStatus[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6037_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net264),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.IStatus[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6038_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net837),
    .RESET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__dfrtp_1 _6039_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(net270),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.BTR_r ));
 sky130_fd_sc_hd__dfrtp_1 _6040_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0163_),
    .RESET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6041_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net680),
    .RESET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6042_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0165_),
    .RESET_B(net183),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6043_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0166_),
    .RESET_B(net183),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6044_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0167_),
    .RESET_B(net183),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6045_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net410),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.Z16_r ));
 sky130_fd_sc_hd__dfrtp_4 _6046_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net712),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.Arith16_r ));
 sky130_fd_sc_hd__dfrtp_4 _6047_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0023_),
    .RESET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.BusReq_s ));
 sky130_fd_sc_hd__dfrtp_4 _6048_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(net505),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.NMICycle ));
 sky130_fd_sc_hd__dfrtp_1 _6049_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(net750),
    .RESET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.BusAck ));
 sky130_fd_sc_hd__dfrtp_4 _6050_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(net747),
    .RESET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.IntCycle ));
 sky130_fd_sc_hd__dfrtp_1 _6051_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(net508),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.XY_State[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6052_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net577),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.XY_State[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6053_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0175_),
    .RESET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.Alternate ));
 sky130_fd_sc_hd__dfrtp_4 _6054_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net745),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6055_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net766),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6056_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net760),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6057_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(net758),
    .RESET_B(net183),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6058_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(net764),
    .RESET_B(net183),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6059_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(net777),
    .RESET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6060_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(net770),
    .RESET_B(net183),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6061_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net752),
    .RESET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sky130_fd_sc_hd__dfrtp_2 _6062_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net608),
    .RESET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[8] ));
 sky130_fd_sc_hd__dfrtp_2 _6063_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net672),
    .RESET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[9] ));
 sky130_fd_sc_hd__dfrtp_4 _6064_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net738),
    .RESET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[10] ));
 sky130_fd_sc_hd__dfrtp_2 _6065_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net698),
    .RESET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[11] ));
 sky130_fd_sc_hd__dfrtp_4 _6066_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net719),
    .RESET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[12] ));
 sky130_fd_sc_hd__dfrtp_4 _6067_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net728),
    .RESET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[13] ));
 sky130_fd_sc_hd__dfrtp_2 _6068_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net641),
    .RESET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[14] ));
 sky130_fd_sc_hd__dfrtp_2 _6069_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net676),
    .RESET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[15] ));
 sky130_fd_sc_hd__dfrtp_4 _6070_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net825),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6071_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net827),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.ALU_Op_r[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6072_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_0194_),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6073_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net832),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6074_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_0196_),
    .RESET_B(net175),
    .Q(\z80.tv80s.i_tv80_core.Save_ALU_r ));
 sky130_fd_sc_hd__dfrtp_1 _6075_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net268),
    .RESET_B(net170),
    .Q(_0033_));
 sky130_fd_sc_hd__dfrtp_1 _6076_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net252),
    .RESET_B(net170),
    .Q(_0034_));
 sky130_fd_sc_hd__dfrtp_1 _6077_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0031_),
    .RESET_B(net170),
    .Q(_0035_));
 sky130_fd_sc_hd__dfrtp_1 _6078_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net600),
    .RESET_B(net174),
    .Q(net51));
 sky130_fd_sc_hd__dfrtp_1 _6079_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net559),
    .RESET_B(net174),
    .Q(net52));
 sky130_fd_sc_hd__dfrtp_1 _6080_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net527),
    .RESET_B(net174),
    .Q(net23));
 sky130_fd_sc_hd__dfrtp_1 _6081_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net569),
    .RESET_B(net174),
    .Q(net24));
 sky130_fd_sc_hd__dfrtp_1 _6082_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net546),
    .RESET_B(net174),
    .Q(net25));
 sky130_fd_sc_hd__dfrtp_1 _6083_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net565),
    .RESET_B(net174),
    .Q(net26));
 sky130_fd_sc_hd__dfrtp_1 _6084_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net548),
    .RESET_B(net175),
    .Q(net27));
 sky130_fd_sc_hd__dfrtp_1 _6085_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net531),
    .RESET_B(net175),
    .Q(net28));
 sky130_fd_sc_hd__dfrtp_1 _6086_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net529),
    .RESET_B(net175),
    .Q(net29));
 sky130_fd_sc_hd__dfrtp_2 _6087_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net575),
    .RESET_B(net181),
    .Q(net30));
 sky130_fd_sc_hd__dfrtp_2 _6088_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net614),
    .RESET_B(net182),
    .Q(net31));
 sky130_fd_sc_hd__dfrtp_2 _6089_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net561),
    .RESET_B(net181),
    .Q(net32));
 sky130_fd_sc_hd__dfrtp_2 _6090_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net583),
    .RESET_B(net182),
    .Q(net34));
 sky130_fd_sc_hd__dfrtp_2 _6091_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net557),
    .RESET_B(net181),
    .Q(net35));
 sky130_fd_sc_hd__dfrtp_2 _6092_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net563),
    .RESET_B(net182),
    .Q(net36));
 sky130_fd_sc_hd__dfrtp_2 _6093_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net537),
    .RESET_B(net182),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_1 _6094_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net486),
    .Q(\z80.tv80s.i_tv80_core.IncDecZ ));
 sky130_fd_sc_hd__dfrtp_1 _6095_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(net792),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.No_BTR ));
 sky130_fd_sc_hd__dfxtp_1 _6096_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0214_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6097_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net229),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6098_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net225),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6099_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net237),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6100_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net231),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6101_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net235),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6102_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net219),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6103_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net221),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6104_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net239),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6105_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net254),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6106_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net233),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6107_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net227),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6108_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net247),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6109_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net249),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6110_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net223),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6111_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net243),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[15] ));
 sky130_fd_sc_hd__dfxtp_2 _6112_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0230_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrC[0] ));
 sky130_fd_sc_hd__dfxtp_4 _6113_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net581),
    .Q(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6114_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net702),
    .Q(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6115_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net653),
    .Q(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__dfxtp_2 _6116_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net628),
    .Q(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6117_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net591),
    .Q(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__dfxtp_4 _6118_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net606),
    .Q(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__dfxtp_2 _6119_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net602),
    .Q(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__dfxtp_4 _6120_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net626),
    .Q(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__dfrtp_2 _6121_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0025_),
    .RESET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.INT_s ));
 sky130_fd_sc_hd__dfrtp_1 _6122_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net516),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.Auto_Wait_t1 ));
 sky130_fd_sc_hd__dfrtp_1 _6123_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_0022_),
    .RESET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.Auto_Wait_t2 ));
 sky130_fd_sc_hd__dfstp_1 _6124_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0239_),
    .SET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6125_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net863),
    .RESET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6126_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net861),
    .RESET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6127_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net822),
    .RESET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6128_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net715),
    .RESET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6129_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net736),
    .RESET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6130_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net804),
    .RESET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6131_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0246_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6132_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net525),
    .Q(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6133_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net520),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.NMI_s ));
 sky130_fd_sc_hd__dfrtp_1 _6134_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net10),
    .RESET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.Oldnmi_n ));
 sky130_fd_sc_hd__dfxtp_4 _6135_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net726),
    .Q(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__dfxtp_4 _6136_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net740),
    .Q(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__dfxtp_4 _6137_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net637),
    .Q(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__dfxtp_4 _6138_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net618),
    .Q(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__dfxtp_4 _6139_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net634),
    .Q(\z80.tv80s.i_tv80_core.BusA[4] ));
 sky130_fd_sc_hd__dfxtp_4 _6140_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net624),
    .Q(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__dfxtp_4 _6141_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net700),
    .Q(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6142_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net872),
    .Q(\z80.tv80s.i_tv80_core.BusA[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6143_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net266),
    .Q(\z80.tv80s.i_tv80_core.RegAddrA_r[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6144_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(net241),
    .Q(\z80.tv80s.i_tv80_core.RegAddrA_r[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6145_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net302),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6146_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0260_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6147_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net292),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6148_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net330),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6149_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net278),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6150_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0264_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6151_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net397),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6152_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net294),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][7] ));
 sky130_fd_sc_hd__dfstp_1 _6153_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net722),
    .SET_B(net173),
    .Q(net44));
 sky130_fd_sc_hd__dfrtp_4 _6154_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0267_),
    .RESET_B(net179),
    .Q(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6155_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(_0268_),
    .RESET_B(net180),
    .Q(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6156_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0269_),
    .RESET_B(net179),
    .Q(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6157_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net841),
    .RESET_B(net180),
    .Q(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6158_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0271_),
    .RESET_B(net179),
    .Q(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6159_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0272_),
    .RESET_B(net179),
    .Q(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6160_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0273_),
    .RESET_B(net179),
    .Q(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6161_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0274_),
    .RESET_B(net179),
    .Q(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__dfstp_1 _6162_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net498),
    .SET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.ts[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6163_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net717),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.ts[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6164_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net657),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.ts[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6165_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_0278_),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.ts[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6166_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(_0279_),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.ts[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6167_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net399),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.ts[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6168_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net256),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.ts[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6169_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net664),
    .RESET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.IntE ));
 sky130_fd_sc_hd__dfrtp_1 _6170_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net830),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.IntE_FF2 ));
 sky130_fd_sc_hd__dfrtp_1 _6171_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net620),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.Halt_FF ));
 sky130_fd_sc_hd__dfstp_4 _6172_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net867),
    .SET_B(net181),
    .Q(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__dfstp_4 _6173_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0283_),
    .SET_B(net181),
    .Q(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__dfstp_4 _6174_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net785),
    .SET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__dfstp_1 _6175_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(_0285_),
    .SET_B(net183),
    .Q(\z80.tv80s.i_tv80_core.F[3] ));
 sky130_fd_sc_hd__dfstp_4 _6176_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net834),
    .SET_B(net181),
    .Q(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__dfstp_2 _6177_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net794),
    .SET_B(net183),
    .Q(\z80.tv80s.i_tv80_core.F[5] ));
 sky130_fd_sc_hd__dfstp_2 _6178_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0288_),
    .SET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__dfstp_2 _6179_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net819),
    .SET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6180_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net589),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.I[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6181_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net630),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.I[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6182_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net567),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.I[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6183_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net616),
    .RESET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.I[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6184_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net645),
    .RESET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.I[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6185_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net598),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.I[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6186_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net550),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.I[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6187_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net579),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.I[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6188_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0298_),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.PC[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6189_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net730),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.PC[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6190_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net610),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.PC[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6191_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(net643),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.PC[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6192_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net649),
    .RESET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.PC[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6193_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net639),
    .RESET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.PC[5] ));
 sky130_fd_sc_hd__dfrtp_2 _6194_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net632),
    .RESET_B(net184),
    .Q(\z80.tv80s.i_tv80_core.PC[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6195_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net678),
    .RESET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.PC[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6196_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net779),
    .RESET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__dfrtp_4 _6197_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net762),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__dfrtp_4 _6198_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net754),
    .RESET_B(net184),
    .Q(\z80.tv80s.i_tv80_core.PC[10] ));
 sky130_fd_sc_hd__dfrtp_4 _6199_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net743),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.PC[11] ));
 sky130_fd_sc_hd__dfrtp_4 _6200_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net684),
    .RESET_B(net184),
    .Q(\z80.tv80s.i_tv80_core.PC[12] ));
 sky130_fd_sc_hd__dfrtp_4 _6201_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net708),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.PC[13] ));
 sky130_fd_sc_hd__dfrtp_2 _6202_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net612),
    .RESET_B(net184),
    .Q(\z80.tv80s.i_tv80_core.PC[14] ));
 sky130_fd_sc_hd__dfrtp_2 _6203_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net668),
    .RESET_B(net184),
    .Q(\z80.tv80s.i_tv80_core.PC[15] ));
 sky130_fd_sc_hd__dfstp_2 _6204_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net796),
    .SET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.SP[0] ));
 sky130_fd_sc_hd__dfstp_2 _6205_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net724),
    .SET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.SP[1] ));
 sky130_fd_sc_hd__dfstp_2 _6206_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net688),
    .SET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.SP[2] ));
 sky130_fd_sc_hd__dfstp_2 _6207_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net670),
    .SET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.SP[3] ));
 sky130_fd_sc_hd__dfstp_1 _6208_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net781),
    .SET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.SP[4] ));
 sky130_fd_sc_hd__dfstp_1 _6209_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net787),
    .SET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.SP[5] ));
 sky130_fd_sc_hd__dfstp_1 _6210_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net768),
    .SET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.SP[6] ));
 sky130_fd_sc_hd__dfstp_1 _6211_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net801),
    .SET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.SP[7] ));
 sky130_fd_sc_hd__dfstp_1 _6212_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net704),
    .SET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.SP[8] ));
 sky130_fd_sc_hd__dfstp_1 _6213_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net756),
    .SET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.SP[9] ));
 sky130_fd_sc_hd__dfstp_1 _6214_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net775),
    .SET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.SP[10] ));
 sky130_fd_sc_hd__dfstp_1 _6215_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net789),
    .SET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.SP[11] ));
 sky130_fd_sc_hd__dfstp_1 _6216_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net783),
    .SET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.SP[12] ));
 sky130_fd_sc_hd__dfstp_2 _6217_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net682),
    .SET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.SP[13] ));
 sky130_fd_sc_hd__dfstp_1 _6218_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net475),
    .SET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.SP[14] ));
 sky130_fd_sc_hd__dfstp_1 _6219_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net772),
    .SET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.SP[15] ));
 sky130_fd_sc_hd__dfstp_1 _6220_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net659),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.Ap[0] ));
 sky130_fd_sc_hd__dfstp_1 _6221_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net710),
    .SET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.Ap[1] ));
 sky130_fd_sc_hd__dfstp_1 _6222_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net655),
    .SET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.Ap[2] ));
 sky130_fd_sc_hd__dfstp_1 _6223_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net706),
    .SET_B(net181),
    .Q(\z80.tv80s.i_tv80_core.Ap[3] ));
 sky130_fd_sc_hd__dfstp_1 _6224_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net666),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.Ap[4] ));
 sky130_fd_sc_hd__dfstp_1 _6225_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net694),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.Ap[5] ));
 sky130_fd_sc_hd__dfstp_1 _6226_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net690),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.Ap[6] ));
 sky130_fd_sc_hd__dfstp_1 _6227_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net686),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.Ap[7] ));
 sky130_fd_sc_hd__dfstp_1 _6228_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net674),
    .SET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.Fp[0] ));
 sky130_fd_sc_hd__dfstp_1 _6229_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net696),
    .SET_B(net181),
    .Q(\z80.tv80s.i_tv80_core.Fp[1] ));
 sky130_fd_sc_hd__dfstp_1 _6230_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net647),
    .SET_B(net181),
    .Q(\z80.tv80s.i_tv80_core.Fp[2] ));
 sky130_fd_sc_hd__dfstp_1 _6231_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net622),
    .SET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.Fp[3] ));
 sky130_fd_sc_hd__dfstp_1 _6232_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net732),
    .SET_B(net181),
    .Q(\z80.tv80s.i_tv80_core.Fp[4] ));
 sky130_fd_sc_hd__dfstp_1 _6233_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net661),
    .SET_B(net181),
    .Q(\z80.tv80s.i_tv80_core.Fp[5] ));
 sky130_fd_sc_hd__dfstp_1 _6234_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net651),
    .SET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.Fp[6] ));
 sky130_fd_sc_hd__dfstp_1 _6235_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net692),
    .SET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.Fp[7] ));
 sky130_fd_sc_hd__dfstp_2 _6236_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0346_),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__dfstp_2 _6237_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0347_),
    .SET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__dfstp_2 _6238_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0348_),
    .SET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__dfstp_2 _6239_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net817),
    .SET_B(net181),
    .Q(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__dfstp_2 _6240_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0350_),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__dfstp_2 _6241_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net814),
    .SET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__dfstp_2 _6242_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(_0352_),
    .SET_B(net182),
    .Q(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__dfstp_2 _6243_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0353_),
    .SET_B(net183),
    .Q(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6244_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net554),
    .RESET_B(net183),
    .Q(net38));
 sky130_fd_sc_hd__dfrtp_1 _6245_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net533),
    .RESET_B(net183),
    .Q(net39));
 sky130_fd_sc_hd__dfrtp_1 _6246_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net535),
    .RESET_B(net181),
    .Q(net40));
 sky130_fd_sc_hd__dfrtp_1 _6247_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net573),
    .RESET_B(net181),
    .Q(net41));
 sky130_fd_sc_hd__dfrtp_1 _6248_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net552),
    .RESET_B(net181),
    .Q(net42));
 sky130_fd_sc_hd__dfrtp_1 _6249_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net541),
    .RESET_B(net181),
    .Q(net43));
 sky130_fd_sc_hd__dfrtp_1 _6250_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net593),
    .RESET_B(net183),
    .Q(net45));
 sky130_fd_sc_hd__dfrtp_1 _6251_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net604),
    .RESET_B(net183),
    .Q(net46));
 sky130_fd_sc_hd__dfrtp_1 _6252_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(net571),
    .RESET_B(net175),
    .Q(\z80.tv80s.i_tv80_core.IR[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6253_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(net858),
    .RESET_B(net175),
    .Q(\z80.tv80s.i_tv80_core.IR[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6254_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(net856),
    .RESET_B(net175),
    .Q(\z80.tv80s.i_tv80_core.IR[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6255_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(net843),
    .RESET_B(net175),
    .Q(\z80.tv80s.i_tv80_core.IR[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6256_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_0366_),
    .RESET_B(net175),
    .Q(\z80.tv80s.i_tv80_core.IR[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6257_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_0367_),
    .RESET_B(net175),
    .Q(\z80.tv80s.i_tv80_core.IR[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6258_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(net851),
    .RESET_B(net175),
    .Q(\z80.tv80s.i_tv80_core.IR[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6259_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(net839),
    .RESET_B(net175),
    .Q(\z80.tv80s.i_tv80_core.IR[7] ));
 sky130_fd_sc_hd__buf_1 _6293_ (.A(net21),
    .X(net14));
 sky130_fd_sc_hd__buf_1 _6294_ (.A(net21),
    .X(net15));
 sky130_fd_sc_hd__buf_1 _6295_ (.A(net21),
    .X(net16));
 sky130_fd_sc_hd__buf_1 _6296_ (.A(net21),
    .X(net17));
 sky130_fd_sc_hd__buf_1 _6297_ (.A(net21),
    .X(net18));
 sky130_fd_sc_hd__buf_1 _6298_ (.A(net21),
    .X(net19));
 sky130_fd_sc_hd__buf_1 _6299_ (.A(net21),
    .X(net20));
 sky130_fd_sc_hd__conb_1 ci2406_z80_185 (.LO(net185));
 sky130_fd_sc_hd__conb_1 ci2406_z80_186 (.LO(net186));
 sky130_fd_sc_hd__conb_1 ci2406_z80_187 (.LO(net187));
 sky130_fd_sc_hd__conb_1 ci2406_z80_188 (.LO(net188));
 sky130_fd_sc_hd__conb_1 ci2406_z80_189 (.LO(net189));
 sky130_fd_sc_hd__conb_1 ci2406_z80_190 (.LO(net190));
 sky130_fd_sc_hd__conb_1 ci2406_z80_191 (.LO(net191));
 sky130_fd_sc_hd__conb_1 ci2406_z80_192 (.LO(net192));
 sky130_fd_sc_hd__conb_1 ci2406_z80_193 (.LO(net193));
 sky130_fd_sc_hd__conb_1 ci2406_z80_194 (.LO(net194));
 sky130_fd_sc_hd__conb_1 ci2406_z80_195 (.LO(net195));
 sky130_fd_sc_hd__conb_1 ci2406_z80_196 (.LO(net196));
 sky130_fd_sc_hd__conb_1 ci2406_z80_197 (.LO(net197));
 sky130_fd_sc_hd__conb_1 ci2406_z80_198 (.LO(net198));
 sky130_fd_sc_hd__conb_1 ci2406_z80_199 (.LO(net199));
 sky130_fd_sc_hd__conb_1 ci2406_z80_200 (.LO(net200));
 sky130_fd_sc_hd__conb_1 ci2406_z80_201 (.LO(net201));
 sky130_fd_sc_hd__conb_1 ci2406_z80_202 (.LO(net202));
 sky130_fd_sc_hd__conb_1 ci2406_z80_203 (.LO(net203));
 sky130_fd_sc_hd__conb_1 ci2406_z80_204 (.LO(net204));
 sky130_fd_sc_hd__conb_1 ci2406_z80_205 (.LO(net205));
 sky130_fd_sc_hd__conb_1 ci2406_z80_206 (.LO(net206));
 sky130_fd_sc_hd__conb_1 ci2406_z80_207 (.LO(net207));
 sky130_fd_sc_hd__conb_1 ci2406_z80_208 (.LO(net208));
 sky130_fd_sc_hd__conb_1 ci2406_z80_209 (.LO(net209));
 sky130_fd_sc_hd__conb_1 ci2406_z80_210 (.LO(net210));
 sky130_fd_sc_hd__conb_1 ci2406_z80_211 (.LO(net211));
 sky130_fd_sc_hd__conb_1 ci2406_z80_212 (.LO(net212));
 sky130_fd_sc_hd__conb_1 ci2406_z80_213 (.HI(net213));
 sky130_fd_sc_hd__conb_1 ci2406_z80_214 (.HI(net214));
 sky130_fd_sc_hd__conb_1 ci2406_z80_215 (.HI(net215));
 sky130_fd_sc_hd__conb_1 ci2406_z80_216 (.HI(net216));
 sky130_fd_sc_hd__conb_1 ci2406_z80_217 (.HI(net217));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_37_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_39_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_40_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_41_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_42_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_43_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_44_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_45_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_46_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_47_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_48_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_49_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_50_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 fanout100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_8 fanout101 (.A(_0541_),
    .X(net101));
 sky130_fd_sc_hd__buf_4 fanout102 (.A(net103),
    .X(net102));
 sky130_fd_sc_hd__buf_8 fanout103 (.A(_0540_),
    .X(net103));
 sky130_fd_sc_hd__buf_6 fanout104 (.A(_0444_),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_8 fanout105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_8 fanout106 (.A(_0378_),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_8 fanout107 (.A(_0377_),
    .X(net107));
 sky130_fd_sc_hd__buf_4 fanout108 (.A(_2723_),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_8 fanout109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_8 fanout110 (.A(net114),
    .X(net110));
 sky130_fd_sc_hd__buf_6 fanout111 (.A(net114),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_8 fanout112 (.A(net114),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_4 fanout113 (.A(net114),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_8 fanout114 (.A(net33),
    .X(net114));
 sky130_fd_sc_hd__buf_6 fanout115 (.A(_2707_),
    .X(net115));
 sky130_fd_sc_hd__buf_6 fanout116 (.A(_2706_),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_8 fanout117 (.A(_2705_),
    .X(net117));
 sky130_fd_sc_hd__buf_4 fanout118 (.A(_2701_),
    .X(net118));
 sky130_fd_sc_hd__buf_4 fanout119 (.A(_2701_),
    .X(net119));
 sky130_fd_sc_hd__buf_4 fanout120 (.A(net121),
    .X(net120));
 sky130_fd_sc_hd__buf_2 fanout121 (.A(net122),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_8 fanout122 (.A(net797),
    .X(net122));
 sky130_fd_sc_hd__buf_4 fanout123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__buf_4 fanout124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__buf_4 fanout125 (.A(net791),
    .X(net125));
 sky130_fd_sc_hd__buf_4 fanout126 (.A(net130),
    .X(net126));
 sky130_fd_sc_hd__buf_4 fanout127 (.A(net128),
    .X(net127));
 sky130_fd_sc_hd__buf_4 fanout128 (.A(net130),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_8 fanout129 (.A(net130),
    .X(net129));
 sky130_fd_sc_hd__buf_2 fanout130 (.A(net842),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_8 fanout131 (.A(\z80.tv80s.i_tv80_core.IR[2] ),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_4 fanout132 (.A(net855),
    .X(net132));
 sky130_fd_sc_hd__buf_4 fanout133 (.A(\z80.tv80s.i_tv80_core.IR[1] ),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_4 fanout134 (.A(net857),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_8 fanout135 (.A(\z80.tv80s.i_tv80_core.IR[0] ),
    .X(net135));
 sky130_fd_sc_hd__buf_8 fanout136 (.A(net773),
    .X(net136));
 sky130_fd_sc_hd__buf_4 fanout137 (.A(\z80.tv80s.i_tv80_core.ts[3] ),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_4 fanout138 (.A(\z80.tv80s.i_tv80_core.ts[3] ),
    .X(net138));
 sky130_fd_sc_hd__buf_4 fanout139 (.A(net871),
    .X(net139));
 sky130_fd_sc_hd__buf_4 fanout140 (.A(net873),
    .X(net140));
 sky130_fd_sc_hd__buf_4 fanout141 (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ),
    .X(net141));
 sky130_fd_sc_hd__buf_4 fanout142 (.A(net869),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_8 fanout143 (.A(net144),
    .X(net143));
 sky130_fd_sc_hd__buf_4 fanout144 (.A(net860),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_8 fanout145 (.A(net146),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_8 fanout146 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ),
    .X(net146));
 sky130_fd_sc_hd__buf_4 fanout147 (.A(net149),
    .X(net147));
 sky130_fd_sc_hd__buf_4 fanout148 (.A(net149),
    .X(net148));
 sky130_fd_sc_hd__buf_4 fanout149 (.A(net151),
    .X(net149));
 sky130_fd_sc_hd__buf_4 fanout150 (.A(net151),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_4 fanout151 (.A(net809),
    .X(net151));
 sky130_fd_sc_hd__buf_6 fanout152 (.A(\z80.tv80s.i_tv80_core.RegAddrC[0] ),
    .X(net152));
 sky130_fd_sc_hd__buf_6 fanout153 (.A(net865),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_8 fanout154 (.A(net826),
    .X(net154));
 sky130_fd_sc_hd__buf_6 fanout155 (.A(net160),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_8 fanout156 (.A(net157),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_8 fanout157 (.A(net160),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_8 fanout158 (.A(net159),
    .X(net158));
 sky130_fd_sc_hd__buf_4 fanout159 (.A(net160),
    .X(net159));
 sky130_fd_sc_hd__buf_4 fanout160 (.A(net824),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_8 fanout161 (.A(\z80.tv80s.i_tv80_core.RegAddrC[1] ),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_8 fanout162 (.A(net864),
    .X(net162));
 sky130_fd_sc_hd__buf_6 fanout163 (.A(net805),
    .X(net163));
 sky130_fd_sc_hd__buf_6 fanout164 (.A(net167),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_8 fanout165 (.A(net167),
    .X(net165));
 sky130_fd_sc_hd__buf_2 fanout166 (.A(net167),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_4 fanout167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__buf_4 fanout168 (.A(\z80.tv80s.i_tv80_core.ISet[0] ),
    .X(net168));
 sky130_fd_sc_hd__buf_6 fanout169 (.A(net807),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_8 fanout170 (.A(net171),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_4 fanout171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__buf_4 fanout172 (.A(net13),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_8 fanout173 (.A(net176),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_8 fanout174 (.A(net175),
    .X(net174));
 sky130_fd_sc_hd__buf_4 fanout175 (.A(net176),
    .X(net175));
 sky130_fd_sc_hd__buf_4 fanout176 (.A(net13),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_8 fanout177 (.A(net184),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_8 fanout178 (.A(net184),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_8 fanout179 (.A(net180),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_8 fanout180 (.A(net183),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_8 fanout181 (.A(net183),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_8 fanout182 (.A(net183),
    .X(net182));
 sky130_fd_sc_hd__buf_6 fanout183 (.A(net184),
    .X(net183));
 sky130_fd_sc_hd__buf_4 fanout184 (.A(net13),
    .X(net184));
 sky130_fd_sc_hd__buf_6 fanout53 (.A(_1389_),
    .X(net53));
 sky130_fd_sc_hd__buf_6 fanout54 (.A(net55),
    .X(net54));
 sky130_fd_sc_hd__buf_6 fanout55 (.A(_0517_),
    .X(net55));
 sky130_fd_sc_hd__buf_4 fanout57 (.A(_1744_),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_8 fanout58 (.A(_0441_),
    .X(net58));
 sky130_fd_sc_hd__buf_6 fanout59 (.A(_2377_),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_8 fanout60 (.A(_1741_),
    .X(net60));
 sky130_fd_sc_hd__buf_2 fanout61 (.A(_1741_),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_8 fanout62 (.A(_2388_),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_8 fanout63 (.A(net64),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_8 fanout64 (.A(_1739_),
    .X(net64));
 sky130_fd_sc_hd__buf_4 fanout65 (.A(_0718_),
    .X(net65));
 sky130_fd_sc_hd__buf_4 fanout66 (.A(_2572_),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_8 fanout67 (.A(_1734_),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_8 fanout68 (.A(_1734_),
    .X(net68));
 sky130_fd_sc_hd__buf_4 fanout69 (.A(_0726_),
    .X(net69));
 sky130_fd_sc_hd__buf_4 fanout70 (.A(_0725_),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_8 fanout71 (.A(_0722_),
    .X(net71));
 sky130_fd_sc_hd__buf_4 fanout72 (.A(_0721_),
    .X(net72));
 sky130_fd_sc_hd__buf_4 fanout73 (.A(_1577_),
    .X(net73));
 sky130_fd_sc_hd__buf_4 fanout74 (.A(_0737_),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_8 fanout76 (.A(_2471_),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_8 fanout77 (.A(_0855_),
    .X(net77));
 sky130_fd_sc_hd__buf_2 fanout78 (.A(_0855_),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_8 fanout79 (.A(_0733_),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_8 fanout80 (.A(net81),
    .X(net80));
 sky130_fd_sc_hd__buf_6 fanout81 (.A(_0732_),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_8 fanout82 (.A(net85),
    .X(net82));
 sky130_fd_sc_hd__buf_4 fanout83 (.A(net85),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_4 fanout84 (.A(net85),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_4 fanout85 (.A(_0730_),
    .X(net85));
 sky130_fd_sc_hd__buf_4 fanout86 (.A(_1239_),
    .X(net86));
 sky130_fd_sc_hd__buf_4 fanout87 (.A(_1239_),
    .X(net87));
 sky130_fd_sc_hd__buf_4 fanout88 (.A(_1237_),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_8 fanout89 (.A(_0678_),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_8 fanout90 (.A(_0675_),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_4 fanout91 (.A(_0675_),
    .X(net91));
 sky130_fd_sc_hd__buf_4 fanout92 (.A(_1238_),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_8 fanout94 (.A(_2859_),
    .X(net94));
 sky130_fd_sc_hd__buf_4 fanout95 (.A(_2852_),
    .X(net95));
 sky130_fd_sc_hd__buf_4 fanout96 (.A(_2851_),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_8 fanout98 (.A(_1743_),
    .X(net98));
 sky130_fd_sc_hd__buf_4 fanout99 (.A(_1743_),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[6] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0225_),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][2] ),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(_0099_),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][5] ),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(_0126_),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][5] ),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_0110_),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][7] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_0112_),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][3] ),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_0132_),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[1] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][7] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_0080_),
    .X(net328));
 sky130_fd_sc_hd__buf_1 hold112 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][3] ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(_0262_),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_0127_),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_0036_),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][7] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_0043_),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0215_),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][4] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(_0050_),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_0153_),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(_0059_),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\z80.tv80s.i_tv80_core.mcycles[5] ),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_0016_),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_0107_),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[4] ),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(_0129_),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][6] ),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(_0151_),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_0134_),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_0061_),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0218_),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(_0092_),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_0060_),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_0058_),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][0] ),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_0097_),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][5] ),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_0118_),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][1] ),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[10] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(_0106_),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][0] ),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_0145_),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][7] ),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(_0071_),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_0040_),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_0062_),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][3] ),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_0224_),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(_0067_),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][6] ),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_0111_),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][3] ),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_0049_),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[0] ),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(_0086_),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][7] ),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][0] ),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[5] ),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_0073_),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][4] ),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_0149_),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][3] ),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(_0156_),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][5] ),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(_0069_),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_0056_),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][6] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_0219_),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(_0265_),
    .X(net397));
 sky130_fd_sc_hd__buf_2 hold181 (.A(\z80.tv80s.i_tv80_core.ts[4] ),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(_0280_),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(_0158_),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][2] ),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(_0094_),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][0] ),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[3] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(_0113_),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][1] ),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\z80.tv80s.i_tv80_core.Z16_r ),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(_0168_),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(_0124_),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[4] ),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][3] ),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(_0116_),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0220_),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_0217_),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(_0133_),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][1] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_0146_),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\z80.tv80s.i_tv80_core.mcycles[4] ),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(_0015_),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][4] ),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][4] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(_0157_),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(net877),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[8] ),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_0057_),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][7] ),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(_0063_),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][7] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(_0152_),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][5] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][0] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(_0105_),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0222_),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(_0095_),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(_0039_),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(_0159_),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][7] ),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][5] ),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(_0150_),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\z80.tv80s.i_tv80_core.RegAddrA_r[1] ),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(_0142_),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\z80.tv80s.i_tv80_core.Auto_Wait_t1 ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][4] ),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\z80.tv80s.i_tv80_core.mcycles[1] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(_0013_),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][3] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][1] ),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][0] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_0258_),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][7] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][7] ),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(_0160_),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[5] ),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(_0010_),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(_0143_),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][3] ),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(_0100_),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[15] ),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][7] ),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(_0104_),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][5] ),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][6] ),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ),
    .X(net472));
 sky130_fd_sc_hd__buf_1 hold256 (.A(\z80.tv80s.i_tv80_core.SP[14] ),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(_2614_),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(_0328_),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_0229_),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][6] ),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(_0119_),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][4] ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ),
    .X(net484));
 sky130_fd_sc_hd__buf_1 hold268 (.A(\z80.tv80s.i_tv80_core.IncDecZ ),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(_0213_),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\z80.tv80s.i_tv80_core.RegAddrA_r[2] ),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][6] ),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(_0042_),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[7] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(_0012_),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(_0084_),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][7] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(_0088_),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0044_),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\z80.tv80s.i_tv80_core.ts[6] ),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(_0275_),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][6] ),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][3] ),
    .X(net503));
 sky130_fd_sc_hd__buf_1 hold287 (.A(\z80.tv80s.i_tv80_core.NMI_s ),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(_0170_),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[12] ),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\z80.tv80s.i_tv80_core.XY_State[0] ),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(_0173_),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(_0121_),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][7] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(_0144_),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(_0089_),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\z80.tv80s.i_tv80_core.Auto_Wait_t2 ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(_0021_),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[7] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0226_),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\z80.tv80s.i_tv80_core.IStatus[1] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(_0004_),
    .X(net518));
 sky130_fd_sc_hd__clkbuf_2 hold302 (.A(\z80.tv80s.i_tv80_core.NMICycle ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(_0248_),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[0] ),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(_0122_),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(_0247_),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(net23),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[13] ),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(_0199_),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(net29),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(_0205_),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(net28),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(_0204_),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(net39),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(_0355_),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(net40),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(_0356_),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(net37),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0227_),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(_0212_),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(_0090_),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(net43),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(_0359_),
    .X(net541));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold325 (.A(net878),
    .X(net542));
 sky130_fd_sc_hd__buf_1 hold326 (.A(\z80.tv80s.i_tv80_core.PreserveC_r ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(_0055_),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(net25),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(_0201_),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[6] ),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(net27),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(_0203_),
    .X(net548));
 sky130_fd_sc_hd__buf_1 hold332 (.A(\z80.tv80s.i_tv80_core.I[6] ),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(_0296_),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(net42),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(_0358_),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(net38),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(_0354_),
    .X(net554));
 sky130_fd_sc_hd__clkbuf_4 hold338 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(net35),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0539_),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(_0210_),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(net52),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(_0198_),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(net32),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(_0208_),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(net36),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(_0211_),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(net26),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(_0202_),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\z80.tv80s.i_tv80_core.I[2] ),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(_0030_),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(_0292_),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(net24),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(_0200_),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\z80.tv80s.i_tv80_core.IR[0] ),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(_0362_),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(net41),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(_0357_),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(net30),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(_0206_),
    .X(net575));
 sky130_fd_sc_hd__buf_1 hold359 (.A(\z80.tv80s.i_tv80_core.XY_State[1] ),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[9] ),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(_0174_),
    .X(net577));
 sky130_fd_sc_hd__buf_1 hold361 (.A(\z80.tv80s.i_tv80_core.I[7] ),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(_0297_),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\z80.tv80s.i_tv80_core.BusB[0] ),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(_0231_),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(net34),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(_0209_),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[2] ),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(_0045_),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\z80.tv80s.i_tv80_core.ISet[1] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(_0223_),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(_0001_),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\z80.tv80s.i_tv80_core.I[0] ),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(_0290_),
    .X(net589));
 sky130_fd_sc_hd__buf_1 hold373 (.A(\z80.tv80s.i_tv80_core.BusB[4] ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(_0235_),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(net45),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(_0360_),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\z80.tv80s.i_tv80_core.mcycles[2] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(_0580_),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(_0014_),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\z80.tv80s.i_tv80_core.ts[5] ),
    .X(net255));
 sky130_fd_sc_hd__buf_1 hold380 (.A(\z80.tv80s.i_tv80_core.I[5] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(_0295_),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(net51),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(_0197_),
    .X(net600));
 sky130_fd_sc_hd__buf_1 hold384 (.A(\z80.tv80s.i_tv80_core.BusB[6] ),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(_0237_),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(net46),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(_0361_),
    .X(net604));
 sky130_fd_sc_hd__buf_1 hold388 (.A(\z80.tv80s.i_tv80_core.BusB[5] ),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(_0236_),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(_0281_),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(_0184_),
    .X(net608));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold392 (.A(\z80.tv80s.i_tv80_core.PC[2] ),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(_0300_),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\z80.tv80s.i_tv80_core.PC[14] ),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(_0312_),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(net31),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(_0207_),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(\z80.tv80s.i_tv80_core.I[3] ),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(_0293_),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0221_),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[1] ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(\z80.tv80s.i_tv80_core.BusA[3] ),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(_0252_),
    .X(net618));
 sky130_fd_sc_hd__buf_1 hold402 (.A(\z80.tv80s.i_tv80_core.Halt_FF ),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(_0024_),
    .X(net620));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold404 (.A(\z80.tv80s.i_tv80_core.F[3] ),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(_0341_),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\z80.tv80s.i_tv80_core.BusA[5] ),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(_0254_),
    .X(net624));
 sky130_fd_sc_hd__clkbuf_2 hold408 (.A(\z80.tv80s.i_tv80_core.BusB[7] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(_0238_),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_0006_),
    .X(net258));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold410 (.A(\z80.tv80s.i_tv80_core.BusB[3] ),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(_0234_),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(\z80.tv80s.i_tv80_core.I[1] ),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(_0291_),
    .X(net630));
 sky130_fd_sc_hd__buf_1 hold414 (.A(\z80.tv80s.i_tv80_core.PC[6] ),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(_0304_),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(_0253_),
    .X(net634));
 sky130_fd_sc_hd__clkbuf_2 hold418 (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\z80.tv80s.i_tv80_core.BusA[2] ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[2] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(_0251_),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\z80.tv80s.i_tv80_core.PC[5] ),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(_0303_),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(_0190_),
    .X(net641));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold425 (.A(\z80.tv80s.i_tv80_core.PC[3] ),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(_0301_),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\z80.tv80s.i_tv80_core.I[4] ),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(_0294_),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\z80.tv80s.i_tv80_core.Fp[2] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(_0007_),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(_0340_),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\z80.tv80s.i_tv80_core.PC[4] ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(_0302_),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\z80.tv80s.i_tv80_core.Fp[6] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(_0344_),
    .X(net651));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold435 (.A(\z80.tv80s.i_tv80_core.BusB[2] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(_0233_),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\z80.tv80s.i_tv80_core.Ap[2] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(_0332_),
    .X(net655));
 sky130_fd_sc_hd__buf_2 hold439 (.A(\z80.tv80s.i_tv80_core.ts[1] ),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[4] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(_0277_),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\z80.tv80s.i_tv80_core.Ap[0] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(_0330_),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\z80.tv80s.i_tv80_core.Fp[5] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(_0343_),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\z80.tv80s.i_tv80_core.IntE ),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(_0660_),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(_0026_),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(\z80.tv80s.i_tv80_core.Ap[4] ),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(_0334_),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_0009_),
    .X(net262));
 sky130_fd_sc_hd__buf_1 hold450 (.A(\z80.tv80s.i_tv80_core.PC[15] ),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(_0313_),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\z80.tv80s.i_tv80_core.SP[3] ),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(_0317_),
    .X(net670));
 sky130_fd_sc_hd__clkbuf_2 hold454 (.A(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(_0185_),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\z80.tv80s.i_tv80_core.Fp[0] ),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(_0338_),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\z80.tv80s.i_tv80_core.TmpAddr[15] ),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(_0191_),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\z80.tv80s.i_tv80_core.IStatus[2] ),
    .X(net263));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold460 (.A(\z80.tv80s.i_tv80_core.PC[7] ),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(_0305_),
    .X(net678));
 sky130_fd_sc_hd__clkbuf_2 hold462 (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(_0164_),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\z80.tv80s.i_tv80_core.SP[13] ),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(_0327_),
    .X(net682));
 sky130_fd_sc_hd__buf_1 hold466 (.A(\z80.tv80s.i_tv80_core.PC[12] ),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(_0310_),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\z80.tv80s.i_tv80_core.Ap[7] ),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(_0337_),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_0005_),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(\z80.tv80s.i_tv80_core.SP[2] ),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(_0316_),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\z80.tv80s.i_tv80_core.Ap[6] ),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(_0336_),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\z80.tv80s.i_tv80_core.Fp[7] ),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(_0345_),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\z80.tv80s.i_tv80_core.Ap[5] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(_0335_),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\z80.tv80s.i_tv80_core.Fp[1] ),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(_0339_),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\z80.tv80s.i_tv80_core.RegAddrA_r[0] ),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(_0187_),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\z80.tv80s.i_tv80_core.BusA[6] ),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(_0255_),
    .X(net700));
 sky130_fd_sc_hd__buf_1 hold484 (.A(\z80.tv80s.i_tv80_core.BusB[1] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(_0232_),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\z80.tv80s.i_tv80_core.SP[8] ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(_0322_),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\z80.tv80s.i_tv80_core.Ap[3] ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(_0333_),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(_0257_),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\z80.tv80s.i_tv80_core.PC[13] ),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(_0311_),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\z80.tv80s.i_tv80_core.Ap[1] ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(_0331_),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\z80.tv80s.i_tv80_core.Arith16_r ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(_0169_),
    .X(net712));
 sky130_fd_sc_hd__clkbuf_2 hold496 (.A(_0035_),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(_2165_),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(_0243_),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\z80.tv80s.i_tv80_core.ts[0] ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[14] ),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_2 hold50 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(_0276_),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(_0188_),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(net44),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(_0651_),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(_0032_),
    .X(net722));
 sky130_fd_sc_hd__buf_1 hold506 (.A(\z80.tv80s.i_tv80_core.SP[1] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(_0315_),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\z80.tv80s.i_tv80_core.BusA[0] ),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(_0249_),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_0029_),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(_0189_),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(\z80.tv80s.i_tv80_core.PC[1] ),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(_0299_),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(\z80.tv80s.i_tv80_core.Fp[4] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(_0342_),
    .X(net732));
 sky130_fd_sc_hd__buf_1 hold516 (.A(_0033_),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(_2160_),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(_2166_),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(_0244_),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\z80.tv80s.i_tv80_core.BTR_r ),
    .X(net269));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold520 (.A(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(_0186_),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(\z80.tv80s.i_tv80_core.BusA[1] ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(_0250_),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(\z80.tv80s.i_tv80_core.Alternate ),
    .X(net741));
 sky130_fd_sc_hd__buf_1 hold525 (.A(\z80.tv80s.i_tv80_core.PC[11] ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(_0309_),
    .X(net743));
 sky130_fd_sc_hd__buf_1 hold527 (.A(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(_0176_),
    .X(net745));
 sky130_fd_sc_hd__clkbuf_2 hold529 (.A(\z80.tv80s.i_tv80_core.IntCycle ),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(_0162_),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(_0172_),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\z80.tv80s.i_tv80_core.PC[0] ),
    .X(net748));
 sky130_fd_sc_hd__buf_2 hold532 (.A(\z80.tv80s.i_tv80_core.BusReq_s ),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(_0171_),
    .X(net750));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold534 (.A(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(_0183_),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(\z80.tv80s.i_tv80_core.PC[10] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(_0308_),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(\z80.tv80s.i_tv80_core.SP[9] ),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(_0323_),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][2] ),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(_0179_),
    .X(net758));
 sky130_fd_sc_hd__buf_1 hold542 (.A(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(_0178_),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_2 hold544 (.A(\z80.tv80s.i_tv80_core.PC[9] ),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(_0307_),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(_0180_),
    .X(net764));
 sky130_fd_sc_hd__buf_1 hold548 (.A(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(_0177_),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(_0066_),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(\z80.tv80s.i_tv80_core.SP[6] ),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(_0320_),
    .X(net768));
 sky130_fd_sc_hd__buf_1 hold552 (.A(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(_0182_),
    .X(net770));
 sky130_fd_sc_hd__buf_1 hold554 (.A(\z80.tv80s.i_tv80_core.SP[15] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(_0329_),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(\z80.tv80s.i_tv80_core.ts[3] ),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\z80.tv80s.i_tv80_core.SP[10] ),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(_0324_),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[3] ),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(_0181_),
    .X(net777));
 sky130_fd_sc_hd__buf_1 hold561 (.A(\z80.tv80s.i_tv80_core.PC[8] ),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(_0306_),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(\z80.tv80s.i_tv80_core.SP[4] ),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(_0318_),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\z80.tv80s.i_tv80_core.SP[12] ),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(_0326_),
    .X(net783));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold567 (.A(\z80.tv80s.i_tv80_core.F[2] ),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(_0284_),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\z80.tv80s.i_tv80_core.SP[5] ),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(_0008_),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(_0319_),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\z80.tv80s.i_tv80_core.SP[11] ),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(_0325_),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\z80.tv80s.i_tv80_core.BusB[3] ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(\z80.tv80s.i_tv80_core.IR[4] ),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(_0028_),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(\z80.tv80s.i_tv80_core.F[5] ),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(_0287_),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(\z80.tv80s.i_tv80_core.SP[0] ),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(_0314_),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][7] ),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(\z80.tv80s.i_tv80_core.IR[5] ),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(_0553_),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(_0000_),
    .X(net799));
 sky130_fd_sc_hd__buf_1 hold583 (.A(\z80.tv80s.i_tv80_core.SP[7] ),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(_0321_),
    .X(net801));
 sky130_fd_sc_hd__buf_1 hold585 (.A(_0034_),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(_2167_),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(_0245_),
    .X(net804));
 sky130_fd_sc_hd__clkbuf_2 hold588 (.A(\z80.tv80s.i_tv80_core.ISet[2] ),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(_0019_),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_0053_),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(\z80.tv80s.i_tv80_core.RegAddrC[2] ),
    .X(net807));
 sky130_fd_sc_hd__clkbuf_2 hold591 (.A(\z80.tv80s.i_tv80_core.ACC[7] ),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[0] ),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(\z80.tv80s.i_tv80_core.ACC[2] ),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(\z80.tv80s.i_tv80_core.ACC[4] ),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\z80.tv80s.i_tv80_core.ACC[6] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(\z80.tv80s.i_tv80_core.ACC[5] ),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(_0351_),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(\z80.tv80s.i_tv80_core.ACC[0] ),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\z80.tv80s.i_tv80_core.ACC[3] ),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0228_),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][4] ),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(_0349_),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\z80.tv80s.i_tv80_core.F[7] ),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(_0289_),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\z80.tv80s.i_tv80_core.ACC[1] ),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(_0242_),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(\z80.tv80s.i_tv80_core.F[6] ),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\z80.tv80s.i_tv80_core.BusAck ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(_0192_),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[1] ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(_0263_),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(_0193_),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\z80.tv80s.i_tv80_core.IntE_FF2 ),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(_0662_),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(_0027_),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(_0195_),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(\z80.tv80s.i_tv80_core.F[4] ),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(_0286_),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][1] ),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(_0161_),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\z80.tv80s.i_tv80_core.IR[7] ),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(_0369_),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\z80.tv80s.di_reg[3] ),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(_0270_),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\z80.tv80s.i_tv80_core.IR[3] ),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(_0365_),
    .X(net843));
 sky130_fd_sc_hd__buf_2 hold627 (.A(\z80.tv80s.i_tv80_core.ts[2] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\z80.tv80s.di_reg[4] ),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_0074_),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(\z80.tv80s.di_reg[6] ),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\z80.tv80s.di_reg[2] ),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(\z80.tv80s.di_reg[1] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\z80.tv80s.i_tv80_core.IR[6] ),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(_0368_),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(\z80.tv80s.di_reg[5] ),
    .X(net852));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold636 (.A(\z80.tv80s.di_reg[7] ),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\z80.tv80s.di_reg[0] ),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(\z80.tv80s.i_tv80_core.IR[2] ),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(_0364_),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][6] ),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(\z80.tv80s.i_tv80_core.IR[1] ),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(_0363_),
    .X(net858));
 sky130_fd_sc_hd__buf_1 hold642 (.A(\z80.tv80s.i_tv80_core.ts[2] ),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(_0241_),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\z80.tv80s.i_tv80_core.No_BTR ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(_0240_),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\z80.tv80s.i_tv80_core.RegAddrC[1] ),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(\z80.tv80s.i_tv80_core.RegAddrC[0] ),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\z80.tv80s.i_tv80_core.F[0] ),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_0079_),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(_0282_),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\z80.tv80s.i_tv80_core.F[1] ),
    .X(net868));
 sky130_fd_sc_hd__clkbuf_2 hold652 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(\z80.tv80s.i_tv80_core.ts[2] ),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(\z80.tv80s.i_tv80_core.BusA[7] ),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(_0256_),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\z80.tv80s.i_tv80_core.ts[6] ),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][1] ),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(_0816_),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][2] ),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][1] ),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[2] ),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(_0075_),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][4] ),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_0068_),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[2] ),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][4] ),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_0077_),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][5] ),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_0078_),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_0261_),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][7] ),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(_0266_),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][1] ),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(_0065_),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0216_),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][6] ),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(_0070_),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][3] ),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(_0076_),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(_0259_),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(_0046_),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_0115_),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[11] ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][1] ),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\z80.tv80s.i_tv80_core.ISet[3] ),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_0003_),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(_0048_),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][4] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_0117_),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][5] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_0051_),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(io_in[24]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(io_in[33]),
    .X(net10));
 sky130_fd_sc_hd__buf_4 input11 (.A(io_in[34]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(io_in[35]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input13 (.A(rst_n),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(io_in[25]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(io_in[26]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(io_in[27]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(io_in[28]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(io_in[29]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(io_in[30]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(io_in[31]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(io_in[32]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 max_cap56 (.A(_1746_),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 max_cap75 (.A(_0715_),
    .X(net75));
 sky130_fd_sc_hd__buf_2 max_cap97 (.A(_2768_),
    .X(net97));
 sky130_fd_sc_hd__buf_12 output14 (.A(net14),
    .X(io_oeb[24]));
 sky130_fd_sc_hd__buf_12 output15 (.A(net15),
    .X(io_oeb[25]));
 sky130_fd_sc_hd__buf_12 output16 (.A(net16),
    .X(io_oeb[26]));
 sky130_fd_sc_hd__buf_12 output17 (.A(net17),
    .X(io_oeb[27]));
 sky130_fd_sc_hd__buf_12 output18 (.A(net18),
    .X(io_oeb[28]));
 sky130_fd_sc_hd__buf_12 output19 (.A(net19),
    .X(io_oeb[29]));
 sky130_fd_sc_hd__buf_12 output20 (.A(net20),
    .X(io_oeb[30]));
 sky130_fd_sc_hd__buf_12 output21 (.A(net21),
    .X(io_oeb[31]));
 sky130_fd_sc_hd__buf_12 output22 (.A(net22),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_12 output23 (.A(net23),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_12 output24 (.A(net24),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_12 output25 (.A(net25),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_12 output26 (.A(net26),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_12 output27 (.A(net27),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_12 output28 (.A(net28),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_12 output29 (.A(net29),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_12 output30 (.A(net30),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_12 output31 (.A(net31),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_12 output32 (.A(net32),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_12 output33 (.A(net110),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_12 output34 (.A(net34),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_12 output35 (.A(net35),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_12 output36 (.A(net36),
    .X(io_out[22]));
 sky130_fd_sc_hd__buf_12 output37 (.A(net37),
    .X(io_out[23]));
 sky130_fd_sc_hd__buf_12 output38 (.A(net38),
    .X(io_out[24]));
 sky130_fd_sc_hd__buf_12 output39 (.A(net39),
    .X(io_out[25]));
 sky130_fd_sc_hd__buf_12 output40 (.A(net40),
    .X(io_out[26]));
 sky130_fd_sc_hd__buf_12 output41 (.A(net41),
    .X(io_out[27]));
 sky130_fd_sc_hd__buf_12 output42 (.A(net42),
    .X(io_out[28]));
 sky130_fd_sc_hd__buf_12 output43 (.A(net43),
    .X(io_out[29]));
 sky130_fd_sc_hd__buf_12 output44 (.A(net44),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_12 output45 (.A(net45),
    .X(io_out[30]));
 sky130_fd_sc_hd__buf_12 output46 (.A(net46),
    .X(io_out[31]));
 sky130_fd_sc_hd__buf_12 output47 (.A(net47),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_12 output48 (.A(net48),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_12 output49 (.A(net49),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_12 output50 (.A(net50),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_12 output51 (.A(net51),
    .X(io_out[8]));
 sky130_fd_sc_hd__buf_12 output52 (.A(net52),
    .X(io_out[9]));
 sky130_fd_sc_hd__clkbuf_2 wire93 (.A(_2882_),
    .X(net93));
 assign io_oeb[0] = net185;
 assign io_oeb[10] = net195;
 assign io_oeb[11] = net196;
 assign io_oeb[12] = net197;
 assign io_oeb[13] = net198;
 assign io_oeb[14] = net199;
 assign io_oeb[15] = net200;
 assign io_oeb[16] = net201;
 assign io_oeb[17] = net202;
 assign io_oeb[18] = net203;
 assign io_oeb[19] = net204;
 assign io_oeb[1] = net186;
 assign io_oeb[20] = net205;
 assign io_oeb[21] = net206;
 assign io_oeb[22] = net207;
 assign io_oeb[23] = net208;
 assign io_oeb[2] = net187;
 assign io_oeb[32] = net213;
 assign io_oeb[33] = net214;
 assign io_oeb[34] = net215;
 assign io_oeb[35] = net216;
 assign io_oeb[3] = net188;
 assign io_oeb[4] = net189;
 assign io_oeb[5] = net190;
 assign io_oeb[6] = net191;
 assign io_oeb[7] = net192;
 assign io_oeb[8] = net193;
 assign io_oeb[9] = net194;
 assign io_out[32] = net209;
 assign io_out[33] = net210;
 assign io_out[34] = net211;
 assign io_out[35] = net212;
 assign io_out[7] = net217;
endmodule

