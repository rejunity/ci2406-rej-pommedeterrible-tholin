* NGSPICE file created from execution_unit.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

.subckt execution_unit busy curr_PC[0] curr_PC[10] curr_PC[11] curr_PC[12] curr_PC[13]
+ curr_PC[14] curr_PC[15] curr_PC[16] curr_PC[17] curr_PC[18] curr_PC[19] curr_PC[1]
+ curr_PC[20] curr_PC[21] curr_PC[22] curr_PC[23] curr_PC[24] curr_PC[25] curr_PC[26]
+ curr_PC[27] curr_PC[2] curr_PC[3] curr_PC[4] curr_PC[5] curr_PC[6] curr_PC[7] curr_PC[8]
+ curr_PC[9] dest_idx[0] dest_idx[1] dest_idx[2] dest_idx[3] dest_idx[4] dest_idx[5]
+ dest_mask[0] dest_mask[1] dest_pred[0] dest_pred[1] dest_pred[2] dest_pred_val dest_val[0]
+ dest_val[10] dest_val[11] dest_val[12] dest_val[13] dest_val[14] dest_val[15] dest_val[16]
+ dest_val[17] dest_val[18] dest_val[19] dest_val[1] dest_val[20] dest_val[21] dest_val[22]
+ dest_val[23] dest_val[24] dest_val[25] dest_val[26] dest_val[27] dest_val[28] dest_val[29]
+ dest_val[2] dest_val[30] dest_val[31] dest_val[3] dest_val[4] dest_val[5] dest_val[6]
+ dest_val[7] dest_val[8] dest_val[9] instruction[0] instruction[10] instruction[11]
+ instruction[12] instruction[13] instruction[14] instruction[15] instruction[16]
+ instruction[17] instruction[18] instruction[19] instruction[1] instruction[20] instruction[21]
+ instruction[22] instruction[23] instruction[24] instruction[25] instruction[26]
+ instruction[27] instruction[28] instruction[29] instruction[2] instruction[30] instruction[31]
+ instruction[32] instruction[33] instruction[34] instruction[35] instruction[36]
+ instruction[37] instruction[38] instruction[39] instruction[3] instruction[40] instruction[41]
+ instruction[4] instruction[5] instruction[6] instruction[7] instruction[8] instruction[9]
+ int_return is_load is_store loadstore_address[0] loadstore_address[10] loadstore_address[11]
+ loadstore_address[12] loadstore_address[13] loadstore_address[14] loadstore_address[15]
+ loadstore_address[16] loadstore_address[17] loadstore_address[18] loadstore_address[19]
+ loadstore_address[1] loadstore_address[20] loadstore_address[21] loadstore_address[22]
+ loadstore_address[23] loadstore_address[24] loadstore_address[25] loadstore_address[26]
+ loadstore_address[27] loadstore_address[28] loadstore_address[29] loadstore_address[2]
+ loadstore_address[30] loadstore_address[31] loadstore_address[3] loadstore_address[4]
+ loadstore_address[5] loadstore_address[6] loadstore_address[7] loadstore_address[8]
+ loadstore_address[9] loadstore_dest[0] loadstore_dest[1] loadstore_dest[2] loadstore_dest[3]
+ loadstore_dest[4] loadstore_dest[5] loadstore_size[0] loadstore_size[1] new_PC[0]
+ new_PC[10] new_PC[11] new_PC[12] new_PC[13] new_PC[14] new_PC[15] new_PC[16] new_PC[17]
+ new_PC[18] new_PC[19] new_PC[1] new_PC[20] new_PC[21] new_PC[22] new_PC[23] new_PC[24]
+ new_PC[25] new_PC[26] new_PC[27] new_PC[2] new_PC[3] new_PC[4] new_PC[5] new_PC[6]
+ new_PC[7] new_PC[8] new_PC[9] pred_idx[0] pred_idx[1] pred_idx[2] pred_val reg1_idx[0]
+ reg1_idx[1] reg1_idx[2] reg1_idx[3] reg1_idx[4] reg1_idx[5] reg1_val[0] reg1_val[10]
+ reg1_val[11] reg1_val[12] reg1_val[13] reg1_val[14] reg1_val[15] reg1_val[16] reg1_val[17]
+ reg1_val[18] reg1_val[19] reg1_val[1] reg1_val[20] reg1_val[21] reg1_val[22] reg1_val[23]
+ reg1_val[24] reg1_val[25] reg1_val[26] reg1_val[27] reg1_val[28] reg1_val[29] reg1_val[2]
+ reg1_val[30] reg1_val[31] reg1_val[3] reg1_val[4] reg1_val[5] reg1_val[6] reg1_val[7]
+ reg1_val[8] reg1_val[9] reg2_idx[0] reg2_idx[1] reg2_idx[2] reg2_idx[3] reg2_idx[4]
+ reg2_idx[5] reg2_val[0] reg2_val[10] reg2_val[11] reg2_val[12] reg2_val[13] reg2_val[14]
+ reg2_val[15] reg2_val[16] reg2_val[17] reg2_val[18] reg2_val[19] reg2_val[1] reg2_val[20]
+ reg2_val[21] reg2_val[22] reg2_val[23] reg2_val[24] reg2_val[25] reg2_val[26] reg2_val[27]
+ reg2_val[28] reg2_val[29] reg2_val[2] reg2_val[30] reg2_val[31] reg2_val[3] reg2_val[4]
+ reg2_val[5] reg2_val[6] reg2_val[7] reg2_val[8] reg2_val[9] rst sign_extend take_branch
+ vccd1 vssd1 wb_clk_i
XFILLER_0_94_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09523__A2 _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06883_ _06672_/A _06882_/X _06870_/X vssd1 vssd1 vccd1 vccd1 _06883_/X sky130_fd_sc_hd__a21o_1
X_09671_ _09671_/A _09672_/B vssd1 vssd1 vccd1 vccd1 _09671_/Y sky130_fd_sc_hd__nor2_1
X_08622_ _08611_/Y _08620_/Y _08621_/Y _08603_/X vssd1 vssd1 vccd1 vccd1 _08624_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_77_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12815__C1 _13147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08553_ _08553_/A _08553_/B vssd1 vssd1 vccd1 vccd1 _08556_/A sky130_fd_sc_hd__or2_1
XANTENNA__09287__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout162_A _12322_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08484_ _09404_/S _08484_/B vssd1 vssd1 vccd1 vccd1 _08524_/A sky130_fd_sc_hd__or2_1
X_07504_ _07505_/B _07505_/A vssd1 vssd1 vccd1 vccd1 _07504_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__09287__B2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10841__A1 _11868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07435_ _07435_/A _07435_/B vssd1 vssd1 vccd1 vccd1 _07440_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10974__A _10974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10841__B2 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07366_ _07366_/A _07366_/B vssd1 vssd1 vccd1 vccd1 _07368_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11397__A2 _07171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07297_ _10246_/A _07297_/B vssd1 vssd1 vccd1 vccd1 _07298_/B sky130_fd_sc_hd__or2_1
XFILLER_0_33_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09105_ _07172_/Y _08877_/B fanout6/X _09325_/A vssd1 vssd1 vccd1 vccd1 _09106_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_32_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09036_ _09037_/A _09549_/A vssd1 vssd1 vccd1 vccd1 _09036_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07470__B1 _07238_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06812__A3 _12650_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10357__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10109__B1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09938_ _09938_/A _09938_/B vssd1 vssd1 vccd1 vccd1 _09939_/B sky130_fd_sc_hd__or2_1
XANTENNA__07773__B2 _08627_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07773__A1 _08641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10214__A _11179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09869_ _09869_/A _09869_/B vssd1 vssd1 vccd1 vccd1 _09909_/B sky130_fd_sc_hd__or2_2
X_12880_ _12878_/X _12880_/B vssd1 vssd1 vccd1 vccd1 _13225_/A sky130_fd_sc_hd__nand2b_1
X_11900_ _06860_/A _11898_/X _11899_/Y vssd1 vssd1 vccd1 vccd1 _11900_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _06984_/B _09257_/S _11830_/X _06698_/Y vssd1 vssd1 vccd1 vccd1 _11831_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _11762_/A _11762_/B vssd1 vssd1 vccd1 vccd1 _11763_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_95_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12821__A2 _13101_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11693_ _11785_/A _11693_/B vssd1 vssd1 vccd1 vccd1 _11695_/B sky130_fd_sc_hd__nor2_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10713_ _07097_/X _07417_/B fanout42/X _07256_/Y vssd1 vssd1 vccd1 vccd1 _10714_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10832__A1 _10950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10644_ _10645_/A _10645_/B _10645_/C vssd1 vssd1 vccd1 vccd1 _10646_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10575_ _10165_/S _10164_/X _09251_/A vssd1 vssd1 vccd1 vccd1 _10575_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_63_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13363_ _13365_/CLK _13363_/D vssd1 vssd1 vccd1 vccd1 hold295/A sky130_fd_sc_hd__dfxtp_1
X_12314_ _12313_/A _12313_/B _12313_/Y _09225_/Y vssd1 vssd1 vccd1 vccd1 _12331_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09884__S _10297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09450__A1 _07554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09450__B2 _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08253__A2 _10221_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13294_ _13296_/CLK _13294_/D vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__dfxtp_1
X_12245_ _12300_/B _12299_/A vssd1 vssd1 vccd1 vccd1 _12350_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12176_ _12177_/A _12177_/B _12177_/C vssd1 vssd1 vccd1 vccd1 _12178_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__09753__A2 _09257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11127_ _11809_/A _08751_/A _08751_/B _08751_/C vssd1 vssd1 vccd1 vccd1 _11127_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__07764__A1 _08540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07764__B2 _08515_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07417__B _07417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11058_ _11058_/A _11058_/B vssd1 vssd1 vccd1 vccd1 _11060_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_64_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10009_ _11630_/A _10010_/B _10010_/C vssd1 vssd1 vccd1 vccd1 _10009_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__08529__A _08664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13065__A2 _13101_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12273__B1 _11554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12485__S _12520_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07220_ _07283_/A _06972_/C _07117_/C _07133_/A _07215_/B vssd1 vssd1 vccd1 vccd1
+ _07221_/B sky130_fd_sc_hd__o41ai_4
XFILLER_0_27_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07151_ reg1_val[24] _08870_/C _07585_/B1 reg1_val[25] vssd1 vssd1 vccd1 vccd1 _07155_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_42_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09441__A1 _09440_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07082_ _09944_/A _07082_/B vssd1 vssd1 vccd1 vccd1 _07442_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12514__A _12680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07608__A _07608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12233__B _12233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout105 _07299_/X vssd1 vssd1 vccd1 vccd1 _09479_/B1 sky130_fd_sc_hd__buf_8
Xfanout138 _09794_/A vssd1 vssd1 vccd1 vccd1 _10207_/A sky130_fd_sc_hd__buf_12
Xfanout127 _07135_/X vssd1 vssd1 vccd1 vccd1 _08561_/B1 sky130_fd_sc_hd__clkbuf_8
X_07984_ _07985_/B _07985_/C _08664_/A vssd1 vssd1 vccd1 vccd1 _07988_/A sky130_fd_sc_hd__a21oi_1
Xfanout149 _07037_/X vssd1 vssd1 vccd1 vccd1 _08649_/A2 sky130_fd_sc_hd__buf_8
X_06935_ instruction[18] _06590_/X _06934_/X _06716_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[0]
+ sky130_fd_sc_hd__o211a_4
X_09723_ _09721_/X _09722_/X _10295_/S vssd1 vssd1 vccd1 vccd1 _09723_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_97_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06866_ reg1_val[29] _06866_/B vssd1 vssd1 vccd1 vccd1 _06877_/A sky130_fd_sc_hd__nand2_1
X_09654_ _09653_/B _09653_/C _09653_/A vssd1 vssd1 vccd1 vccd1 _09655_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08605_ _08605_/A _08605_/B vssd1 vssd1 vccd1 vccd1 _08677_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__06730__A2 _12796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06797_ reg2_val[3] _06810_/B vssd1 vssd1 vccd1 vccd1 _06797_/X sky130_fd_sc_hd__and2_2
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09585_ reg1_val[1] _07149_/A _07959_/A _12642_/A vssd1 vssd1 vccd1 vccd1 _09586_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08536_ _08557_/A _08557_/B _08532_/X vssd1 vssd1 vccd1 vccd1 _08543_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_49_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08467_ _08467_/A _08467_/B _08467_/C vssd1 vssd1 vccd1 vccd1 _08687_/B sky130_fd_sc_hd__and3_1
XFILLER_0_108_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12016__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08398_ _08406_/B _08406_/A vssd1 vssd1 vccd1 vccd1 _08399_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07418_ _09779_/A _07418_/B vssd1 vssd1 vccd1 vccd1 _07420_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_107_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07349_ _07349_/A _07349_/B vssd1 vssd1 vccd1 vccd1 _07353_/A sky130_fd_sc_hd__xor2_1
XANTENNA__10209__A _10209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10360_ _12224_/A _10360_/B vssd1 vssd1 vccd1 vccd1 _10362_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_5_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10291_ _10291_/A _10291_/B vssd1 vssd1 vccd1 vccd1 _10291_/Y sky130_fd_sc_hd__nand2_1
X_09019_ _08900_/A _08900_/B _08899_/A vssd1 vssd1 vccd1 vccd1 _09029_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_14_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12030_ _12030_/A _12030_/B _12030_/C vssd1 vssd1 vccd1 vccd1 _12031_/B sky130_fd_sc_hd__nand3_1
Xhold170 hold170/A vssd1 vssd1 vccd1 vccd1 hold170/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09196__A0 _09218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold181 hold181/A vssd1 vssd1 vccd1 vccd1 hold181/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 hold192/A vssd1 vssd1 vccd1 vccd1 hold192/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09499__A1 _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09499__B2 _09669_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12932_ hold94/X hold288/A vssd1 vssd1 vccd1 vccd1 _13158_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__10598__B _12087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07253__A _10749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12863_ _07051_/X _12863_/A2 hold61/X _13246_/A vssd1 vssd1 vccd1 vccd1 _13292_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13047__A2 _12820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ _11814_/A _11814_/B vssd1 vssd1 vccd1 vccd1 _11814_/Y sky130_fd_sc_hd__xnor2_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12255__B1 _11637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12794_ _12791_/B _12793_/B _12789_/X vssd1 vssd1 vccd1 vccd1 _12795_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _10159_/A _10803_/X _11733_/B _09222_/Y _11744_/X vssd1 vssd1 vccd1 vccd1
+ _11745_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_56_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09120__B1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08474__A2 _08561_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11676_ _12009_/A fanout23/X fanout15/X fanout58/X vssd1 vssd1 vccd1 vccd1 _11677_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_83_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10627_ _10627_/A _10627_/B vssd1 vssd1 vccd1 vccd1 _10631_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10558_ reg1_val[9] curr_PC[9] vssd1 vssd1 vccd1 vccd1 _10558_/Y sky130_fd_sc_hd__nor2_1
X_13346_ _13396_/CLK hold102/X vssd1 vssd1 vccd1 vccd1 hold100/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10033__A2 _12144_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09974__A2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13277_ _13392_/CLK _13277_/D vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12334__A _12335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10489_ _12157_/A _10489_/B vssd1 vssd1 vccd1 vccd1 _10498_/A sky130_fd_sc_hd__xnor2_1
X_12228_ _12228_/A vssd1 vssd1 vccd1 vccd1 _12230_/B sky130_fd_sc_hd__inv_2
X_12159_ _07158_/X _12158_/B _12158_/Y _12224_/A vssd1 vssd1 vccd1 vccd1 _12161_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07147__B _07147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12089__A3 _12084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06986__B _07014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06720_ reg1_val[17] _07097_/A vssd1 vssd1 vccd1 vccd1 _06721_/B sky130_fd_sc_hd__nand2b_1
X_06651_ reg1_val[25] _06998_/A vssd1 vssd1 vccd1 vccd1 _06652_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13038__A2 _13254_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06582_ instruction[41] vssd1 vssd1 vccd1 vccd1 _06582_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_87_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09370_ _09371_/A _09371_/B vssd1 vssd1 vccd1 vccd1 _09370_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08321_ _08328_/B _08328_/A vssd1 vssd1 vccd1 vccd1 _08321_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_24_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08252_ _08454_/A _08252_/B vssd1 vssd1 vccd1 vccd1 _08255_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07203_ _07191_/X _07195_/X _10725_/A _07202_/Y vssd1 vssd1 vccd1 vccd1 _07204_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09414__A1 _12064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08183_ _08779_/A _08790_/B vssd1 vssd1 vccd1 vccd1 _08183_/X sky130_fd_sc_hd__or2_1
X_07134_ _08613_/B _08613_/C vssd1 vssd1 vccd1 vccd1 _07134_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_42_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07065_ reg1_val[6] _07065_/B vssd1 vssd1 vccd1 vccd1 _07073_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07338__A _10479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07967_ _07918_/A _07918_/B _07915_/Y vssd1 vssd1 vccd1 vccd1 _07970_/B sky130_fd_sc_hd__o21bai_1
X_06918_ _06783_/A _06610_/X _09239_/B instruction[4] _06917_/Y vssd1 vssd1 vccd1
+ vccd1 _12805_/B sky130_fd_sc_hd__a221oi_4
X_09706_ _09707_/A _09707_/B vssd1 vssd1 vccd1 vccd1 _09706_/X sky130_fd_sc_hd__and2_1
XANTENNA__07073__A _09947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07898_ _09677_/A _08112_/B fanout25/X _07172_/Y vssd1 vssd1 vccd1 vccd1 _07899_/B
+ sky130_fd_sc_hd__o22a_1
X_06849_ reg1_val[16] _07094_/A vssd1 vssd1 vccd1 vccd1 _06849_/Y sky130_fd_sc_hd__nand2_1
X_09637_ _09638_/A _09638_/B vssd1 vssd1 vccd1 vccd1 _09850_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09568_ _09566_/X _09567_/X _10295_/S vssd1 vssd1 vccd1 vccd1 _09568_/X sky130_fd_sc_hd__mux2_1
X_08519_ _08553_/A _08523_/B _08512_/Y vssd1 vssd1 vccd1 vccd1 _08522_/B sky130_fd_sc_hd__a21bo_1
X_11530_ _11335_/X _11712_/A _11529_/X vssd1 vssd1 vccd1 vccd1 _11530_/X sky130_fd_sc_hd__a21o_1
XANTENNA__11996__C1 _12421_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11460__A1 _09221_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09499_ _09301_/A fanout14/X fanout13/X _09669_/B2 vssd1 vssd1 vccd1 vccd1 _09500_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_108_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11461_ hold204/A _11461_/B vssd1 vssd1 vccd1 vccd1 _11557_/B sky130_fd_sc_hd__or2_1
XANTENNA__11748__C1 _11747_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13200_ hold274/X _13223_/A2 _13199_/X _13223_/B2 vssd1 vssd1 vccd1 vccd1 _13201_/B
+ sky130_fd_sc_hd__a22o_1
X_11392_ _12233_/B _07131_/Y fanout46/X _12233_/A vssd1 vssd1 vccd1 vccd1 _11393_/B
+ sky130_fd_sc_hd__o22a_1
X_10412_ _10413_/A _10413_/B _10413_/C vssd1 vssd1 vccd1 vccd1 _10538_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08632__A _09673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10343_ _10343_/A _10343_/B vssd1 vssd1 vccd1 vccd1 _10344_/B sky130_fd_sc_hd__nand2_1
X_13131_ hold260/X _13254_/A2 _13130_/X _06577_/A vssd1 vssd1 vccd1 vccd1 hold261/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11366__A1_N _09221_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10274_ _10274_/A _10274_/B vssd1 vssd1 vccd1 vccd1 _10275_/B sky130_fd_sc_hd__xor2_4
X_13062_ hold82/X _13094_/A2 _13101_/A2 _13341_/Q _13259_/A vssd1 vssd1 vccd1 vccd1
+ hold83/A sky130_fd_sc_hd__o221a_1
X_12013_ _12013_/A _12013_/B vssd1 vssd1 vccd1 vccd1 _12033_/A sky130_fd_sc_hd__and2_1
XANTENNA__08144__B2 _09940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08144__A1 _09770_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12915_ _13110_/A _13111_/A _13110_/B vssd1 vssd1 vccd1 vccd1 _13116_/A sky130_fd_sc_hd__a21bo_1
X_12846_ hold96/X _12862_/B vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__or2_1
XFILLER_0_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06972__D _07117_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12777_ reg1_val[28] _12790_/B vssd1 vssd1 vccd1 vccd1 _12778_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_126_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11728_ reg1_val[20] curr_PC[20] vssd1 vssd1 vccd1 vccd1 _11730_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_83_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11659_ curr_PC[19] _11749_/C _12471_/S vssd1 vssd1 vccd1 vccd1 _11659_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12400__B1 _11892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11754__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13329_ _13360_/CLK _13329_/D vssd1 vssd1 vccd1 vccd1 hold119/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11506__A2 _12017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12999__A _13001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06997__A _06998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08870_ reg1_val[28] reg1_val[29] _08870_/C _12779_/B vssd1 vssd1 vccd1 vccd1 _08985_/B
+ sky130_fd_sc_hd__or4_1
X_07821_ _07874_/A _07874_/B vssd1 vssd1 vccd1 vccd1 _07877_/A sky130_fd_sc_hd__nand2_1
X_07752_ _07752_/A _07752_/B vssd1 vssd1 vccd1 vccd1 _07754_/B sky130_fd_sc_hd__xnor2_2
X_06703_ _06703_/A _12660_/B vssd1 vssd1 vccd1 vccd1 _06703_/Y sky130_fd_sc_hd__nor2_1
X_07683_ fanout72/X _08484_/B _09479_/B1 _10595_/A1 vssd1 vssd1 vccd1 vccd1 _07684_/B
+ sky130_fd_sc_hd__o22a_1
X_06634_ _06703_/A _12719_/B vssd1 vssd1 vccd1 vccd1 _06634_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12219__B1 _12631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09422_ _09728_/S _09422_/B _12644_/A vssd1 vssd1 vccd1 vccd1 _09422_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_35_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09353_ _09354_/A _09354_/B vssd1 vssd1 vccd1 vccd1 _09355_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11978__C1 _12359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout242_A _12471_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08304_ _08598_/B _10221_/B2 _09770_/B2 _08538_/A1 vssd1 vssd1 vccd1 vccd1 _08305_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07110__A2 _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10245__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09284_ _09284_/A _09284_/B vssd1 vssd1 vccd1 vccd1 _09286_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08235_ _08235_/A _08235_/B vssd1 vssd1 vccd1 vccd1 _08272_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09548__A _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08166_ _08227_/B _08227_/A vssd1 vssd1 vccd1 vccd1 _08166_/Y sky130_fd_sc_hd__nand2b_1
X_07117_ _12438_/A _07147_/B _07117_/C vssd1 vssd1 vccd1 vccd1 _07133_/B sky130_fd_sc_hd__and3_1
XFILLER_0_43_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08097_ _08098_/A _08098_/B vssd1 vssd1 vccd1 vccd1 _08097_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_101_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07048_ _07070_/A _07048_/B _07048_/C vssd1 vssd1 vccd1 vccd1 _08973_/D sky130_fd_sc_hd__or3_4
X_08999_ _09000_/A _09000_/B vssd1 vssd1 vccd1 vccd1 _08999_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12458__B1 _06958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10222__A _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08126__B2 _08613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08126__A1 _06992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10961_ _10962_/A _10962_/B vssd1 vssd1 vccd1 vccd1 _10963_/A sky130_fd_sc_hd__and2_1
XFILLER_0_97_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11752__S _11752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12700_ _12705_/B _12700_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[11] sky130_fd_sc_hd__and2_4
X_10892_ _10892_/A _10892_/B vssd1 vssd1 vccd1 vccd1 _10894_/B sky130_fd_sc_hd__xor2_1
X_12631_ reg1_val[26] curr_PC[26] _12631_/S vssd1 vssd1 vccd1 vccd1 _12633_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_38_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12562_ _11242_/A curr_PC[15] _12638_/S vssd1 vssd1 vccd1 vccd1 _12564_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_80_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11513_ _11514_/A _11514_/B vssd1 vssd1 vccd1 vccd1 _11612_/A sky130_fd_sc_hd__or2_1
X_12493_ _12665_/B _12494_/B vssd1 vssd1 vccd1 vccd1 _12504_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_65_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13186__B2 _13223_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11444_ _11630_/A _11444_/B _11444_/C vssd1 vssd1 vccd1 vccd1 _11444_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_104_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10944__B1 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11375_ curr_PC[16] curr_PC[17] _11375_/C vssd1 vssd1 vccd1 vccd1 _11564_/B sky130_fd_sc_hd__and3_1
XFILLER_0_1_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13114_ _13147_/A _13114_/B vssd1 vssd1 vccd1 vccd1 _13363_/D sky130_fd_sc_hd__and2_1
X_10326_ _11893_/A _10453_/A vssd1 vssd1 vccd1 vccd1 _10326_/X sky130_fd_sc_hd__or2_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10257_ _10257_/A _10257_/B _10257_/C vssd1 vssd1 vccd1 vccd1 _10259_/A sky130_fd_sc_hd__and3_1
X_13045_ _09673_/A _12820_/B hold40/X vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__a21oi_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12331__B _12331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10188_ _10135_/A _10135_/B _10133_/X vssd1 vssd1 vccd1 vccd1 _10276_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__06847__A_N _07262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06695__A2_N _06766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10475__A2 _07608_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12829_ _07232_/X _12871_/A2 hold23/X _13246_/A vssd1 vssd1 vccd1 vccd1 _13275_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09093__A2 _10476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08020_ _08540_/B _08457_/A2 _08501_/B1 _08515_/A2 vssd1 vssd1 vccd1 vccd1 _08021_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_25_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout7 fanout8/X vssd1 vssd1 vccd1 vccd1 fanout7/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__10935__B1 _11752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09971_ _11770_/A _09971_/B vssd1 vssd1 vccd1 vccd1 _09973_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08922_ _08807_/B _08920_/X _08921_/X _08805_/X _08919_/X vssd1 vssd1 vccd1 vccd1
+ _10138_/A sky130_fd_sc_hd__o221a_2
XFILLER_0_110_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12522__A _12685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout192_A _12416_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11360__B1 _12421_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08853_ _08854_/A _08854_/B vssd1 vssd1 vccd1 vccd1 _08943_/B sky130_fd_sc_hd__or2_1
XANTENNA__11138__A _11138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08784_ _11893_/B _08784_/B vssd1 vssd1 vccd1 vccd1 _08784_/Y sky130_fd_sc_hd__nand2_1
X_07804_ _07804_/A _07804_/B vssd1 vssd1 vccd1 vccd1 _07807_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13101__B2 _13101_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09305__B1 _09672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07735_ _07735_/A _07735_/B vssd1 vssd1 vccd1 vccd1 _07737_/B sky130_fd_sc_hd__and2_1
XANTENNA__11663__A1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11663__B2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09405_ _09403_/X _09404_/X _09725_/S vssd1 vssd1 vccd1 vccd1 _10022_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07331__A2 _10473_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07666_ _07666_/A _07666_/B vssd1 vssd1 vccd1 vccd1 _07667_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__07351__A _09922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06617_ _06927_/A _06617_/B vssd1 vssd1 vccd1 vccd1 _06617_/Y sky130_fd_sc_hd__nand2_1
X_07597_ _09325_/A _07362_/B fanout16/X _12808_/A vssd1 vssd1 vccd1 vccd1 _07598_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09336_ _09336_/A _09336_/B vssd1 vssd1 vccd1 vccd1 _09352_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08292__B1 fanout72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ _07175_/A _10337_/A _07238_/Y _07554_/B vssd1 vssd1 vccd1 vccd1 _09268_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08218_ _08218_/A _08218_/B vssd1 vssd1 vccd1 vccd1 _08222_/B sky130_fd_sc_hd__and2_1
XANTENNA__12376__C1 _12376_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09198_ _09194_/X _09197_/X _09725_/S vssd1 vssd1 vccd1 vccd1 _09198_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10926__B1 _12376_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08149_ _10207_/A _08149_/B vssd1 vssd1 vccd1 vccd1 _08220_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08044__B1 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11160_ curr_PC[13] _11159_/C curr_PC[14] vssd1 vssd1 vccd1 vccd1 _11161_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11091_ _11476_/A _07362_/B fanout16/X _11406_/A vssd1 vssd1 vccd1 vccd1 _11092_/B
+ sky130_fd_sc_hd__o22a_1
X_10111_ _10112_/A _10112_/B vssd1 vssd1 vccd1 vccd1 _10113_/A sky130_fd_sc_hd__and2_1
XFILLER_0_31_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10042_ _09225_/Y _10014_/Y _10016_/Y _12379_/B2 _10041_/X vssd1 vssd1 vccd1 vccd1
+ _10042_/X sky130_fd_sc_hd__a221o_1
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12578__S _12638_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11993_ _11650_/B _12068_/B hold254/A vssd1 vssd1 vccd1 vccd1 _11993_/Y sky130_fd_sc_hd__a21oi_1
X_10944_ _11592_/A fanout43/X fanout41/X _10944_/B2 vssd1 vssd1 vccd1 vccd1 _10945_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11654__A1 _07078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07261__A _07262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07858__B1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10875_ _10875_/A _10875_/B vssd1 vssd1 vccd1 vccd1 _10877_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12614_ _12621_/B _12614_/B vssd1 vssd1 vccd1 vccd1 new_PC[22] sky130_fd_sc_hd__xnor2_4
XFILLER_0_54_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12545_ _12546_/A _12546_/B _12546_/C vssd1 vssd1 vccd1 vccd1 _12553_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_93_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12476_ _12476_/A _12476_/B _12476_/C vssd1 vssd1 vccd1 vccd1 _12477_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_53_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08092__A _08575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ _11322_/A _11322_/B _11323_/Y vssd1 vssd1 vccd1 vccd1 _11429_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_111_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_5 instruction[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11358_ hold292/A _11650_/B _11549_/C _12376_/C1 vssd1 vssd1 vccd1 vccd1 _11359_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07389__A2 _10599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10309_ _10179_/A _10176_/Y _10178_/B vssd1 vssd1 vccd1 vccd1 _10313_/A sky130_fd_sc_hd__o21a_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11289_ _11387_/A _11289_/B vssd1 vssd1 vccd1 vccd1 _11291_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_67_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13028_ hold229/A _13223_/B2 _13209_/A2 hold224/X vssd1 vssd1 vccd1 vccd1 hold225/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11342__B1 _12356_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07520_ _09947_/A _07520_/B vssd1 vssd1 vccd1 vccd1 _07526_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07171__A _07171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09370__B _09371_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07451_ _07451_/A _07451_/B vssd1 vssd1 vccd1 vccd1 _07530_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07382_ fanout86/X fanout76/X fanout72/X fanout82/X vssd1 vssd1 vccd1 vccd1 _07383_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09121_ _11770_/A _09121_/B vssd1 vssd1 vccd1 vccd1 _09122_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__13112__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09052_ _09922_/A _09052_/B vssd1 vssd1 vccd1 vccd1 _09053_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_114_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08003_ _08003_/A _08003_/B vssd1 vssd1 vccd1 vccd1 _08004_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout205_A _07604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10908__B1 _10788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10384__A1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10384__B2 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09954_ fanout58/X fanout78/X fanout74/X _11868_/A vssd1 vssd1 vccd1 vccd1 _09955_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_0_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09885_ _09739_/X _09884_/X _11138_/A vssd1 vssd1 vccd1 vccd1 _09885_/X sky130_fd_sc_hd__mux2_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08905_ _08904_/A _08904_/B _08906_/A vssd1 vssd1 vccd1 vccd1 _08905_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10687__A2 _11990_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _10749_/A _08836_/B vssd1 vssd1 vccd1 vccd1 _08840_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_99_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07552__A2 _09325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08767_ _11538_/B _11538_/C vssd1 vssd1 vccd1 vccd1 _11630_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10500__A _10500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07718_ _08501_/B1 _08289_/B fanout75/X _10221_/B2 vssd1 vssd1 vccd1 vccd1 _07719_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07304__A2 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08698_ _08176_/Y _08180_/Y _08181_/X _08790_/A _08794_/A vssd1 vssd1 vccd1 vccd1
+ _08698_/X sky130_fd_sc_hd__a2111o_1
XANTENNA__08501__A1 _08613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07649_ fanout80/X fanout78/X fanout76/X fanout74/X vssd1 vssd1 vccd1 vccd1 _07650_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08501__B2 _06992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10660_ _10328_/Y _10902_/A _10658_/X vssd1 vssd1 vccd1 vccd1 _10660_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout20_A _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09319_ _09319_/A _09319_/B vssd1 vssd1 vccd1 vccd1 _09321_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_118_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10591_ _10592_/B _10591_/B vssd1 vssd1 vccd1 vccd1 _10593_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_63_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12330_ _12322_/Y _12323_/X _12326_/X _12329_/Y vssd1 vssd1 vccd1 vccd1 _12330_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13010__B1 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12261_ reg1_val[27] curr_PC[27] vssd1 vssd1 vccd1 vccd1 _12262_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11050__B _11050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11212_ _11212_/A _11212_/B vssd1 vssd1 vccd1 vccd1 _11214_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12192_ _12134_/A _12131_/Y _12133_/B vssd1 vssd1 vccd1 vccd1 _12192_/X sky130_fd_sc_hd__o21a_1
X_11143_ hold270/A _11143_/B vssd1 vssd1 vccd1 vccd1 _11255_/B sky130_fd_sc_hd__or2_1
X_11074_ _12096_/A _11074_/B vssd1 vssd1 vccd1 vccd1 _11076_/B sky130_fd_sc_hd__xor2_2
XANTENNA__07791__A2 _08289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10025_ _11028_/S _10023_/Y _10024_/X vssd1 vssd1 vccd1 vccd1 _10025_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07543__A2 _07959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11976_ _11809_/A _08784_/Y _08786_/Y _10788_/A vssd1 vssd1 vccd1 vccd1 _11977_/B
+ sky130_fd_sc_hd__a31o_1
X_10927_ _12420_/A0 _09422_/B _10927_/S vssd1 vssd1 vccd1 vccd1 _10927_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10858_ _10858_/A _10858_/B vssd1 vssd1 vccd1 vccd1 _10866_/A sky130_fd_sc_hd__xor2_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07141__D _07143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09048__A2 _07362_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12052__A1 _11892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10789_ _11630_/A _08735_/Y _08737_/Y _10788_/Y vssd1 vssd1 vccd1 vccd1 _10818_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_5_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08256__B1 _09940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12528_ _12689_/B _12529_/B vssd1 vssd1 vccd1 vccd1 _12539_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11241__A _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12459_ _12437_/Y _12441_/X _12457_/X _12458_/X vssd1 vssd1 vccd1 vccd1 dest_val[31]
+ sky130_fd_sc_hd__o31a_4
XFILLER_0_41_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08559__B2 _08613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08559__A1 _06992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11563__B1 _11562_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06951_ _09226_/B _09237_/B vssd1 vssd1 vccd1 vccd1 _09221_/B sky130_fd_sc_hd__or2_4
X_09670_ _09670_/A _09670_/B vssd1 vssd1 vccd1 vccd1 _09672_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06882_ _06672_/B _06864_/Y _06871_/X vssd1 vssd1 vccd1 vccd1 _06882_/X sky130_fd_sc_hd__a21o_1
X_08621_ _08603_/A _08603_/B _08610_/A _08603_/D vssd1 vssd1 vccd1 vccd1 _08621_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_89_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13107__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08552_ _08552_/A _08552_/B vssd1 vssd1 vccd1 vccd1 _08553_/B sky130_fd_sc_hd__and2_1
XANTENNA__09287__A2 _09943_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08483_ _08483_/A _08483_/B vssd1 vssd1 vccd1 vccd1 _08498_/A sky130_fd_sc_hd__xnor2_1
X_07503_ _07503_/A _07503_/B vssd1 vssd1 vccd1 vccd1 _07505_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_119_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout155_A _09669_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07434_ _07434_/A _07434_/B vssd1 vssd1 vccd1 vccd1 _07435_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10974__B _12017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10841__A2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08247__B1 fanout72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07365_ _07589_/A _07365_/B vssd1 vssd1 vccd1 vccd1 _07366_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07296_ _10246_/A _07297_/B vssd1 vssd1 vccd1 vccd1 _07298_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09104_ _08982_/A _08982_/B _08980_/X vssd1 vssd1 vccd1 vccd1 _09108_/A sky130_fd_sc_hd__o21ai_2
X_09035_ _07675_/X _08915_/X _08916_/X vssd1 vssd1 vccd1 vccd1 _09035_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_60_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09556__A _10049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10357__B2 _11406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10357__A1 _11476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10109__A1 _10944_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09937_ _09938_/A _09938_/B vssd1 vssd1 vccd1 vccd1 _09939_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07773__A2 _09661_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11306__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10109__B2 _07097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09868_ _10331_/A _09868_/B _09868_/C vssd1 vssd1 vccd1 vccd1 _09869_/B sky130_fd_sc_hd__and3_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ _09799_/A _09799_/B vssd1 vssd1 vccd1 vccd1 _09800_/B sky130_fd_sc_hd__nand2_1
X_08819_ _09779_/A _08819_/B vssd1 vssd1 vccd1 vccd1 _08821_/B sky130_fd_sc_hd__xor2_1
X_11830_ _11829_/A _09422_/B _11829_/Y _12421_/A1 vssd1 vssd1 vccd1 vccd1 _11830_/X
+ sky130_fd_sc_hd__o211a_1
X_11761_ _11760_/B _11761_/B vssd1 vssd1 vccd1 vccd1 _11762_/B sky130_fd_sc_hd__nand2b_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07015__S _09302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _11929_/A _10712_/B vssd1 vssd1 vccd1 vccd1 _10715_/A sky130_fd_sc_hd__xnor2_1
X_11692_ _11692_/A _11692_/B _11692_/C vssd1 vssd1 vccd1 vccd1 _11693_/B sky130_fd_sc_hd__and3_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10643_ _10643_/A _10643_/B vssd1 vssd1 vccd1 vccd1 _10645_/C sky130_fd_sc_hd__xor2_1
XANTENNA__12157__A _12157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08238__B1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10574_ _10566_/Y _10567_/X _10573_/X vssd1 vssd1 vccd1 vccd1 _10574_/Y sky130_fd_sc_hd__o21ai_1
X_13362_ _13365_/CLK _13362_/D vssd1 vssd1 vccd1 vccd1 hold235/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12313_ _12313_/A _12313_/B vssd1 vssd1 vccd1 vccd1 _12313_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09450__A2 _07232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13293_ _13296_/CLK _13293_/D vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__dfxtp_1
X_12244_ _12244_/A _12244_/B vssd1 vssd1 vccd1 vccd1 _12430_/A sky130_fd_sc_hd__nand2_2
X_12175_ _12175_/A _12175_/B vssd1 vssd1 vccd1 vccd1 _12177_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_48_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11126_ _11052_/X _11124_/Y _11125_/Y vssd1 vssd1 vccd1 vccd1 _11126_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07764__A2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11057_ _11055_/A _11055_/B _11058_/B vssd1 vssd1 vccd1 vccd1 _11207_/A sky130_fd_sc_hd__a21o_1
XANTENNA__08713__A1 _08664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10008_ _09910_/Y _10324_/A _10007_/Y vssd1 vssd1 vccd1 vccd1 _10008_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11959_ _11959_/A _11959_/B vssd1 vssd1 vccd1 vccd1 _11960_/B sky130_fd_sc_hd__or2_1
XFILLER_0_86_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10284__B1 _12356_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08477__B1 _08576_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07150_ _11134_/A _11242_/A _07141_/C _07143_/A _07585_/B1 vssd1 vssd1 vccd1 vccd1
+ _07167_/B sky130_fd_sc_hd__o41a_1
XFILLER_0_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07081_ _09943_/B2 fanout53/X _09650_/A fanout51/X vssd1 vssd1 vccd1 vccd1 _07082_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_120_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12328__A2 _11995_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07608__B _07608_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12233__C _12335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout117 _07198_/Y vssd1 vssd1 vccd1 vccd1 _10338_/B2 sky130_fd_sc_hd__buf_8
Xfanout106 _08484_/B vssd1 vssd1 vccd1 vccd1 _10473_/B2 sky130_fd_sc_hd__buf_6
Xfanout128 _07135_/X vssd1 vssd1 vccd1 vccd1 _09822_/A sky130_fd_sc_hd__clkbuf_4
X_09722_ _09390_/X _09400_/X _09727_/S vssd1 vssd1 vccd1 vccd1 _09722_/X sky130_fd_sc_hd__mux2_1
X_07983_ _07983_/A _07983_/B vssd1 vssd1 vccd1 vccd1 _07985_/C sky130_fd_sc_hd__nand2_1
X_06934_ instruction[25] _06944_/B vssd1 vssd1 vccd1 vccd1 _06934_/X sky130_fd_sc_hd__or2_1
XANTENNA__11839__A1 _11752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout272_A _06675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06865_ reg1_val[30] _08860_/A vssd1 vssd1 vccd1 vccd1 _06865_/X sky130_fd_sc_hd__and2_1
X_09653_ _09653_/A _09653_/B _09653_/C vssd1 vssd1 vccd1 vccd1 _09655_/A sky130_fd_sc_hd__and3_1
X_09584_ hold237/A _12322_/A1 _09582_/X _12205_/B1 vssd1 vssd1 vccd1 vccd1 _09584_/X
+ sky130_fd_sc_hd__a31o_1
X_08604_ _08596_/A _08596_/B _08596_/C _08603_/X vssd1 vssd1 vccd1 vccd1 _08677_/A
+ sky130_fd_sc_hd__a31o_1
X_06796_ _06796_/A _06796_/B vssd1 vssd1 vccd1 vccd1 _06898_/C sky130_fd_sc_hd__nand2_2
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08535_ _08535_/A _08535_/B vssd1 vssd1 vccd1 vccd1 _08557_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08466_ _08491_/A _08491_/B vssd1 vssd1 vccd1 vccd1 _08467_/C sky130_fd_sc_hd__nand2_1
XANTENNA__12016__B2 _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12016__A1 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08397_ _08397_/A _08397_/B vssd1 vssd1 vccd1 vccd1 _08406_/B sky130_fd_sc_hd__xor2_2
X_07417_ _07959_/A _07417_/B vssd1 vssd1 vccd1 vccd1 _07418_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09968__B1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07348_ _07349_/A _07349_/B vssd1 vssd1 vccd1 vccd1 _07655_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_122_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10578__A1 _12365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07279_ _07626_/A _07279_/B vssd1 vssd1 vccd1 vccd1 _07292_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_115_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10290_ _10291_/A _10291_/B vssd1 vssd1 vccd1 vccd1 _10290_/X sky130_fd_sc_hd__or2_1
XANTENNA__08190__A _08564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09018_ _09018_/A _09018_/B vssd1 vssd1 vccd1 vccd1 _09031_/A sky130_fd_sc_hd__xor2_4
Xhold171 hold171/A vssd1 vssd1 vccd1 vccd1 hold171/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold160 hold160/A vssd1 vssd1 vccd1 vccd1 hold160/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10225__A _10225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold182 hold182/A vssd1 vssd1 vccd1 vccd1 hold182/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 hold193/A vssd1 vssd1 vccd1 vccd1 hold193/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09499__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12931_ _13153_/A _13154_/A _13153_/B vssd1 vssd1 vccd1 vccd1 _13159_/A sky130_fd_sc_hd__a21bo_1
X_12862_ hold60/X _12862_/B vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__or2_1
X_11813_ _11811_/X _11812_/X _11813_/S vssd1 vssd1 vccd1 vccd1 _11814_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _12793_/A _12793_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[30] sky130_fd_sc_hd__xnor2_4
XANTENNA__09120__A1 _10234_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11744_ _07016_/A _09257_/S _11743_/X _06691_/X vssd1 vssd1 vccd1 vccd1 _11744_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09120__B2 _10725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11675_ _11675_/A _11675_/B vssd1 vssd1 vccd1 vccd1 _11687_/A sky130_fd_sc_hd__nand2_1
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10626_ _10627_/A _10627_/B vssd1 vssd1 vccd1 vccd1 _10709_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_64_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10557_ _10429_/A _10426_/Y _10428_/B vssd1 vssd1 vccd1 vccd1 _10561_/A sky130_fd_sc_hd__o21a_1
X_13345_ _13358_/CLK hold81/X vssd1 vssd1 vccd1 vccd1 _13345_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08631__B1 _07173_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13276_ _13392_/CLK _13276_/D vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__dfxtp_1
X_10488_ _10974_/A fanout23/X fanout15/X _10595_/A1 vssd1 vssd1 vccd1 vccd1 _10489_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12227_ _12336_/A _12227_/B vssd1 vssd1 vccd1 vccd1 _12228_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12158_ _12158_/A _12158_/B vssd1 vssd1 vccd1 vccd1 _12158_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07147__C _07959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11109_ _11109_/A _11109_/B vssd1 vssd1 vccd1 vccd1 _11111_/B sky130_fd_sc_hd__xnor2_1
X_12089_ _12009_/A _12335_/B _12084_/B _12013_/A vssd1 vssd1 vccd1 vccd1 _12103_/A
+ sky130_fd_sc_hd__o31ai_2
XANTENNA__11892__C _12049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_12_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13398_/CLK sky130_fd_sc_hd__clkbuf_8
X_06650_ _06998_/A reg1_val[25] vssd1 vssd1 vccd1 vccd1 _12143_/S sky130_fd_sc_hd__and2b_1
XFILLER_0_59_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06581_ _12642_/A vssd1 vssd1 vccd1 vccd1 _06581_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08320_ _08320_/A _08320_/B vssd1 vssd1 vccd1 vccd1 _08328_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08251_ _08561_/A2 _08484_/B _09479_/B1 _08561_/B1 vssd1 vssd1 vccd1 vccd1 _08252_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07202_ _11381_/A _07192_/B _07200_/X vssd1 vssd1 vccd1 vccd1 _07202_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_40_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08182_ _08182_/A _08182_/B vssd1 vssd1 vccd1 vccd1 _08790_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_70_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07133_ _07133_/A _07133_/B vssd1 vssd1 vccd1 vccd1 _08613_/C sky130_fd_sc_hd__and2_2
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07064_ _07083_/C _07083_/D _07248_/A vssd1 vssd1 vccd1 vccd1 _07065_/B sky130_fd_sc_hd__o21a_1
XANTENNA__07619__A _09944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09834__A _09834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07966_ _07966_/A _08062_/A vssd1 vssd1 vccd1 vccd1 _07996_/A sky130_fd_sc_hd__or2_1
X_06917_ instruction[6] instruction[5] instruction[4] vssd1 vssd1 vccd1 vccd1 _06917_/Y
+ sky130_fd_sc_hd__a21oi_2
X_09705_ _09707_/A _09707_/B vssd1 vssd1 vccd1 vccd1 _09705_/X sky130_fd_sc_hd__or2_1
XFILLER_0_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09636_ _09636_/A _09636_/B vssd1 vssd1 vccd1 vccd1 _09638_/B sky130_fd_sc_hd__xnor2_1
X_07897_ _07897_/A _07897_/B vssd1 vssd1 vccd1 vccd1 _08000_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_97_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06848_ _11239_/A _06846_/X _06847_/X vssd1 vssd1 vccd1 vccd1 _06848_/X sky130_fd_sc_hd__o21ba_1
X_06779_ reg1_val[6] _07283_/A vssd1 vssd1 vccd1 vccd1 _06779_/X sky130_fd_sc_hd__and2_1
X_09567_ _09181_/X _09202_/X _09727_/S vssd1 vssd1 vccd1 vccd1 _09567_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09498_ _09498_/A _09498_/B vssd1 vssd1 vccd1 vccd1 _09507_/A sky130_fd_sc_hd__xnor2_1
X_08518_ _08518_/A _08518_/B vssd1 vssd1 vccd1 vccd1 _08523_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08449_ _08449_/A _08449_/B vssd1 vssd1 vccd1 vccd1 _08450_/B sky130_fd_sc_hd__or2_1
XFILLER_0_108_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08861__B1 _08859_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11460_ _09221_/Y _11455_/B _11459_/X vssd1 vssd1 vccd1 vccd1 _11460_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11271__D_N _11124_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11391_ _12096_/A _11391_/B vssd1 vssd1 vccd1 vccd1 _11395_/A sky130_fd_sc_hd__xor2_1
X_10411_ _10411_/A _10411_/B vssd1 vssd1 vccd1 vccd1 _10413_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_45_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10342_ _10343_/A _10343_/B vssd1 vssd1 vccd1 vccd1 _10468_/B sky130_fd_sc_hd__or2_1
X_13130_ hold248/X _13129_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13130_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13061_ _10748_/A _13101_/B2 hold99/X vssd1 vssd1 vccd1 vccd1 _13340_/D sky130_fd_sc_hd__o21a_1
X_12012_ _12012_/A _12012_/B _12012_/C vssd1 vssd1 vccd1 vccd1 _12013_/B sky130_fd_sc_hd__or3_1
X_10273_ _10274_/A _10274_/B vssd1 vssd1 vccd1 vccd1 _10273_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10723__A1 _07269_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11920__B1 _11895_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10723__B2 _07262_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07264__A _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08144__A2 _08484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12914_ hold70/X hold235/X vssd1 vssd1 vccd1 vccd1 _13110_/B sky130_fd_sc_hd__nand2b_1
X_12845_ _07983_/B _12863_/A2 hold122/X _13210_/A vssd1 vssd1 vccd1 vccd1 _13283_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10239__B1 _10473_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12776_ reg1_val[28] _12790_/B vssd1 vssd1 vccd1 vccd1 _12787_/A sky130_fd_sc_hd__and2_1
XFILLER_0_29_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11727_ _11726_/A _11726_/B _11726_/Y _09225_/Y vssd1 vssd1 vccd1 vccd1 _11747_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11233__B _11271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11658_ _11627_/X _11628_/Y _11631_/Y _10788_/A _11657_/X vssd1 vssd1 vccd1 vccd1
+ _11658_/X sky130_fd_sc_hd__o221a_1
X_11589_ _11946_/C _11589_/B vssd1 vssd1 vccd1 vccd1 _11591_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_114_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10609_ _10609_/A _10609_/B vssd1 vssd1 vccd1 vccd1 _10611_/B sky130_fd_sc_hd__xor2_1
XANTENNA__10564__S _11820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13328_ _13392_/CLK hold139/X vssd1 vssd1 vccd1 vccd1 hold137/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13259_ _13259_/A _13259_/B hold128/X vssd1 vssd1 vccd1 vccd1 hold129/A sky130_fd_sc_hd__and3_1
XANTENNA__12080__A _12631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07820_ _07820_/A _07820_/B vssd1 vssd1 vccd1 vccd1 _07874_/B sky130_fd_sc_hd__xnor2_1
X_07751_ _07751_/A _07751_/B vssd1 vssd1 vccd1 vccd1 _07754_/A sky130_fd_sc_hd__xor2_2
X_06702_ instruction[29] _06716_/B vssd1 vssd1 vccd1 vccd1 _12660_/B sky130_fd_sc_hd__and2_4
XFILLER_0_126_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07682_ _07682_/A _07682_/B vssd1 vssd1 vccd1 vccd1 _07703_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_126_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06633_ instruction[40] _06675_/B vssd1 vssd1 vccd1 vccd1 _12719_/B sky130_fd_sc_hd__and2_4
X_09421_ _09418_/Y _09419_/Y _09420_/Y vssd1 vssd1 vccd1 vccd1 _09429_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09352_ _09352_/A _09352_/B vssd1 vssd1 vccd1 vccd1 _09354_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08303_ _08454_/A _08303_/B vssd1 vssd1 vccd1 vccd1 _08306_/A sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout235_A _09423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11442__A2 _11840_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09283_ _09079_/A _09078_/Y _09074_/Y vssd1 vssd1 vccd1 vccd1 _09284_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_28_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08234_ _08234_/A _08234_/B vssd1 vssd1 vccd1 vccd1 _08282_/A sky130_fd_sc_hd__xor2_4
XANTENNA__09548__B _09548_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08165_ _08165_/A _08165_/B vssd1 vssd1 vccd1 vccd1 _08227_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_27_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07116_ _07168_/A _07168_/B vssd1 vssd1 vccd1 vccd1 _07116_/X sky130_fd_sc_hd__and2_2
XFILLER_0_30_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08096_ _08098_/A _08098_/B vssd1 vssd1 vccd1 vccd1 _08096_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_100_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07047_ _07070_/A _07048_/B _07048_/C vssd1 vssd1 vccd1 vccd1 _07315_/A sky130_fd_sc_hd__nor3_4
XFILLER_0_101_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12702__B _12702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10181__A2 _10165_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07582__B1 _10599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08998_ _08998_/A _08998_/B vssd1 vssd1 vccd1 vccd1 _09000_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__12458__A1 _07147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08126__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07949_ _07948_/A _07948_/B _07948_/C vssd1 vssd1 vccd1 vccd1 _07950_/B sky130_fd_sc_hd__a21o_1
XANTENNA_fanout50_A _11484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ _11582_/A _10960_/B vssd1 vssd1 vccd1 vccd1 _10962_/B sky130_fd_sc_hd__xnor2_1
X_10891_ _10892_/A _10892_/B vssd1 vssd1 vccd1 vccd1 _11006_/A sky130_fd_sc_hd__nand2_1
X_09619_ _09619_/A _09619_/B vssd1 vssd1 vccd1 vccd1 _09621_/C sky130_fd_sc_hd__or2_1
X_12630_ _12630_/A _12630_/B vssd1 vssd1 vccd1 vccd1 new_PC[25] sky130_fd_sc_hd__xnor2_4
XFILLER_0_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12561_ _12567_/B _12561_/B vssd1 vssd1 vccd1 vccd1 new_PC[14] sky130_fd_sc_hd__and2_4
XFILLER_0_81_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11512_ _11419_/A _11418_/B _11416_/X vssd1 vssd1 vccd1 vccd1 _11514_/B sky130_fd_sc_hd__a21oi_1
X_12492_ reg1_val[5] curr_PC[5] _12520_/S vssd1 vssd1 vccd1 vccd1 _12494_/B sky130_fd_sc_hd__mux2_1
XANTENNA__13186__A2 _13223_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11443_ _11377_/Y _11840_/C _11442_/Y vssd1 vssd1 vccd1 vccd1 _11443_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_34_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10944__A1 _11592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10944__B2 _10944_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13113_ hold295/X _13254_/A2 _13112_/X _06577_/A vssd1 vssd1 vccd1 vccd1 _13114_/B
+ sky130_fd_sc_hd__a22o_1
X_11374_ curr_PC[16] _11375_/C curr_PC[17] vssd1 vssd1 vccd1 vccd1 _11374_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10325_ _10581_/A _10581_/B vssd1 vssd1 vccd1 vccd1 _10453_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_0_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10256_ _10255_/B _10255_/C _10255_/A vssd1 vssd1 vccd1 vccd1 _10257_/C sky130_fd_sc_hd__o21ai_1
X_13044_ _06576_/Y _06577_/A _13254_/A2 hold39/X rst vssd1 vssd1 vccd1 vccd1 hold40/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__09474__A _11946_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10187_ _10049_/B _10147_/Y _10049_/A vssd1 vssd1 vccd1 vccd1 _10187_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_88_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12828_ hold22/X _12870_/B vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__or2_1
XFILLER_0_57_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09093__A3 _10476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12759_ _12764_/A _12759_/B vssd1 vssd1 vccd1 vccd1 _12763_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_17_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout8 fanout8/A vssd1 vssd1 vccd1 vccd1 fanout8/X sky130_fd_sc_hd__buf_6
XFILLER_0_110_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09970_ _07097_/X fanout32/X fanout30/X _07256_/Y vssd1 vssd1 vccd1 vccd1 _09971_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08921_ _08799_/B _08799_/C _09037_/A _08920_/B vssd1 vssd1 vccd1 vccd1 _08921_/X
+ sky130_fd_sc_hd__a211o_1
X_08852_ _09667_/A _08852_/B vssd1 vssd1 vccd1 vccd1 _08854_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07803_ _07822_/A _07822_/B _07783_/X vssd1 vssd1 vccd1 vccd1 _07810_/B sky130_fd_sc_hd__a21bo_1
X_08783_ _08783_/A _08783_/B vssd1 vssd1 vccd1 vccd1 _08784_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_79_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07734_ _07734_/A _07734_/B _07734_/C vssd1 vssd1 vccd1 vccd1 _07735_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07665_ _07663_/A _07663_/B _07666_/B vssd1 vssd1 vccd1 vccd1 _07665_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__07632__A _09834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11663__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06616_ instruction[24] _12796_/A _06927_/B instruction[41] _06612_/X vssd1 vssd1
+ vccd1 vccd1 _06617_/B sky130_fd_sc_hd__a221o_1
X_09404_ _09185_/X _09211_/X _09404_/S vssd1 vssd1 vccd1 vccd1 _09404_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07596_ _07596_/A _07596_/B vssd1 vssd1 vccd1 vccd1 _07596_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_47_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08816__B1 _07221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09335_ _09335_/A _09335_/B vssd1 vssd1 vccd1 vccd1 _09336_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08292__A1 _06992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09266_ _09936_/A _09266_/B vssd1 vssd1 vccd1 vccd1 _09270_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08217_ _08217_/A _08217_/B vssd1 vssd1 vccd1 vccd1 _08218_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08292__B2 _08613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09197_ _09195_/X _09196_/X _09419_/B vssd1 vssd1 vccd1 vccd1 _09197_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07079__A _07080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08044__B2 _08649_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08044__A1 _08657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08148_ _08561_/A2 _08411_/B _10476_/A _08561_/B1 vssd1 vssd1 vccd1 vccd1 _08149_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_113_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08079_ _08079_/A _08079_/B vssd1 vssd1 vccd1 vccd1 _08165_/A sky130_fd_sc_hd__nand2_2
X_11090_ _12017_/A _11090_/B vssd1 vssd1 vccd1 vccd1 _11096_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10110_ _11484_/A _10110_/B vssd1 vssd1 vccd1 vccd1 _10112_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout98_A _07096_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09294__A _10479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10041_ _09887_/X _10026_/X _10028_/Y _09236_/Y _10040_/X vssd1 vssd1 vccd1 vccd1
+ _10041_/X sky130_fd_sc_hd__a221o_1
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07555__B1 _09922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ hold266/A _11992_/B vssd1 vssd1 vccd1 vccd1 _12068_/B sky130_fd_sc_hd__or2_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
X_10943_ _10943_/A _10943_/B vssd1 vssd1 vccd1 vccd1 _10947_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07858__A1 _09770_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07542__A _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12851__A1 _11779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11064__A _11582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11654__A2 _09257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07858__B2 _09940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10874_ _10874_/A _10874_/B _10874_/C vssd1 vssd1 vccd1 vccd1 _10875_/B sky130_fd_sc_hd__or3_1
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12613_ _12600_/Y _12621_/C _12623_/B vssd1 vssd1 vccd1 vccd1 _12614_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_38_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12544_ _12553_/A _12544_/B vssd1 vssd1 vccd1 vccd1 _12546_/C sky130_fd_sc_hd__nand2_1
XANTENNA__10614__B1 _10748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12475_ _12476_/A _12476_/B _12476_/C vssd1 vssd1 vccd1 vccd1 _12483_/B sky130_fd_sc_hd__a21o_1
X_11426_ _11426_/A _11426_/B vssd1 vssd1 vccd1 vccd1 _11429_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_6 instruction[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11357_ _11650_/B _11549_/C hold292/A vssd1 vssd1 vccd1 vccd1 _11359_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10308_ _10291_/A _12420_/A0 _10301_/Y _10302_/X _10307_/X vssd1 vssd1 vccd1 vccd1
+ _10308_/Y sky130_fd_sc_hd__o221ai_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11288_ _11288_/A _11288_/B vssd1 vssd1 vccd1 vccd1 _11289_/B sky130_fd_sc_hd__and2_1
X_13027_ _13162_/A hold230/X vssd1 vssd1 vccd1 vccd1 hold231/A sky130_fd_sc_hd__and2_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10239_ _07608_/A _07608_/B _10473_/B2 vssd1 vssd1 vccd1 vccd1 _10242_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_89_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10289__S _12054_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07450_ _10623_/A _07450_/B vssd1 vssd1 vccd1 vccd1 _07530_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07381_ _09667_/A _07381_/B vssd1 vssd1 vccd1 vccd1 _07384_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09120_ _10234_/A2 _07959_/B fanout29/X _10725_/A vssd1 vssd1 vccd1 vccd1 _09121_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09051_ _07554_/B _10337_/A _12823_/A1 _07175_/A vssd1 vssd1 vccd1 vccd1 _09052_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08002_ _08001_/A _08001_/B _08001_/C vssd1 vssd1 vccd1 vccd1 _08004_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_690 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07234__C1 _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout100_A _07088_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10384__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07785__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09953_ _10060_/A _09953_/B vssd1 vssd1 vccd1 vccd1 _09957_/A sky130_fd_sc_hd__xnor2_4
X_09884_ _09191_/X _09213_/X _10297_/S vssd1 vssd1 vccd1 vccd1 _09884_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08904_ _08904_/A _08904_/B vssd1 vssd1 vccd1 vccd1 _08906_/B sky130_fd_sc_hd__nor2_2
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ fanout53/X _10473_/B2 _10240_/A fanout51/X vssd1 vssd1 vccd1 vccd1 _08836_/B
+ sky130_fd_sc_hd__o22a_1
X_08766_ _08766_/A _08766_/B vssd1 vssd1 vccd1 vccd1 _11538_/C sky130_fd_sc_hd__xnor2_2
X_07717_ _07717_/A _07717_/B vssd1 vssd1 vccd1 vccd1 _07755_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07362__A _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08458__A _08502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12833__A1 _07195_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10500__B _12087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08697_ _08176_/Y _08180_/Y _08181_/X vssd1 vssd1 vccd1 vccd1 _08697_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_94_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07648_ _10623_/A _07648_/B vssd1 vssd1 vccd1 vccd1 _07652_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08501__A2 _10221_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07579_ _07580_/A _07580_/B vssd1 vssd1 vccd1 vccd1 _07581_/A sky130_fd_sc_hd__and2_1
X_09318_ _09667_/A _09318_/B vssd1 vssd1 vccd1 vccd1 _09319_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_106_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10590_ _12096_/A _10590_/B vssd1 vssd1 vccd1 vccd1 _10591_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_63_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06837__A_N _07233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09249_ _11138_/A _09250_/B vssd1 vssd1 vccd1 vccd1 _09249_/Y sky130_fd_sc_hd__nor2_1
X_12260_ reg1_val[27] curr_PC[27] vssd1 vssd1 vccd1 vccd1 _12260_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_50_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11050__C _11050_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11211_ _11212_/A _11212_/B vssd1 vssd1 vccd1 vccd1 _11211_/X sky130_fd_sc_hd__and2_1
XFILLER_0_105_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12191_ _06672_/D _12189_/X _12190_/Y vssd1 vssd1 vccd1 vccd1 _12215_/B sky130_fd_sc_hd__o21a_1
X_11142_ _11820_/A _11137_/X _11141_/Y _12446_/C1 vssd1 vssd1 vccd1 vccd1 _11157_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11073_ _11764_/A _07417_/B fanout41/X _11592_/A vssd1 vssd1 vccd1 vccd1 _11074_/B
+ sky130_fd_sc_hd__a22o_1
X_10024_ _11138_/A _10024_/B vssd1 vssd1 vccd1 vccd1 _10024_/X sky130_fd_sc_hd__or2_1
XANTENNA__13077__A1 _11582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11975_ _11809_/A _08784_/Y _08786_/Y vssd1 vssd1 vccd1 vccd1 _11977_/A sky130_fd_sc_hd__a21oi_1
X_10926_ hold285/A _12449_/B1 _11035_/B _12376_/C1 vssd1 vssd1 vccd1 vccd1 _10926_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_0_85_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10857_ _10858_/A _10858_/B vssd1 vssd1 vccd1 vccd1 _10980_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_27_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13213__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ _10788_/A _10788_/B vssd1 vssd1 vccd1 vccd1 _10788_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_6_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08256__A1 _08540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08256__B2 _08515_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12527_ reg1_val[10] curr_PC[10] _12638_/S vssd1 vssd1 vccd1 vccd1 _12529_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_42_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12458_ _07147_/B _09257_/S _06958_/A vssd1 vssd1 vccd1 vccd1 _12458_/X sky130_fd_sc_hd__o21a_1
X_11409_ _11409_/A _11409_/B vssd1 vssd1 vccd1 vccd1 _11410_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09756__A1 _09225_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08559__A2 _09770_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12389_ _12389_/A _12389_/B vssd1 vssd1 vccd1 vccd1 _12390_/B sky130_fd_sc_hd__or2_1
XANTENNA__11563__A1 _10788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07447__A _09667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06950_ _09226_/B _09237_/B vssd1 vssd1 vccd1 vccd1 _09222_/B sky130_fd_sc_hd__nor2_2
XANTENNA__07519__B1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06881_ _06963_/B _06878_/Y _06879_/X _06880_/Y vssd1 vssd1 vccd1 vccd1 _06881_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12499__S _12520_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09662__A _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_10_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08620_ _08630_/A _08625_/B vssd1 vssd1 vccd1 vccd1 _08620_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12815__A1 _07166_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08551_ _08739_/A _08741_/A vssd1 vssd1 vccd1 vccd1 _08681_/A sky130_fd_sc_hd__and2_1
XFILLER_0_76_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08482_ _08483_/B _08483_/A vssd1 vssd1 vccd1 vccd1 _08482_/Y sky130_fd_sc_hd__nand2b_1
X_07502_ _07502_/A _07502_/B vssd1 vssd1 vccd1 vccd1 _07503_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_92_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07433_ _07433_/A _07433_/B vssd1 vssd1 vccd1 vccd1 _07440_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__12528__A _12689_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout148_A _07068_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09103_ _09103_/A _11497_/A vssd1 vssd1 vccd1 vccd1 _09109_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08247__A1 _08649_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08247__B2 _08657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07364_ _07363_/A _07363_/B _07588_/A vssd1 vssd1 vccd1 vccd1 _07365_/B sky130_fd_sc_hd__o21bai_1
XFILLER_0_127_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10054__A1 _07282_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07295_ reg1_val[10] _07295_/B vssd1 vssd1 vccd1 vccd1 _07297_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08798__A2 _08799_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09034_ _09034_/A _09034_/B vssd1 vssd1 vccd1 vccd1 _09708_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__07470__A2 _10337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10357__A2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07758__B1 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11306__A1 _11476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10109__A2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09936_ _09936_/A _09936_/B vssd1 vssd1 vccd1 vccd1 _09938_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11306__B2 _11406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09867_ _09868_/B _09868_/C _10331_/A vssd1 vssd1 vccd1 vccd1 _09869_/A sky130_fd_sc_hd__a21oi_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09798_ _09799_/A _09799_/B vssd1 vssd1 vccd1 vccd1 _09800_/A sky130_fd_sc_hd__or2_1
X_08818_ _07134_/Y _07417_/B fanout42/X _07166_/Y vssd1 vssd1 vccd1 vccd1 _08819_/B
+ sky130_fd_sc_hd__a22o_1
X_08749_ _08749_/A _08757_/B _08749_/C vssd1 vssd1 vccd1 vccd1 _08751_/C sky130_fd_sc_hd__and3_1
X_11760_ _11761_/B _11760_/B vssd1 vssd1 vccd1 vccd1 _11762_/A sky130_fd_sc_hd__nand2b_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ fanout62/X fanout47/X fanout45/X _11671_/A vssd1 vssd1 vccd1 vccd1 _10712_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_67_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11691_ _11692_/A _11692_/B _11692_/C vssd1 vssd1 vccd1 vccd1 _11785_/A sky130_fd_sc_hd__a21oi_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10832__A3 fanout8/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12438__A _12438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10642_ _10634_/B _10499_/B _10516_/B _10515_/B _10515_/A vssd1 vssd1 vccd1 vccd1
+ _10643_/B sky130_fd_sc_hd__a32o_1
XANTENNA__08238__B2 _09404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08238__A1 _08649_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10573_ _06763_/Y _10568_/Y _10570_/Y _10571_/X _10572_/X vssd1 vssd1 vccd1 vccd1
+ _10573_/X sky130_fd_sc_hd__o221a_1
X_13361_ _13365_/CLK _13361_/D vssd1 vssd1 vccd1 vccd1 hold245/A sky130_fd_sc_hd__dfxtp_2
XFILLER_0_36_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13292_ _13390_/CLK _13292_/D vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12312_ _06885_/Y _12311_/Y _12404_/S vssd1 vssd1 vccd1 vccd1 _12313_/B sky130_fd_sc_hd__mux2_1
XANTENNA__12990__B1 _13257_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12243_ _12243_/A _12243_/B _12243_/C vssd1 vssd1 vccd1 vccd1 _12244_/B sky130_fd_sc_hd__or3_1
XFILLER_0_51_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12174_ _12175_/B _12175_/A vssd1 vssd1 vccd1 vccd1 _12243_/B sky130_fd_sc_hd__and2b_1
XANTENNA__07267__A _09794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11125_ _11052_/X _11124_/Y _09150_/X vssd1 vssd1 vccd1 vccd1 _11125_/Y sky130_fd_sc_hd__a21oi_1
X_11056_ _10623_/A _10950_/B _10953_/X vssd1 vssd1 vccd1 vccd1 _11058_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__09482__A _09944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13208__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10007_ _09910_/Y _10324_/A _12356_/B1 vssd1 vssd1 vccd1 vccd1 _10007_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_max_cap113_A _10225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10808__A0 _12420_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08477__A1 _08598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11958_ _11959_/A _11959_/B vssd1 vssd1 vccd1 vccd1 _12040_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12273__A2 _11829_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08477__B2 _08538_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11481__B1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11889_ _11124_/B _11528_/Y _11886_/Y _11888_/Y vssd1 vssd1 vccd1 vccd1 _11890_/B
+ sky130_fd_sc_hd__o31ai_4
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10909_ _06753_/Y _10791_/B _10808_/S vssd1 vssd1 vccd1 vccd1 _10909_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09426__B1 _09257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07080_ _07080_/A _07080_/B vssd1 vssd1 vccd1 vccd1 _11592_/A sky130_fd_sc_hd__nand2_8
XANTENNA__09657__A _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12083__A _12087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07177__A _09922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout107 _07298_/Y vssd1 vssd1 vccd1 vccd1 _08484_/B sky130_fd_sc_hd__buf_8
X_07982_ _07080_/A _07080_/B _06993_/A vssd1 vssd1 vccd1 vccd1 _07985_/B sky130_fd_sc_hd__a21o_1
Xfanout129 _07120_/X vssd1 vssd1 vccd1 vccd1 _08561_/A2 sky130_fd_sc_hd__buf_6
XFILLER_0_10_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06933_ instruction[16] _06933_/B vssd1 vssd1 vccd1 vccd1 dest_idx[5] sky130_fd_sc_hd__and2_4
X_09721_ _09387_/X _09389_/X _09727_/S vssd1 vssd1 vccd1 vccd1 _09721_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07905__A _08334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06864_ _06701_/Y _06856_/Y _06863_/Y vssd1 vssd1 vccd1 vccd1 _06864_/Y sky130_fd_sc_hd__o21ai_2
X_09652_ _09944_/A _09652_/B _09652_/C vssd1 vssd1 vccd1 vccd1 _09653_/C sky130_fd_sc_hd__nand3_1
X_06795_ reg1_val[4] _07117_/C vssd1 vssd1 vccd1 vccd1 _06796_/B sky130_fd_sc_hd__nand2_1
X_09583_ _12322_/A1 _09582_/X hold237/A vssd1 vssd1 vccd1 vccd1 _09583_/Y sky130_fd_sc_hd__a21oi_1
X_08603_ _08603_/A _08603_/B _08610_/A _08603_/D vssd1 vssd1 vccd1 vccd1 _08603_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_89_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout265_A _12796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08534_ _08575_/A _08534_/B vssd1 vssd1 vccd1 vccd1 _08557_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_49_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08465_ _08465_/A _08465_/B vssd1 vssd1 vccd1 vccd1 _08491_/B sky130_fd_sc_hd__xor2_2
XANTENNA__12016__A2 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09417__B1 _12205_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08396_ _08421_/A _08394_/B _08437_/A vssd1 vssd1 vccd1 vccd1 _08406_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07416_ _09834_/A _07416_/B vssd1 vssd1 vccd1 vccd1 _07420_/A sky130_fd_sc_hd__xor2_1
XANTENNA__09968__A1 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09968__B2 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07347_ _09834_/A _07347_/B vssd1 vssd1 vccd1 vccd1 _07349_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07979__B1 _08457_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07278_ _07278_/A _07278_/B vssd1 vssd1 vccd1 vccd1 _07279_/B sky130_fd_sc_hd__and2_1
X_09017_ _09017_/A _09017_/B vssd1 vssd1 vccd1 vccd1 _09018_/B sky130_fd_sc_hd__and2_2
XFILLER_0_21_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10506__A _11398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06703__B _12660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09422__C_N _12644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold161 hold161/A vssd1 vssd1 vccd1 vccd1 hold161/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold150 hold158/X vssd1 vssd1 vccd1 vccd1 hold150/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 hold172/A vssd1 vssd1 vccd1 vccd1 hold172/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 hold183/A vssd1 vssd1 vccd1 vccd1 hold183/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 hold194/A vssd1 vssd1 vccd1 vccd1 hold194/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10225__B _11946_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout80_A _11198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09919_ _09919_/A _09919_/B vssd1 vssd1 vccd1 vccd1 _09920_/B sky130_fd_sc_hd__nor2_1
X_12930_ hold85/X hold279/X vssd1 vssd1 vccd1 vccd1 _13153_/B sky130_fd_sc_hd__nand2b_1
X_12861_ _12169_/A _12863_/A2 hold45/X _13249_/A vssd1 vssd1 vccd1 vccd1 _13291_/D
+ sky130_fd_sc_hd__o211a_1
X_11812_ _11726_/A _11724_/Y _11742_/A vssd1 vssd1 vccd1 vccd1 _11812_/X sky130_fd_sc_hd__a21bo_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12792_ _12786_/A _12788_/B _12786_/B vssd1 vssd1 vccd1 vccd1 _12793_/B sky130_fd_sc_hd__a21bo_2
XANTENNA__09656__B1 _10245_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _11742_/A _09422_/B _11742_/Y _12421_/A1 vssd1 vssd1 vccd1 vccd1 _11743_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09120__A2 _07959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11674_ _11674_/A _11674_/B vssd1 vssd1 vccd1 vccd1 _11675_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11072__A _12093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10625_ _11381_/A _10625_/B vssd1 vssd1 vccd1 vccd1 _10627_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10556_ _06896_/C _10554_/X _10555_/Y vssd1 vssd1 vccd1 vccd1 _10556_/X sky130_fd_sc_hd__o21a_1
X_13344_ _13396_/CLK _13344_/D vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13275_ _13296_/CLK _13275_/D vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__dfxtp_1
X_10487_ _10487_/A _10487_/B vssd1 vssd1 vccd1 vccd1 _10517_/B sky130_fd_sc_hd__and2_1
XANTENNA__10416__A _10416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12226_ fanout15/X fanout12/X fanout8/A fanout23/X vssd1 vssd1 vccd1 vccd1 _12227_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12157_ _12157_/A _12157_/B vssd1 vssd1 vccd1 vccd1 _12160_/B sky130_fd_sc_hd__xnor2_1
X_11108_ _11108_/A _11108_/B vssd1 vssd1 vccd1 vccd1 _11109_/B sky130_fd_sc_hd__and2_1
X_12088_ _12088_/A _12088_/B vssd1 vssd1 vccd1 vccd1 _12105_/A sky130_fd_sc_hd__xnor2_1
X_11039_ _12420_/A0 _09422_/B _11039_/S vssd1 vssd1 vccd1 vccd1 _11039_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06580_ instruction[5] vssd1 vssd1 vccd1 vccd1 _09234_/B sky130_fd_sc_hd__clkinv_4
XANTENNA__09647__B1 _10240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07460__A _09944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10297__S _10297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08250_ _08315_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08250_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_117_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07201_ _11381_/A _07192_/B _07200_/X vssd1 vssd1 vccd1 vccd1 _07201_/X sky130_fd_sc_hd__o21a_2
X_08181_ _08182_/A _08182_/B vssd1 vssd1 vccd1 vccd1 _08181_/X sky130_fd_sc_hd__and2b_1
X_07132_ _07215_/B _07133_/A _07117_/C vssd1 vssd1 vccd1 vccd1 _08613_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_54_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07063_ reg1_val[7] _07063_/B vssd1 vssd1 vccd1 vccd1 _07063_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07965_ _08061_/B _07965_/B vssd1 vssd1 vccd1 vccd1 _08062_/A sky130_fd_sc_hd__and2b_1
XANTENNA__08138__B1 _08457_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06916_ instruction[6] _09234_/B vssd1 vssd1 vccd1 vccd1 _09239_/B sky130_fd_sc_hd__nand2_8
X_09704_ _09704_/A _09704_/B vssd1 vssd1 vccd1 vccd1 _09707_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_4_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11142__C1 _12446_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09635_ _09636_/A _09636_/B vssd1 vssd1 vccd1 vccd1 _09850_/A sky130_fd_sc_hd__nand2b_1
X_07896_ _07896_/A _07896_/B vssd1 vssd1 vccd1 vccd1 _07897_/B sky130_fd_sc_hd__nor2_1
X_06847_ _07262_/A _11242_/A vssd1 vssd1 vccd1 vccd1 _06847_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_78_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06778_ reg1_val[6] _07283_/A vssd1 vssd1 vccd1 vccd1 _06781_/A sky130_fd_sc_hd__or2_1
X_09566_ _09174_/X _09178_/X _09727_/S vssd1 vssd1 vccd1 vccd1 _09566_/X sky130_fd_sc_hd__mux2_1
X_09497_ _09667_/A _09497_/B vssd1 vssd1 vccd1 vccd1 _09498_/B sky130_fd_sc_hd__xnor2_1
X_08517_ _08552_/A _08552_/B vssd1 vssd1 vccd1 vccd1 _08553_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_108_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08448_ _08471_/A _08471_/B _08444_/X vssd1 vssd1 vccd1 vccd1 _08462_/A sky130_fd_sc_hd__o21a_1
XANTENNA__08861__B2 _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10410_ _10411_/A _10411_/B vssd1 vssd1 vccd1 vccd1 _10538_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11748__B2 _12365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08379_ _10748_/A _08379_/B vssd1 vssd1 vccd1 vccd1 _08384_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11390_ _11946_/B _07157_/Y fanout42/X _07013_/X vssd1 vssd1 vccd1 vccd1 _11391_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10341_ _10341_/A _10341_/B vssd1 vssd1 vccd1 vccd1 _10343_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10272_ _10272_/A _10272_/B vssd1 vssd1 vccd1 vccd1 _10274_/B sky130_fd_sc_hd__xnor2_4
X_13060_ hold98/X _13094_/A2 _13101_/A2 hold82/X _13259_/A vssd1 vssd1 vccd1 vccd1
+ hold99/A sky130_fd_sc_hd__o221a_1
X_12011_ _12012_/A _12012_/B _12012_/C vssd1 vssd1 vccd1 vccd1 _12013_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__11920__A1 _09149_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09877__B1 _11637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12913_ _13106_/A _13106_/B _12910_/X vssd1 vssd1 vccd1 vccd1 _13111_/A sky130_fd_sc_hd__a21o_1
X_12844_ hold121/X _12862_/B vssd1 vssd1 vccd1 vccd1 hold122/A sky130_fd_sc_hd__or2_1
XFILLER_0_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10239__A1 _07608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12775_ _12775_/A _12780_/C vssd1 vssd1 vccd1 vccd1 loadstore_address[27] sky130_fd_sc_hd__xnor2_4
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11726_ _11726_/A _11726_/B vssd1 vssd1 vccd1 vccd1 _11726_/Y sky130_fd_sc_hd__nand2_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11657_ _11656_/X _11657_/B _11657_/C _11657_/D vssd1 vssd1 vccd1 vccd1 _11657_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_83_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11588_ fanout62/X fanout10/X fanout5/X _11671_/A vssd1 vssd1 vccd1 vccd1 _11589_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_107_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10608_ _11770_/A _10608_/B vssd1 vssd1 vccd1 vccd1 _10609_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09801__B1 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13327_ _13392_/CLK hold234/X vssd1 vssd1 vccd1 vccd1 hold232/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10539_ _10539_/A _10658_/A vssd1 vssd1 vccd1 vccd1 _10779_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_3_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13258_ hold127/X hold298/A hold305/A hold66/X vssd1 vssd1 vccd1 vccd1 hold128/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08368__B1 _10338_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13189_ _13189_/A _13189_/B vssd1 vssd1 vccd1 vccd1 _13189_/Y sky130_fd_sc_hd__xnor2_1
X_12209_ _07046_/B _09257_/S _12208_/X vssd1 vssd1 vccd1 vccd1 _12209_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__06918__A1 _06783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07455__A _10479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07750_ _07750_/A _07750_/B vssd1 vssd1 vccd1 vccd1 _07810_/A sky130_fd_sc_hd__xnor2_1
X_06701_ _06701_/A vssd1 vssd1 vccd1 vccd1 _06701_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09670__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07681_ _07681_/A _07681_/B vssd1 vssd1 vccd1 vccd1 _07743_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06632_ _06630_/X _06632_/B vssd1 vssd1 vccd1 vccd1 _12313_/A sky130_fd_sc_hd__and2b_1
X_09420_ _09418_/Y _09419_/Y _11637_/A vssd1 vssd1 vccd1 vccd1 _09420_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07190__A _09667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09351_ _09351_/A _09351_/B vssd1 vssd1 vccd1 vccd1 _09352_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_59_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08302_ _08561_/B1 _08484_/B _09479_/B1 _08576_/A2 vssd1 vssd1 vccd1 vccd1 _08303_/B
+ sky130_fd_sc_hd__o22a_1
X_09282_ _09122_/A _09122_/B _09118_/X vssd1 vssd1 vccd1 vccd1 _09284_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08233_ _08234_/A _08234_/B vssd1 vssd1 vccd1 vccd1 _08233_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12536__A _12696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07110__A4 _12740_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08164_ _08162_/A _08162_/B _08163_/Y vssd1 vssd1 vccd1 vccd1 _08227_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_125_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07115_ reg1_val[23] _07210_/B _07115_/C vssd1 vssd1 vccd1 vccd1 _07168_/B sky130_fd_sc_hd__or3_1
XFILLER_0_42_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08095_ _08095_/A _08095_/B vssd1 vssd1 vccd1 vccd1 _08098_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_15_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07046_ _07049_/A _07046_/B _07046_/C vssd1 vssd1 vccd1 vccd1 _07048_/C sky130_fd_sc_hd__nand3_2
XFILLER_0_113_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13104__B1 _13254_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07582__A1 _07198_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07582__B2 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ _08997_/A _08997_/B vssd1 vssd1 vccd1 vccd1 _08998_/B sky130_fd_sc_hd__xor2_4
XANTENNA__12458__A2 _09257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07948_ _07948_/A _07948_/B _07948_/C vssd1 vssd1 vccd1 vccd1 _07948_/X sky130_fd_sc_hd__and3_1
X_07879_ _07879_/A _07879_/B vssd1 vssd1 vccd1 vccd1 _07944_/A sky130_fd_sc_hd__nor2_1
X_10890_ _10890_/A _10890_/B vssd1 vssd1 vccd1 vccd1 _10892_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout43_A _07417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09618_ _09617_/B _09618_/B vssd1 vssd1 vccd1 vccd1 _09619_/B sky130_fd_sc_hd__and2b_1
X_09549_ _09549_/A _09708_/A _09863_/A _10004_/A vssd1 vssd1 vccd1 vccd1 _10138_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12560_ _12560_/A _12560_/B _12560_/C vssd1 vssd1 vccd1 vccd1 _12561_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_26_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11511_ _11511_/A _11511_/B vssd1 vssd1 vccd1 vccd1 _11514_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_108_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12491_ _12497_/B _12491_/B vssd1 vssd1 vccd1 vccd1 new_PC[4] sky130_fd_sc_hd__and2_4
XFILLER_0_81_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11442_ _11377_/Y _11840_/C _12356_/B1 vssd1 vssd1 vccd1 vccd1 _11442_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11373_ _12471_/S _11370_/X _11371_/Y _11372_/X vssd1 vssd1 vccd1 vccd1 dest_val[16]
+ sky130_fd_sc_hd__a22o_4
XANTENNA__10944__A2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13112_ hold235/X _13111_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13112_/X sky130_fd_sc_hd__mux2_1
X_10324_ _10324_/A _10324_/B _10324_/C _10324_/D vssd1 vssd1 vccd1 vccd1 _10581_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_34_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12146__A1 _12379_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10255_ _10255_/A _10255_/B _10255_/C vssd1 vssd1 vccd1 vccd1 _10257_/B sky130_fd_sc_hd__or3_1
X_13043_ _07029_/B _12820_/B hold166/X vssd1 vssd1 vccd1 vccd1 _13331_/D sky130_fd_sc_hd__a21boi_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10186_ _10448_/C _10185_/Y _10183_/X vssd1 vssd1 vccd1 vccd1 dest_val[6] sky130_fd_sc_hd__o21ai_4
Xfanout290 reg1_val[15] vssd1 vssd1 vccd1 vccd1 _11242_/A sky130_fd_sc_hd__buf_6
XANTENNA__09490__A _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_15_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06619__A _06723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12827_ _07238_/Y _13101_/B2 hold33/X _13147_/A vssd1 vssd1 vccd1 vccd1 _13274_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12082__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12758_ reg1_val[24] _12790_/B vssd1 vssd1 vccd1 vccd1 _12759_/B sky130_fd_sc_hd__or2_1
X_11709_ _11709_/A _11709_/B vssd1 vssd1 vccd1 vccd1 _11710_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_126_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12689_ reg1_val[10] _12689_/B vssd1 vssd1 vccd1 vccd1 _12690_/B sky130_fd_sc_hd__or2_1
XFILLER_0_126_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12803__B _12803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10604__A _11284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12091__A _12157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10148__B1 _09150_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08920_ _09037_/A _08920_/B vssd1 vssd1 vccd1 vccd1 _08920_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06801__B _07165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08851_ fanout84/X fanout78/X fanout74/X fanout80/X vssd1 vssd1 vccd1 vccd1 _08852_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11360__A2 _12420_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07802_ _07802_/A _07802_/B vssd1 vssd1 vccd1 vccd1 _07822_/B sky130_fd_sc_hd__xnor2_2
X_08782_ _08791_/A _08781_/C _08790_/B vssd1 vssd1 vccd1 vccd1 _08783_/B sky130_fd_sc_hd__a21o_1
X_07733_ _07743_/A _07743_/B vssd1 vssd1 vccd1 vccd1 _07733_/X sky130_fd_sc_hd__or2_1
XANTENNA_fanout178_A _12379_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08513__B1 _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07664_ _07366_/A _07366_/B _07355_/X vssd1 vssd1 vccd1 vccd1 _07666_/B sky130_fd_sc_hd__a21oi_2
X_06615_ instruction[41] _06927_/B _06612_/X vssd1 vssd1 vccd1 vccd1 _06703_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_94_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09403_ _09208_/X _09210_/X _09403_/S vssd1 vssd1 vccd1 vccd1 _09403_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07595_ _12224_/A _07361_/B _11844_/A vssd1 vssd1 vccd1 vccd1 _07596_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__12073__B1 _09221_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08816__B2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08816__A1 _07830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09334_ _09335_/A _09335_/B vssd1 vssd1 vccd1 vccd1 _09334_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_47_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08292__A2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09265_ _09934_/A _07362_/B fanout16/X _09822_/A vssd1 vssd1 vccd1 vccd1 _09266_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_62_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09196_ _09218_/A reg1_val[31] _09211_/S vssd1 vssd1 vccd1 vccd1 _09196_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08216_ _08216_/A _08216_/B vssd1 vssd1 vccd1 vccd1 _08222_/A sky130_fd_sc_hd__or2_1
XFILLER_0_28_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07079__B _07080_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08147_ _08334_/A _08147_/B vssd1 vssd1 vccd1 vccd1 _08150_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08044__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08078_ _08068_/A _08068_/C _08068_/B vssd1 vssd1 vccd1 vccd1 _08079_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_113_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07029_ _08502_/A _07029_/B vssd1 vssd1 vccd1 vccd1 _07031_/B sky130_fd_sc_hd__or2_1
XANTENNA__12713__B _12714_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10040_ _12444_/B _12446_/C1 _10039_/Y _10034_/Y vssd1 vssd1 vccd1 vccd1 _10040_/X
+ sky130_fd_sc_hd__a31o_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07555__A1 _07959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ hold201/A _12447_/B1 _12065_/B _12205_/B1 vssd1 vssd1 vccd1 vccd1 _11991_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_98_623 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
X_10942_ _10943_/A _10943_/B vssd1 vssd1 vccd1 vccd1 _11055_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12851__A2 _12863_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07858__A2 _08289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10873_ _10874_/A _10874_/B _10874_/C vssd1 vssd1 vccd1 vccd1 _10875_/A sky130_fd_sc_hd__o21ai_1
X_12612_ _12612_/A vssd1 vssd1 vccd1 vccd1 _12621_/C sky130_fd_sc_hd__inv_2
XFILLER_0_109_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12543_ _12702_/B _12543_/B vssd1 vssd1 vccd1 vccd1 _12544_/B sky130_fd_sc_hd__or2_1
XFILLER_0_81_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10614__A1 _10240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12474_ _12483_/A _12474_/B vssd1 vssd1 vccd1 vccd1 _12476_/C sky130_fd_sc_hd__nand2_1
X_11425_ _11426_/A _11426_/B vssd1 vssd1 vccd1 vccd1 _11524_/A sky130_fd_sc_hd__nand2_1
XANTENNA_7 instruction[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11356_ hold275/A _11356_/B vssd1 vssd1 vccd1 vccd1 _11549_/C sky130_fd_sc_hd__or2_1
XFILLER_0_22_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10307_ _06773_/Y _12144_/A1 _09422_/B _06775_/B _10306_/X vssd1 vssd1 vccd1 vccd1
+ _10307_/X sky130_fd_sc_hd__o221a_1
XANTENNA__08991__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11287_ _11288_/A _11288_/B vssd1 vssd1 vccd1 vccd1 _11387_/A sky130_fd_sc_hd__nor2_1
X_13026_ _13322_/Q _13171_/B2 _13209_/A2 hold229/X vssd1 vssd1 vccd1 vccd1 hold230/A
+ sky130_fd_sc_hd__a22o_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10238_ _10066_/A _10064_/Y _10063_/Y vssd1 vssd1 vccd1 vccd1 _10249_/A sky130_fd_sc_hd__a21o_1
XANTENNA__11342__A2 _11567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10169_ _10169_/A _10169_/B vssd1 vssd1 vccd1 vccd1 _10169_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10550__B1 _10581_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12827__C1 _13147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13095__A2 _13101_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10302__B1 _12205_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12055__B1 _11637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07380_ _10871_/A fanout78/X fanout74/X _07198_/Y vssd1 vssd1 vccd1 vccd1 _07381_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08564__A _08564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07482__B1 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09050_ _09053_/A vssd1 vssd1 vccd1 vccd1 _09050_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_60_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08001_ _08001_/A _08001_/B _08001_/C vssd1 vssd1 vccd1 vccd1 _08005_/A sky130_fd_sc_hd__and3_1
XFILLER_0_13_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09952_ fanout56/X _08484_/B _10240_/A _12233_/A vssd1 vssd1 vccd1 vccd1 _09953_/B
+ sky130_fd_sc_hd__o22a_2
XANTENNA__07785__B2 _08501_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07785__A1 _08457_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08903_ _07644_/A _07644_/B _07641_/X vssd1 vssd1 vccd1 vccd1 _08906_/A sky130_fd_sc_hd__a21o_2
X_09883_ _09881_/X _09882_/X _11246_/S vssd1 vssd1 vccd1 vccd1 _09883_/X sky130_fd_sc_hd__mux2_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ _08834_/A _08834_/B vssd1 vssd1 vccd1 vccd1 _08883_/A sky130_fd_sc_hd__xnor2_1
X_08765_ _08765_/A _08765_/B vssd1 vssd1 vccd1 vccd1 _08766_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11165__A _12087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07716_ _07717_/A _07717_/B vssd1 vssd1 vccd1 vccd1 _07716_/X sky130_fd_sc_hd__or2_1
XANTENNA__07362__B _07362_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12833__A2 _12863_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08696_ _08013_/A _08013_/B _08695_/X vssd1 vssd1 vccd1 vccd1 _08696_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07647_ fanout98/X fanout86/X fanout84/X fanout82/X vssd1 vssd1 vccd1 vccd1 _07648_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_94_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07578_ _09836_/A _07578_/B vssd1 vssd1 vccd1 vccd1 _07580_/B sky130_fd_sc_hd__xnor2_1
X_09317_ fanout51/X fanout78/X fanout74/X _09661_/B2 vssd1 vssd1 vccd1 vccd1 _09318_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12708__B _12708_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06706__B _07078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09248_ _09248_/A _09248_/B vssd1 vssd1 vccd1 vccd1 _11247_/B sky130_fd_sc_hd__and2_1
XFILLER_0_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13010__A2 _13171_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09179_ _11134_/A reg1_val[17] _09180_/S vssd1 vssd1 vccd1 vccd1 _09179_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11050__D _11050_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11210_ _11210_/A vssd1 vssd1 vccd1 vccd1 _11212_/B sky130_fd_sc_hd__inv_2
X_12190_ _06672_/D _12189_/X _11637_/A vssd1 vssd1 vccd1 vccd1 _12190_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11141_ _11820_/A _11141_/B vssd1 vssd1 vccd1 vccd1 _11141_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11072_ _12093_/A _11072_/B vssd1 vssd1 vccd1 vccd1 _11076_/A sky130_fd_sc_hd__xor2_1
X_10023_ _10297_/S _09396_/X _10022_/X vssd1 vssd1 vccd1 vccd1 _10023_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07553__A _09834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13077__A2 _13101_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11974_ _11973_/A _12049_/B _09150_/X vssd1 vssd1 vccd1 vccd1 _11974_/X sky130_fd_sc_hd__a21o_1
X_10925_ _12449_/B1 _11035_/B hold285/A vssd1 vssd1 vccd1 vccd1 _10925_/X sky130_fd_sc_hd__a21o_1
X_10856_ _11582_/A _10856_/B vssd1 vssd1 vccd1 vccd1 _10858_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10787_ _11630_/A _08735_/Y _08737_/Y vssd1 vssd1 vccd1 vccd1 _10788_/B sky130_fd_sc_hd__o21a_1
XANTENNA__08256__A2 _09770_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12526_ _12532_/B _12526_/B vssd1 vssd1 vccd1 vccd1 new_PC[9] sky130_fd_sc_hd__and2_4
XANTENNA__11260__A1 _12421_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12457_ _12442_/Y _12443_/X _12446_/X _12456_/X vssd1 vssd1 vccd1 vccd1 _12457_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_41_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11408_ _11409_/A _11409_/B vssd1 vssd1 vccd1 vccd1 _11408_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_112_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11012__A1 _10546_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12388_ _12389_/A _12389_/B vssd1 vssd1 vccd1 vccd1 _12390_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11339_ _11526_/A _11340_/B vssd1 vssd1 vccd1 vccd1 _11840_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_94_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07519__A1 _09669_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13009_ _13019_/A hold178/X vssd1 vssd1 vccd1 vccd1 hold179/A sky130_fd_sc_hd__and2_1
XFILLER_0_94_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06880_ _06902_/A _06864_/Y instruction[6] vssd1 vssd1 vccd1 vccd1 _06880_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07519__B2 _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12276__B1 _09886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12815__A2 _13101_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08550_ _08550_/A _08550_/B _08550_/C vssd1 vssd1 vccd1 vccd1 _08741_/A sky130_fd_sc_hd__or3_2
XFILLER_0_49_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07501_ _07501_/A _07501_/B vssd1 vssd1 vccd1 vccd1 _07502_/B sky130_fd_sc_hd__xor2_4
X_08481_ _08479_/Y _08511_/B _08476_/X vssd1 vssd1 vccd1 vccd1 _08483_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07432_ _07678_/A _07431_/B _07403_/Y vssd1 vssd1 vccd1 vccd1 _07505_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_85_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08247__A2 _10595_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07363_ _07363_/A _07363_/B _07588_/A vssd1 vssd1 vccd1 vccd1 _07589_/A sky130_fd_sc_hd__or3b_1
XFILLER_0_17_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09102_ _09102_/A _09102_/B vssd1 vssd1 vccd1 vccd1 _09111_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_127_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10054__A2 _11946_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07294_ reg1_val[8] reg1_val[9] _07105_/D _07248_/A vssd1 vssd1 vccd1 vccd1 _07295_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_45_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout210_A _06946_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09033_ _09034_/A _09034_/B vssd1 vssd1 vccd1 vccd1 _09552_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_5_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08955__B1 _10245_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07758__B2 _08538_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07758__A1 _08598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09935_ _10337_/A _07596_/A _07596_/B _07238_/Y _07360_/X vssd1 vssd1 vccd1 vccd1
+ _09936_/B sky130_fd_sc_hd__a32o_1
XFILLER_0_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11306__A2 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09866_ _10137_/A _09551_/X _10137_/B _09865_/X vssd1 vssd1 vccd1 vccd1 _09868_/C
+ sky130_fd_sc_hd__o31a_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08817_ _09834_/A _08817_/B vssd1 vssd1 vccd1 vccd1 _08821_/A sky130_fd_sc_hd__xnor2_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09797_ _09797_/A _09797_/B vssd1 vssd1 vccd1 vccd1 _09799_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13059__A2 _12826_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08748_ _08749_/A _08749_/C _08757_/B vssd1 vssd1 vccd1 vccd1 _08751_/B sky130_fd_sc_hd__a21oi_2
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10817__B2 _09242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10817__A1 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08679_ _08678_/A _08678_/B _08678_/C _08589_/Y _08588_/X vssd1 vssd1 vccd1 vccd1
+ _08681_/C sky130_fd_sc_hd__a311o_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _10882_/B _10710_/B vssd1 vssd1 vccd1 vccd1 _10742_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_67_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07694__B1 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11690_ _11593_/A _11593_/B _11590_/Y vssd1 vssd1 vccd1 vccd1 _11692_/C sky130_fd_sc_hd__o21a_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06717__A _06723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10641_ _10487_/A _10487_/B _10484_/Y vssd1 vssd1 vccd1 vccd1 _10643_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__09435__A1 _07172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08238__A2 _08289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10572_ _07238_/A _09257_/S _09234_/X _06765_/B _06958_/A vssd1 vssd1 vccd1 vccd1
+ _10572_/X sky130_fd_sc_hd__o221a_1
X_13360_ _13360_/CLK hold17/X vssd1 vssd1 vccd1 vccd1 hold302/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07446__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13291_ _13390_/CLK _13291_/D vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__dfxtp_1
X_12311_ _06874_/A _06672_/D _12188_/X _12310_/X vssd1 vssd1 vccd1 vccd1 _12311_/Y
+ sky130_fd_sc_hd__o31ai_2
XFILLER_0_121_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12242_ _12244_/A vssd1 vssd1 vccd1 vccd1 _12242_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07548__A _09341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12173_ _12243_/A _12173_/B vssd1 vssd1 vccd1 vccd1 _12175_/B sky130_fd_sc_hd__or2_1
XANTENNA__07267__B _07267_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11124_ _11333_/A _11124_/B vssd1 vssd1 vccd1 vccd1 _11124_/Y sky130_fd_sc_hd__xnor2_4
X_11055_ _11055_/A _11055_/B vssd1 vssd1 vccd1 vccd1 _11058_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10505__B1 _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10006_ _10542_/A _10006_/B vssd1 vssd1 vccd1 vccd1 _10324_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__08379__A _10748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11957_ _11957_/A _11957_/B vssd1 vssd1 vccd1 vccd1 _11959_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_98_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10808__A1 _09422_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11481__A1 _12169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10284__A2 _10581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10908_ _11809_/A _08744_/A _08744_/B _10788_/A _10907_/Y vssd1 vssd1 vccd1 vccd1
+ _10933_/B sky130_fd_sc_hd__a311oi_1
XANTENNA__07685__B1 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08477__A2 _08561_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11481__B2 _06998_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11888_ _11714_/X _12043_/A _11886_/A _11530_/X _11887_/Y vssd1 vssd1 vccd1 vccd1
+ _11888_/Y sky130_fd_sc_hd__a221oi_2
XANTENNA__06627__A _06723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10839_ _10944_/B2 fanout43/X fanout42/X _07097_/X vssd1 vssd1 vccd1 vccd1 _10840_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09426__B2 _09728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09426__A1 _12416_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08842__A _10479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12509_ _12518_/A _12509_/B vssd1 vssd1 vccd1 vccd1 _12511_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_54_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10744__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout119 _07194_/Y vssd1 vssd1 vccd1 vccd1 _10595_/A1 sky130_fd_sc_hd__buf_8
XANTENNA__09673__A _09673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout108 _07283_/X vssd1 vssd1 vccd1 vccd1 _09940_/B2 sky130_fd_sc_hd__buf_8
X_07981_ _08023_/A _08023_/B vssd1 vssd1 vccd1 vccd1 _07993_/B sky130_fd_sc_hd__or2_1
X_06932_ instruction[15] _06933_/B vssd1 vssd1 vccd1 vccd1 dest_idx[4] sky130_fd_sc_hd__and2_4
X_09720_ _09718_/X _09719_/X _10294_/S vssd1 vssd1 vccd1 vccd1 _09720_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08289__A _09404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06863_ reg1_val[23] _07036_/A _06862_/Y vssd1 vssd1 vccd1 vccd1 _06863_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09901__A2 _07117_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ _09652_/B _09652_/C _09944_/A vssd1 vssd1 vccd1 vccd1 _09653_/B sky130_fd_sc_hd__a21o_1
X_06794_ reg1_val[4] _07117_/C vssd1 vssd1 vccd1 vccd1 _06796_/A sky130_fd_sc_hd__or2_1
X_09582_ hold301/A hold293/A vssd1 vssd1 vccd1 vccd1 _09582_/X sky130_fd_sc_hd__or2_1
X_08602_ _12808_/A _08598_/B _08580_/A vssd1 vssd1 vccd1 vccd1 _08603_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__07921__A _10243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09114__B1 _10974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08533_ _08649_/A2 _08561_/A2 _09940_/B2 _08657_/B vssd1 vssd1 vccd1 vccd1 _08534_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08464_ _08464_/A _08464_/B vssd1 vssd1 vccd1 vccd1 _08491_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_92_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08395_ _08436_/A _08436_/B vssd1 vssd1 vccd1 vccd1 _08437_/A sky130_fd_sc_hd__or2_1
X_07415_ _07830_/B _09822_/A fanout46/X _08576_/A2 vssd1 vssd1 vccd1 vccd1 _07416_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09968__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07346_ _09934_/A fanout46/X _07283_/X _07830_/B vssd1 vssd1 vccd1 vccd1 _07347_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_73_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07979__A1 _08540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07979__B2 _08515_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07277_ _07278_/A _07278_/B vssd1 vssd1 vccd1 vccd1 _07626_/A sky130_fd_sc_hd__nor2_1
X_09016_ _09016_/A _09016_/B vssd1 vssd1 vccd1 vccd1 _09017_/B sky130_fd_sc_hd__or2_1
XFILLER_0_115_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_458 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold162 hold206/X vssd1 vssd1 vccd1 vccd1 hold162/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10735__B1 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold140 hold305/X vssd1 vssd1 vccd1 vccd1 hold140/X sky130_fd_sc_hd__clkbuf_2
Xhold151 hold151/A vssd1 vssd1 vccd1 vccd1 hold151/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08928__B1 _10500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold173 hold173/A vssd1 vssd1 vccd1 vccd1 hold173/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 hold184/A vssd1 vssd1 vccd1 vccd1 hold184/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 hold195/A vssd1 vssd1 vccd1 vccd1 hold195/X sky130_fd_sc_hd__dlygate4sd3_1
X_09918_ _09919_/A _09919_/B vssd1 vssd1 vccd1 vccd1 _09920_/A sky130_fd_sc_hd__and2_1
XFILLER_0_95_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout73_A _07273_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08199__A _09404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09849_ _09623_/A _09623_/B _09622_/A vssd1 vssd1 vccd1 vccd1 _09854_/A sky130_fd_sc_hd__a21o_1
X_12860_ hold44/X _12862_/B vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__or2_1
XFILLER_0_87_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11811_ _11726_/A _06856_/Y _06858_/Y vssd1 vssd1 vccd1 vccd1 _11811_/X sky130_fd_sc_hd__o21a_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09105__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _12789_/X _12791_/B vssd1 vssd1 vccd1 vccd1 _12793_/A sky130_fd_sc_hd__nand2b_2
XANTENNA__09656__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09656__B2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11742_ _11742_/A _11829_/B vssd1 vssd1 vccd1 vccd1 _11742_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_83_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11673_ _11674_/A _11674_/B vssd1 vssd1 vccd1 vccd1 _11675_/A sky130_fd_sc_hd__or2_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10624_ _12233_/A fanout36/X fanout34/X _12087_/A vssd1 vssd1 vccd1 vccd1 _10625_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_107_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13343_ _13358_/CLK _13343_/D vssd1 vssd1 vccd1 vccd1 hold152/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10555_ _06896_/C _10554_/X _11637_/A vssd1 vssd1 vccd1 vccd1 _10555_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08631__A2 _07148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10486_ _10487_/A _10487_/B vssd1 vssd1 vccd1 vccd1 _10517_/A sky130_fd_sc_hd__nor2_1
X_13274_ _13398_/CLK _13274_/D vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__dfxtp_1
X_12225_ _12284_/A _12225_/B vssd1 vssd1 vccd1 vccd1 _12230_/A sky130_fd_sc_hd__and2_1
XFILLER_0_32_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12156_ fanout15/X _12335_/A fanout12/X fanout23/X vssd1 vssd1 vccd1 vccd1 _12157_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09592__B1 _12416_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11107_ _11107_/A _11107_/B vssd1 vssd1 vccd1 vccd1 _11109_/A sky130_fd_sc_hd__xnor2_2
X_12087_ _12087_/A _12087_/B vssd1 vssd1 vccd1 vccd1 _12088_/B sky130_fd_sc_hd__nor2_1
X_11038_ _11038_/A _12422_/A vssd1 vssd1 vccd1 vccd1 _11038_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_91_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12359__A _12359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12989_ _13001_/A hold216/X vssd1 vssd1 vccd1 vccd1 _13304_/D sky130_fd_sc_hd__and2_1
XANTENNA__09647__A1 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09647__B2 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07200_ _10092_/A _09667_/A _07200_/C vssd1 vssd1 vccd1 vccd1 _07200_/X sky130_fd_sc_hd__or3_2
XFILLER_0_6_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08180_ _08182_/B _08182_/A vssd1 vssd1 vccd1 vccd1 _08180_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_125_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12806__B _12870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07131_ _07136_/B _11854_/A vssd1 vssd1 vccd1 vccd1 _07131_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07062_ reg1_val[6] _07083_/C _07083_/D _07248_/A vssd1 vssd1 vccd1 vccd1 _07063_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_30_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11390__B1 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07964_ _09341_/A _07964_/B vssd1 vssd1 vccd1 vccd1 _07965_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08138__A1 _08598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06915_ reg1_idx[2] reg1_idx[3] _06915_/C _06915_/D vssd1 vssd1 vccd1 vccd1 int_return
+ sky130_fd_sc_hd__and4_4
XANTENNA__13131__B2 _06577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09703_ _09703_/A _09703_/B vssd1 vssd1 vccd1 vccd1 _09704_/B sky130_fd_sc_hd__xor2_4
X_07895_ _07896_/A _07896_/B vssd1 vssd1 vccd1 vccd1 _07897_/A sky130_fd_sc_hd__and2_1
XFILLER_0_4_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08138__B2 _08538_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06846_ _11131_/A _06844_/Y _06845_/Y vssd1 vssd1 vccd1 vccd1 _06846_/X sky130_fd_sc_hd__o21a_1
X_09634_ _09478_/A _09477_/B _09475_/X vssd1 vssd1 vccd1 vccd1 _09636_/B sky130_fd_sc_hd__a21o_1
X_06777_ _06815_/A _06817_/B1 _12675_/B _06776_/X vssd1 vssd1 vccd1 vccd1 _07283_/A
+ sky130_fd_sc_hd__a31o_4
X_09565_ _09563_/X _09564_/X _10294_/S vssd1 vssd1 vccd1 vccd1 _09565_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_93_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09496_ fanout53/X fanout78/X fanout74/X fanout51/X vssd1 vssd1 vccd1 vccd1 _09497_/B
+ sky130_fd_sc_hd__o22a_1
X_08516_ _08564_/A _08516_/B vssd1 vssd1 vccd1 vccd1 _08552_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07649__B1 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11996__A2 _09228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08447_ _08447_/A _08447_/B vssd1 vssd1 vccd1 vccd1 _08471_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08861__A2 _07608_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08378_ _08576_/A2 _10473_/B2 _09479_/B1 _07172_/Y vssd1 vssd1 vccd1 vccd1 _08379_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_45_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07329_ _10479_/A _07329_/B vssd1 vssd1 vccd1 vccd1 _07387_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10340_ _10341_/A _10341_/B vssd1 vssd1 vccd1 vccd1 _10468_/A sky130_fd_sc_hd__or2_1
XFILLER_0_21_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10271_ _10272_/B _10272_/A vssd1 vssd1 vccd1 vccd1 _10413_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12010_ _12084_/B _12010_/B vssd1 vssd1 vccd1 vccd1 _12012_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__13122__B2 _06577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07037__S _09673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09326__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12912_ hold16/X hold11/X vssd1 vssd1 vccd1 vccd1 _13106_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_69_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08657__A _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12843_ _07097_/X _12863_/A2 hold88/X _13210_/A vssd1 vssd1 vccd1 vccd1 _13282_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10239__A2 _07608_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12774_ reg1_val[27] _12790_/B vssd1 vssd1 vccd1 vccd1 _12780_/C sky130_fd_sc_hd__xnor2_4
X_11725_ _06856_/Y _11724_/Y _11813_/S vssd1 vssd1 vccd1 vccd1 _11726_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_96_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11656_ _09238_/Y _11650_/Y _11651_/X _11655_/X vssd1 vssd1 vccd1 vccd1 _11656_/X
+ sky130_fd_sc_hd__a31o_1
Xfanout90 _09922_/A vssd1 vssd1 vccd1 vccd1 _12093_/A sky130_fd_sc_hd__buf_8
XFILLER_0_52_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11587_ _11692_/B _11587_/B vssd1 vssd1 vccd1 vccd1 _11594_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10607_ _07013_/X fanout32/X fanout30/X _11779_/A vssd1 vssd1 vccd1 vccd1 _10608_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09801__B2 _11406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09801__A1 _11476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13326_ _13392_/CLK _13326_/D vssd1 vssd1 vccd1 vccd1 hold241/A sky130_fd_sc_hd__dfxtp_1
X_10538_ _10538_/A _10538_/B _10538_/C vssd1 vssd1 vccd1 vccd1 _10658_/A sky130_fd_sc_hd__or3_2
XFILLER_0_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13257_ hold66/X _13257_/A2 _12800_/Y _12804_/A vssd1 vssd1 vccd1 vccd1 _13259_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12208_ _12421_/A1 _12207_/X _06671_/B vssd1 vssd1 vccd1 vccd1 _12208_/X sky130_fd_sc_hd__a21o_1
X_10469_ _10645_/A _10469_/B vssd1 vssd1 vccd1 vccd1 _10471_/B sky130_fd_sc_hd__or2_1
XANTENNA__12642__A _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08368__A1 _06992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08368__B2 _08613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13188_ _12888_/X _13188_/B vssd1 vssd1 vccd1 vccd1 _13189_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_86_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11372__B1 _11752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12139_ _12139_/A _12139_/B vssd1 vssd1 vccd1 vccd1 _12139_/X sky130_fd_sc_hd__or2_1
XANTENNA__09951__A _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13113__B2 _06577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09317__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06700_ _06700_/A _06860_/A _11726_/A _11814_/A vssd1 vssd1 vccd1 vccd1 _06701_/A
+ sky130_fd_sc_hd__nor4_1
XFILLER_0_126_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07680_ _07745_/A _07745_/B vssd1 vssd1 vccd1 vccd1 _07680_/X sky130_fd_sc_hd__and2_1
XANTENNA__07471__A _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06631_ reg1_val[28] _08973_/B vssd1 vssd1 vccd1 vccd1 _06632_/B sky130_fd_sc_hd__or2_1
XFILLER_0_35_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09350_ _09350_/A _09350_/B vssd1 vssd1 vccd1 vccd1 _09351_/B sky130_fd_sc_hd__xor2_1
X_08301_ _08311_/A _08311_/B vssd1 vssd1 vccd1 vccd1 _08301_/Y sky130_fd_sc_hd__nor2_1
X_09281_ _09084_/X _09281_/B vssd1 vssd1 vccd1 vccd1 _09286_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_51_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08232_ _08232_/A _08232_/B vssd1 vssd1 vccd1 vccd1 _08234_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_90_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10938__B1 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10337__A _10337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08163_ _08186_/A _08186_/B vssd1 vssd1 vccd1 vccd1 _08163_/Y sky130_fd_sc_hd__nand2b_1
X_07114_ _07210_/B _07115_/C reg1_val[23] vssd1 vssd1 vccd1 vccd1 _07168_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08094_ _08094_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08095_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_113_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07045_ _07046_/B _06987_/A _06987_/B _07046_/C _07049_/A vssd1 vssd1 vccd1 vccd1
+ _07045_/X sky130_fd_sc_hd__a41o_1
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08996_ _08997_/A _08997_/B vssd1 vssd1 vccd1 vccd1 _08996_/X sky130_fd_sc_hd__and2b_1
XANTENNA__13104__A1 _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07582__A2 _08112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07947_ _07947_/A _07947_/B vssd1 vssd1 vccd1 vccd1 _07948_/C sky130_fd_sc_hd__nand2_1
XANTENNA__11666__A1 _11584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07381__A _09667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07878_ _07878_/A _07878_/B vssd1 vssd1 vccd1 vccd1 _07879_/B sky130_fd_sc_hd__and2_1
X_06829_ _07283_/A reg1_val[6] vssd1 vssd1 vccd1 vccd1 _06829_/Y sky130_fd_sc_hd__nand2b_1
X_09617_ _09618_/B _09617_/B vssd1 vssd1 vccd1 vccd1 _09619_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_78_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09548_ _09548_/A _09548_/B vssd1 vssd1 vccd1 vccd1 _10137_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_38_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout36_A _07192_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11510_ _11510_/A _11510_/B vssd1 vssd1 vccd1 vccd1 _11511_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_65_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09479_ fanout59/X _10473_/B2 _09479_/B1 fanout57/X vssd1 vssd1 vccd1 vccd1 _09480_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_93_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12490_ _12490_/A _12490_/B _12490_/C vssd1 vssd1 vccd1 vccd1 _12491_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_81_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11441_ _11840_/C vssd1 vssd1 vccd1 vccd1 _11567_/C sky130_fd_sc_hd__inv_2
XFILLER_0_33_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09795__B1 _10245_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11372_ curr_PC[16] _11375_/C _11752_/S vssd1 vssd1 vccd1 vccd1 _11372_/X sky130_fd_sc_hd__o21a_1
X_13111_ _13111_/A _13111_/B vssd1 vssd1 vccd1 vccd1 _13111_/Y sky130_fd_sc_hd__xnor2_1
X_10323_ _10146_/A _10146_/B _09715_/B vssd1 vssd1 vccd1 vccd1 _10324_/D sky130_fd_sc_hd__a21boi_1
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12146__A2 _10165_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12462__A _12642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10254_ _10383_/B _10253_/C _10253_/A vssd1 vssd1 vccd1 vccd1 _10255_/C sky130_fd_sc_hd__a21oi_1
X_13042_ hold125/X _13094_/A2 _13101_/A2 hold165/X _13039_/A vssd1 vssd1 vccd1 vccd1
+ hold166/A sky130_fd_sc_hd__o221a_1
XFILLER_0_100_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10185_ curr_PC[6] _10184_/B _11752_/S vssd1 vssd1 vccd1 vccd1 _10185_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__09771__A _09936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout280 _13259_/A vssd1 vssd1 vccd1 vccd1 _13039_/A sky130_fd_sc_hd__buf_4
Xfanout291 reg1_val[14] vssd1 vssd1 vccd1 vccd1 _11134_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__06619__B _12714_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12826_ hold32/X _12826_/B vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__or2_1
XFILLER_0_29_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12082__A1 _12233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12082__B2 _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10093__B1 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ reg1_val[24] _12790_/B vssd1 vssd1 vccd1 vccd1 _12764_/A sky130_fd_sc_hd__nand2_1
X_11708_ _11709_/A _11709_/B vssd1 vssd1 vccd1 vccd1 _11710_/A sky130_fd_sc_hd__or2_2
XFILLER_0_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12688_ reg1_val[10] _12689_/B vssd1 vssd1 vccd1 vccd1 _12699_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_126_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11639_ reg1_val[19] curr_PC[19] vssd1 vssd1 vccd1 vccd1 _11640_/B sky130_fd_sc_hd__or2_1
XFILLER_0_71_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09946__A _10479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13309_ _13309_/CLK _13309_/D vssd1 vssd1 vccd1 vccd1 hold198/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08850_ _08850_/A _08850_/B vssd1 vssd1 vccd1 vccd1 _08854_/A sky130_fd_sc_hd__xor2_1
X_07801_ _07869_/A _07869_/B _07794_/X vssd1 vssd1 vccd1 vccd1 _07822_/A sky130_fd_sc_hd__a21o_1
XANTENNA__06772__B1 _06771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13098__B1 _13254_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08781_ _08790_/B _08791_/A _08781_/C vssd1 vssd1 vccd1 vccd1 _08783_/A sky130_fd_sc_hd__nand3_1
XANTENNA__08513__A1 _08598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07732_ _07750_/A _07730_/Y _07711_/Y vssd1 vssd1 vccd1 vccd1 _07743_/B sky130_fd_sc_hd__o21a_1
XANTENNA__08513__B2 _08538_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07663_ _07663_/A _07663_/B vssd1 vssd1 vccd1 vccd1 _07666_/A sky130_fd_sc_hd__or2_2
X_06614_ instruction[41] _06927_/B _06612_/X vssd1 vssd1 vccd1 vccd1 _06783_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_94_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09402_ _09400_/X _09401_/X _09727_/S vssd1 vssd1 vccd1 vccd1 _09402_/X sky130_fd_sc_hd__mux2_1
X_07594_ _12224_/A _07361_/B _11844_/A vssd1 vssd1 vccd1 vccd1 _07596_/A sky130_fd_sc_hd__a21o_1
X_09333_ _09335_/A _09335_/B vssd1 vssd1 vccd1 vccd1 _09333_/X sky130_fd_sc_hd__or2_1
XFILLER_0_63_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08816__A2 _07217_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09264_ _09281_/B _09090_/B _09101_/B _09102_/B _09102_/A vssd1 vssd1 vccd1 vccd1
+ _09280_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_118_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13022__B1 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09195_ _12644_/A reg1_val[30] _09211_/S vssd1 vssd1 vccd1 vccd1 _09195_/X sky130_fd_sc_hd__mux2_1
X_08215_ _08215_/A _08215_/B vssd1 vssd1 vccd1 vccd1 _08216_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_43_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08146_ _08576_/A2 _08289_/B fanout75/X _09472_/A vssd1 vssd1 vccd1 vccd1 _08147_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_113_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12282__A _12335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08077_ _08794_/A _08790_/A vssd1 vssd1 vccd1 vccd1 _08077_/X sky130_fd_sc_hd__or2_1
X_07028_ _09672_/A _07029_/B vssd1 vssd1 vccd1 vccd1 _07030_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_11_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__buf_1
XANTENNA__07555__A2 _07554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ _09947_/A _08979_/B vssd1 vssd1 vccd1 vccd1 _08981_/B sky130_fd_sc_hd__xnor2_4
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ _11990_/A1 _12065_/B hold201/A vssd1 vssd1 vccd1 vccd1 _11990_/Y sky130_fd_sc_hd__a21oi_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11626__A _11841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10941_ _12093_/A _10941_/B vssd1 vssd1 vccd1 vccd1 _10943_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_98_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12611_ _12611_/A _12611_/B vssd1 vssd1 vccd1 vccd1 _12612_/A sky130_fd_sc_hd__nor2_1
X_10872_ _10872_/A _10872_/B vssd1 vssd1 vccd1 vccd1 _10874_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12542_ _12702_/B _12543_/B vssd1 vssd1 vccd1 vccd1 _12553_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10614__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11080__B fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12473_ _12650_/B _12473_/B vssd1 vssd1 vccd1 vccd1 _12474_/B sky130_fd_sc_hd__or2_1
X_11424_ _11424_/A _11424_/B vssd1 vssd1 vccd1 vccd1 _11426_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_123_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11575__B1 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_8 reg1_val[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11355_ _11262_/X _11354_/Y _12064_/S vssd1 vssd1 vccd1 vccd1 _11355_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08440__B1 _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10306_ _07222_/A _12422_/A _10304_/Y _10305_/X vssd1 vssd1 vccd1 vccd1 _10306_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_11286_ _07200_/X fanout8/X _11285_/Y vssd1 vssd1 vccd1 vccd1 _11288_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__08991__A1 _09325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08991__B2 _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13025_ _13249_/A hold163/X vssd1 vssd1 vccd1 vccd1 hold164/A sky130_fd_sc_hd__and2_1
X_10237_ _10237_/A _10237_/B vssd1 vssd1 vccd1 vccd1 _10253_/A sky130_fd_sc_hd__xnor2_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10168_ hold211/A _11538_/A _10300_/B _12205_/B1 vssd1 vssd1 vccd1 vccd1 _10169_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09940__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10099_ _10100_/A _10100_/B vssd1 vssd1 vccd1 vccd1 _10265_/A sky130_fd_sc_hd__and2_1
XANTENNA__09006__A _09836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12809_ hold11/X _12820_/B _12808_/Y _13039_/A vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__o211a_1
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13004__B1 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07482__A1 _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07482__B2 _08613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08000_ _08000_/A _08000_/B vssd1 vssd1 vccd1 vccd1 _08001_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_13_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12814__B _12820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08580__A _08580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09951_ _10623_/A _09951_/B vssd1 vssd1 vccd1 vccd1 _09959_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__07785__A2 fanout86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08902_ _07592_/A _07591_/B _07591_/A vssd1 vssd1 vccd1 vccd1 _08907_/A sky130_fd_sc_hd__o21bai_4
X_09882_ _09182_/X _09206_/X _10295_/S vssd1 vssd1 vccd1 vccd1 _09882_/X sky130_fd_sc_hd__mux2_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ _08833_/A _08833_/B vssd1 vssd1 vccd1 vccd1 _08834_/B sky130_fd_sc_hd__xor2_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08764_ _08759_/B _08759_/C _08759_/A _08761_/B vssd1 vssd1 vccd1 vccd1 _08765_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07715_ _10092_/A _07715_/B vssd1 vssd1 vccd1 vccd1 _07717_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08695_ _08013_/A _08013_/B _08076_/A _08076_/B vssd1 vssd1 vccd1 vccd1 _08695_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07646_ _07241_/A _07241_/B _07227_/A vssd1 vssd1 vccd1 vccd1 _07658_/A sky130_fd_sc_hd__a21oi_2
X_07577_ _10337_/A fanout29/X _07238_/Y _07959_/B vssd1 vssd1 vccd1 vccd1 _07578_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10057__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09316_ _09316_/A _09316_/B vssd1 vssd1 vccd1 vccd1 _09319_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_90_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09247_ _10297_/S _09250_/B vssd1 vssd1 vccd1 vccd1 _09248_/B sky130_fd_sc_hd__or2_1
XFILLER_0_35_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09178_ _09176_/X _09177_/X _09403_/S vssd1 vssd1 vccd1 vccd1 _09178_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08129_ _08575_/A _08129_/B vssd1 vssd1 vccd1 vccd1 _08198_/B sky130_fd_sc_hd__xnor2_1
X_11140_ _10165_/S _09437_/Y _11139_/X vssd1 vssd1 vccd1 vccd1 _11141_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_31_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11071_ _07013_/X _07171_/A fanout38/X _11779_/A vssd1 vssd1 vccd1 vccd1 _11072_/B
+ sky130_fd_sc_hd__a22o_1
X_10022_ _10295_/S _10022_/B vssd1 vssd1 vccd1 vccd1 _10022_/X sky130_fd_sc_hd__or2_1
XFILLER_0_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11973_ _11973_/A _12049_/B vssd1 vssd1 vccd1 vccd1 _11973_/Y sky130_fd_sc_hd__nor2_1
X_10924_ hold288/A _10924_/B vssd1 vssd1 vccd1 vccd1 _11035_/B sky130_fd_sc_hd__or2_1
XFILLER_0_58_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10855_ _12233_/A fanout28/X fanout26/X _12087_/A vssd1 vssd1 vccd1 vccd1 _10856_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_94_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08384__B _08384_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12525_ _12525_/A _12525_/B _12525_/C vssd1 vssd1 vccd1 vccd1 _12526_/B sky130_fd_sc_hd__nand3_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ _10703_/X _11050_/B _10785_/Y vssd1 vssd1 vccd1 vccd1 _10818_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12456_ _09236_/Y _12448_/Y _12455_/X vssd1 vssd1 vccd1 vccd1 _12456_/X sky130_fd_sc_hd__a21o_1
X_11407_ _11407_/A _11407_/B vssd1 vssd1 vccd1 vccd1 _11409_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12387_ _08859_/Y _11946_/C _12385_/X _12434_/S vssd1 vssd1 vccd1 vccd1 _12389_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11338_ _10416_/A _10902_/X _11334_/X _11337_/X vssd1 vssd1 vccd1 vccd1 _11340_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_9_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13369_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11269_ _12471_/S _11375_/C vssd1 vssd1 vccd1 vccd1 _11269_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08716__A1 _08575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07519__A2 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13008_ hold204/A _13171_/B2 _13209_/A2 hold177/X vssd1 vssd1 vccd1 vccd1 hold178/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12276__A1 _09221_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12276__B2 _12379_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07500_ _07501_/A _07501_/B vssd1 vssd1 vccd1 vccd1 _07500_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08575__A _08575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08480_ _08480_/A _08480_/B vssd1 vssd1 vccd1 vccd1 _08511_/B sky130_fd_sc_hd__xnor2_2
X_07431_ _07403_/Y _07431_/B vssd1 vssd1 vccd1 vccd1 _07678_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_85_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06807__B _07172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07362_ _12808_/A _07362_/B vssd1 vssd1 vccd1 vccd1 _07588_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_72_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09101_ _09101_/A _09101_/B vssd1 vssd1 vccd1 vccd1 _09102_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_127_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07293_ _07663_/A _07293_/B vssd1 vssd1 vccd1 vccd1 _07310_/A sky130_fd_sc_hd__nor2_1
X_09032_ _09032_/A _09032_/B vssd1 vssd1 vccd1 vccd1 _09034_/B sky130_fd_sc_hd__xor2_4
Xhold300 hold300/A vssd1 vssd1 vccd1 vccd1 hold300/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08955__A1 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07758__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08955__B2 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07357__C _07357_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09934_ _09934_/A _11497_/A vssd1 vssd1 vccd1 vccd1 _09938_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_0_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09904__B1 _09886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09865_ _09546_/X _09705_/X _09706_/X vssd1 vssd1 vccd1 vccd1 _09865_/X sky130_fd_sc_hd__a21o_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08816_ _07830_/B _07217_/Y _07221_/X fanout46/X vssd1 vssd1 vccd1 vccd1 _08817_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ _10246_/A _09796_/B vssd1 vssd1 vccd1 vccd1 _09797_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07391__B1 _07282_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12267__A1 _12447_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08747_ _08741_/A _08741_/B _08741_/C _08683_/B _08492_/X vssd1 vssd1 vccd1 vccd1
+ _08749_/C sky130_fd_sc_hd__a311o_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08678_ _08678_/A _08678_/B _08678_/C vssd1 vssd1 vccd1 vccd1 _08730_/A sky130_fd_sc_hd__and3_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12719__B _12719_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07694__A1 _06993_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07629_ _07417_/B _07166_/Y _07173_/Y fanout42/X vssd1 vssd1 vccd1 vccd1 _07630_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06717__B _12650_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10640_ _10528_/A _10528_/B _10526_/X vssd1 vssd1 vccd1 vccd1 _10647_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07694__B2 _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10571_ hold294/A _09425_/C _10690_/B _12416_/C1 vssd1 vssd1 vccd1 vccd1 _10571_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__07446__B2 _10599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07446__A1 _07198_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13290_ _13390_/CLK _13290_/D vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12310_ _06645_/B _06669_/Y _06643_/X vssd1 vssd1 vccd1 vccd1 _12310_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12990__A2 _13000_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12241_ _12243_/A _12243_/B _12243_/C vssd1 vssd1 vccd1 vccd1 _12244_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__06957__B1 _06723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12172_ _12172_/A _12172_/B vssd1 vssd1 vccd1 vccd1 _12173_/B sky130_fd_sc_hd__and2_1
XFILLER_0_102_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11123_ max_cap3/X _11122_/X _11121_/X vssd1 vssd1 vccd1 vccd1 _11124_/B sky130_fd_sc_hd__a21oi_4
X_11054_ _10966_/A _10966_/B _10963_/A vssd1 vssd1 vccd1 vccd1 _11060_/A sky130_fd_sc_hd__a21o_1
XANTENNA__10505__B2 _07256_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10505__A1 _07097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10005_ _09376_/B _10004_/Y _10003_/X vssd1 vssd1 vccd1 vccd1 _10006_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07382__B1 fanout72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11956_ _11957_/A _11957_/B vssd1 vssd1 vccd1 vccd1 _12040_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10907_ _11809_/A _08744_/A _08744_/B vssd1 vssd1 vccd1 vccd1 _10907_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07685__A1 _09943_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11887_ _11710_/A _11796_/X _11798_/B vssd1 vssd1 vccd1 vccd1 _11887_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__11481__A2 _07171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06627__B _12708_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07685__B2 _08538_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10838_ _10838_/A _10838_/B vssd1 vssd1 vccd1 vccd1 _10879_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10769_ _10770_/B _10770_/A vssd1 vssd1 vccd1 vccd1 _10769_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13240__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12508_ _12675_/B _12508_/B vssd1 vssd1 vccd1 vccd1 _12509_/B sky130_fd_sc_hd__or2_1
XFILLER_0_89_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12439_ _12438_/A _06888_/X _12406_/X _12438_/Y vssd1 vssd1 vccd1 vccd1 _12439_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10744__B2 _08411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10744__A1 _10476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07980_ _08564_/A _07980_/B vssd1 vssd1 vccd1 vccd1 _08023_/B sky130_fd_sc_hd__xnor2_1
Xfanout109 _07237_/Y vssd1 vssd1 vccd1 vccd1 _08501_/B1 sky130_fd_sc_hd__buf_6
X_06931_ instruction[14] _06933_/B vssd1 vssd1 vccd1 vccd1 dest_idx[3] sky130_fd_sc_hd__and2_4
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09650_ _09650_/A _10476_/B _10476_/C vssd1 vssd1 vccd1 vccd1 _09652_/C sky130_fd_sc_hd__or3_1
XANTENNA__08289__B _08289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06862_ _06860_/X _06861_/Y _06700_/A vssd1 vssd1 vccd1 vccd1 _06862_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09901__A3 _11995_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08601_ _08609_/A _08609_/B vssd1 vssd1 vccd1 vccd1 _08610_/A sky130_fd_sc_hd__nand2_1
X_06793_ _06815_/A _06817_/B1 _12665_/B _06791_/X vssd1 vssd1 vccd1 vccd1 _06793_/Y
+ sky130_fd_sc_hd__a31oi_2
X_09581_ _09581_/A _09581_/B vssd1 vssd1 vccd1 vccd1 _09581_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__09114__B2 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09114__A1 _08112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08532_ _08535_/A _08535_/B vssd1 vssd1 vccd1 vccd1 _08532_/X sky130_fd_sc_hd__or2_1
XANTENNA__06818__A _06992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08463_ _08469_/A _08469_/B vssd1 vssd1 vccd1 vccd1 _08464_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_77_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout153_A _07015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07414_ _07414_/A _07414_/B vssd1 vssd1 vccd1 vccd1 _07426_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_92_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08394_ _08421_/A _08394_/B vssd1 vssd1 vccd1 vccd1 _08436_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12421__A1 _12421_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07345_ _09779_/A _07345_/B vssd1 vssd1 vccd1 vccd1 _07349_/A sky130_fd_sc_hd__xor2_1
XANTENNA__13150__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07276_ _09667_/A _07276_/B vssd1 vssd1 vccd1 vccd1 _07278_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07979__A2 _10338_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09015_ _09016_/A _09016_/B vssd1 vssd1 vccd1 vccd1 _09017_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12185__B1 _11892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08928__A1 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10735__A1 _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold141 hold141/A vssd1 vssd1 vccd1 vccd1 hold141/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 hold152/A vssd1 vssd1 vccd1 vccd1 hold152/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 hold130/A vssd1 vssd1 vccd1 vccd1 hold130/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12724__A2 _12719_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08928__B2 _07830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold163 hold163/A vssd1 vssd1 vccd1 vccd1 hold163/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 hold174/A vssd1 vssd1 vccd1 vccd1 hold174/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10735__B2 _12009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold185 hold185/A vssd1 vssd1 vccd1 vccd1 hold185/X sky130_fd_sc_hd__dlygate4sd3_1
X_09917_ _11393_/A _09917_/B vssd1 vssd1 vccd1 vccd1 _09919_/B sky130_fd_sc_hd__xnor2_1
Xhold196 hold196/A vssd1 vssd1 vccd1 vccd1 hold196/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08199__B _08199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout66_A _06997_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09848_ _09690_/A _09689_/B _09687_/Y vssd1 vssd1 vccd1 vccd1 _09858_/A sky130_fd_sc_hd__a21o_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _09779_/A _09779_/B vssd1 vssd1 vccd1 vccd1 _09780_/B sky130_fd_sc_hd__xor2_1
XANTENNA__11634__A _12359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12790_ reg1_val[30] _12790_/B vssd1 vssd1 vccd1 vccd1 _12791_/B sky130_fd_sc_hd__or2_1
XANTENNA__09105__A1 _07172_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11810_ _11810_/A _11810_/B vssd1 vssd1 vccd1 vccd1 _11810_/X sky130_fd_sc_hd__xor2_1
XANTENNA__09105__B2 _09325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11741_ hold274/A _11650_/B _11822_/B _12376_/C1 vssd1 vssd1 vccd1 vccd1 _11741_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_96_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09656__A2 _10245_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11672_ _11764_/C _11672_/B vssd1 vssd1 vccd1 vccd1 _11674_/B sky130_fd_sc_hd__xnor2_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10623_ _10623_/A _10623_/B vssd1 vssd1 vccd1 vccd1 _10627_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__12465__A _12645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08616__B1 _07173_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10554_ _06834_/X _10553_/X _12054_/S vssd1 vssd1 vccd1 vccd1 _10554_/X sky130_fd_sc_hd__mux2_1
X_13342_ _13360_/CLK hold132/X vssd1 vssd1 vccd1 vccd1 hold130/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10485_ _10485_/A _10485_/B vssd1 vssd1 vccd1 vccd1 _10487_/B sky130_fd_sc_hd__xnor2_1
X_13273_ _13369_/CLK _13273_/D vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12224_ _12224_/A _12224_/B vssd1 vssd1 vccd1 vccd1 _12225_/B sky130_fd_sc_hd__nand2_1
X_12155_ _12086_/B _12088_/B _12086_/A vssd1 vssd1 vccd1 vccd1 _12167_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__12404__S _12404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11106_ _11106_/A _11106_/B vssd1 vssd1 vccd1 vccd1 _11107_/B sky130_fd_sc_hd__xor2_2
X_12086_ _12086_/A _12086_/B vssd1 vssd1 vccd1 vccd1 _12088_/A sky130_fd_sc_hd__nand2_1
X_11037_ hold270/A _11650_/B _11143_/B _12376_/C1 vssd1 vssd1 vccd1 vccd1 _11037_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11151__A1 _12421_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12988_ hold211/X _13000_/A2 _13257_/A2 hold215/X vssd1 vssd1 vccd1 vccd1 hold216/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09647__A2 _10473_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11939_ _11939_/A _11939_/B vssd1 vssd1 vccd1 vccd1 _11940_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07122__A3 _12740_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07130_ _07129_/A _07129_/B _07129_/C _07129_/D vssd1 vssd1 vccd1 vccd1 _11854_/A
+ sky130_fd_sc_hd__o22ai_2
XFILLER_0_15_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07061_ reg1_val[4] reg1_val[5] vssd1 vssd1 vccd1 vccd1 _07083_/D sky130_fd_sc_hd__or2_1
XFILLER_0_11_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11719__A _11884_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12822__B _12826_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09583__A1 _12322_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11390__B2 _07013_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11390__A1 _11946_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10623__A _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07594__B1 _11844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07963_ _09472_/A _08112_/B fanout25/X _08649_/B1 vssd1 vssd1 vccd1 vccd1 _07964_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08138__A2 _10338_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06914_ reg1_idx[5] _12218_/A vssd1 vssd1 vccd1 vccd1 _06915_/D sky130_fd_sc_hd__and2_1
XANTENNA__11142__A1 _11820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13131__A2 _13254_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09702_ _09703_/A _09703_/B vssd1 vssd1 vccd1 vccd1 _09702_/X sky130_fd_sc_hd__and2_1
X_07894_ _09836_/A _07894_/B vssd1 vssd1 vccd1 vccd1 _07896_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07346__B1 _07283_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06845_ _07270_/A _11134_/A vssd1 vssd1 vccd1 vccd1 _06845_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_65_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09633_ _09633_/A _09633_/B vssd1 vssd1 vccd1 vccd1 _09636_/A sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout270_A _06927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13145__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09564_ _09166_/X _09171_/X _09727_/S vssd1 vssd1 vccd1 vccd1 _09564_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06776_ reg2_val[6] _06810_/B vssd1 vssd1 vccd1 vccd1 _06776_/X sky130_fd_sc_hd__and2_1
X_08515_ _09404_/S _08515_/A2 _08649_/B1 _10245_/B2 vssd1 vssd1 vccd1 vccd1 _08516_/B
+ sky130_fd_sc_hd__o22a_1
X_09495_ _09495_/A _09495_/B vssd1 vssd1 vccd1 vccd1 _09498_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07649__B2 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07649__A1 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08446_ _08580_/A _08446_/B vssd1 vssd1 vccd1 vccd1 _08471_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08377_ _08424_/A _08424_/B _08372_/X vssd1 vssd1 vccd1 vccd1 _08384_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_61_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07379__A _10749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07328_ fanout51/X _10245_/B2 _10245_/A1 _09661_/B2 vssd1 vssd1 vccd1 vccd1 _07329_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07259_ _06974_/X _06978_/C _06978_/D _07215_/B vssd1 vssd1 vccd1 vccd1 _07270_/B
+ sky130_fd_sc_hd__o31ai_4
XFILLER_0_61_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09594__A _12438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10270_ _10270_/A _10270_/B vssd1 vssd1 vccd1 vccd1 _10272_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09326__A1 _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13122__A2 _13254_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09326__B2 _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07337__B1 _10245_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12911_ hold245/X hold154/X vssd1 vssd1 vccd1 vccd1 _13106_/A sky130_fd_sc_hd__xnor2_1
Xmax_cap9 _08974_/Y vssd1 vssd1 vccd1 vccd1 _12158_/B sky130_fd_sc_hd__buf_4
XFILLER_0_69_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08657__B _08657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12842_ hold87/X _12862_/B vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__or2_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _12769_/B _12772_/B _12767_/X vssd1 vssd1 vccd1 vccd1 _12775_/A sky130_fd_sc_hd__a21o_1
XANTENNA__08837__B1 _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11724_ _11636_/A _11634_/B _11652_/S vssd1 vssd1 vccd1 vccd1 _11724_/Y sky130_fd_sc_hd__o21bai_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11655_ _12379_/B2 _10914_/X _11643_/B _09221_/Y _11654_/Y vssd1 vssd1 vccd1 vccd1
+ _11655_/X sky130_fd_sc_hd__a221o_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06863__A2 _07036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout91 _11398_/A vssd1 vssd1 vccd1 vccd1 _09922_/A sky130_fd_sc_hd__buf_8
Xfanout80 _11198_/A vssd1 vssd1 vccd1 vccd1 fanout80/X sky130_fd_sc_hd__buf_6
XANTENNA__07289__A _09341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11586_ _11586_/A _11586_/B vssd1 vssd1 vccd1 vccd1 _11587_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_107_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10606_ _10606_/A _10606_/B vssd1 vssd1 vccd1 vccd1 _10609_/A sky130_fd_sc_hd__xor2_1
XANTENNA__09801__A2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13325_ _13392_/CLK _13325_/D vssd1 vssd1 vccd1 vccd1 hold227/A sky130_fd_sc_hd__dfxtp_1
X_10537_ _10538_/A _10538_/B _10538_/C vssd1 vssd1 vccd1 vccd1 _10539_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_12_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10468_ _10468_/A _10468_/B _10468_/C vssd1 vssd1 vccd1 vccd1 _10469_/B sky130_fd_sc_hd__and3_1
X_13256_ _13259_/A _13256_/B hold306/X vssd1 vssd1 vccd1 vccd1 hold307/A sky130_fd_sc_hd__and3_1
XANTENNA__12149__B1 _12148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12207_ _09228_/X _09234_/X _12207_/S vssd1 vssd1 vccd1 vccd1 _12207_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12642__B _12642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08368__A2 _10595_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06640__B _06675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13187_ _13210_/A hold247/X vssd1 vssd1 vccd1 vccd1 _13378_/D sky130_fd_sc_hd__and2_1
X_10399_ _10260_/A _10259_/B _10259_/A vssd1 vssd1 vccd1 vccd1 _10409_/A sky130_fd_sc_hd__o21bai_1
X_12138_ hold276/A _12449_/B1 _12199_/B _12416_/C1 vssd1 vssd1 vccd1 vccd1 _12139_/B
+ sky130_fd_sc_hd__a31o_1
X_12069_ _12449_/B1 _12136_/B hold278/A vssd1 vssd1 vccd1 vccd1 _12069_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__13113__A2 _13254_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09317__A1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09317__B2 _09661_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07328__B1 _10245_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08848__A _10092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06630_ reg1_val[28] _08973_/B vssd1 vssd1 vccd1 vccd1 _06630_/X sky130_fd_sc_hd__and2_1
XFILLER_0_79_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08300_ _08349_/A _08349_/B _08296_/X vssd1 vssd1 vccd1 vccd1 _08311_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_19_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09280_ _09280_/A _09280_/B vssd1 vssd1 vccd1 vccd1 _09354_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08231_ _08231_/A _08231_/B vssd1 vssd1 vccd1 vccd1 _08234_/A sky130_fd_sc_hd__or2_2
XFILLER_0_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06815__B _12645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10938__A1 _11406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10337__B _12428_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08162_ _08162_/A _08162_/B vssd1 vssd1 vccd1 vccd1 _08186_/B sky130_fd_sc_hd__xor2_2
XANTENNA__10938__B2 _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07113_ _07248_/A _07140_/C vssd1 vssd1 vccd1 vccd1 _07115_/C sky130_fd_sc_hd__and2_1
XFILLER_0_70_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08093_ _08122_/A _08122_/B vssd1 vssd1 vccd1 vccd1 _08098_/A sky130_fd_sc_hd__or2_1
XFILLER_0_42_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07044_ _07604_/A _07044_/B vssd1 vssd1 vccd1 vccd1 _07059_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09005__B1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10072__B fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08995_ _11844_/A _08995_/B vssd1 vssd1 vccd1 vccd1 _08997_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07946_ _07946_/A _07946_/B _07946_/C vssd1 vssd1 vccd1 vccd1 _07947_/B sky130_fd_sc_hd__or3_1
XANTENNA__12863__A1 _07051_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10800__B _11820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07877_ _07877_/A _07947_/A _07877_/C vssd1 vssd1 vccd1 vccd1 _07877_/X sky130_fd_sc_hd__and3_1
X_06828_ _10014_/A _06826_/Y _06827_/Y vssd1 vssd1 vccd1 vccd1 _06828_/X sky130_fd_sc_hd__o21a_1
X_09616_ _09779_/A _09616_/B vssd1 vssd1 vccd1 vccd1 _09617_/B sky130_fd_sc_hd__xor2_1
XANTENNA__12076__C1 _12058_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06759_ _06759_/A _10688_/S vssd1 vssd1 vccd1 vccd1 _10672_/A sky130_fd_sc_hd__nor2_1
X_09547_ _09548_/A _09548_/B vssd1 vssd1 vccd1 vccd1 _09547_/X sky130_fd_sc_hd__and2_1
XFILLER_0_78_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout29_A fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09478_ _09478_/A _09478_/B vssd1 vssd1 vccd1 vccd1 _09510_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12379__B1 _09596_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_11_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13358_/CLK sky130_fd_sc_hd__clkbuf_8
X_08429_ _08435_/B _08435_/A vssd1 vssd1 vccd1 vccd1 _08429_/X sky130_fd_sc_hd__and2b_1
X_11440_ _11618_/A _11440_/B vssd1 vssd1 vccd1 vccd1 _11840_/C sky130_fd_sc_hd__xnor2_4
XANTENNA__10929__A1 _07195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09795__A1 _10245_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09795__B2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11371_ curr_PC[16] _11375_/C vssd1 vssd1 vccd1 vccd1 _11371_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_33_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13110_ _13110_/A _13110_/B vssd1 vssd1 vccd1 vccd1 _13111_/B sky130_fd_sc_hd__nand2_1
X_10322_ _09869_/A _09869_/B _09765_/B vssd1 vssd1 vccd1 vccd1 _10324_/C sky130_fd_sc_hd__o21ba_1
XFILLER_0_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13041_ _08656_/A _13101_/B2 hold126/X vssd1 vssd1 vccd1 vccd1 _13330_/D sky130_fd_sc_hd__o21a_1
X_10253_ _10253_/A _10383_/B _10253_/C vssd1 vssd1 vccd1 vccd1 _10255_/B sky130_fd_sc_hd__and3_1
X_10184_ curr_PC[6] _10184_/B vssd1 vssd1 vccd1 vccd1 _10448_/C sky130_fd_sc_hd__and2_2
Xfanout270 _06927_/A vssd1 vssd1 vccd1 vccd1 _06815_/A sky130_fd_sc_hd__buf_8
Xfanout281 _13142_/A vssd1 vssd1 vccd1 vccd1 _13259_/A sky130_fd_sc_hd__buf_4
Xfanout292 _09218_/A vssd1 vssd1 vccd1 vccd1 _12642_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12825_ _10337_/A _13089_/A2 hold31/X _13142_/A vssd1 vssd1 vccd1 vccd1 _13273_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12082__A2 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10093__A1 _11671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _12756_/A _12760_/D vssd1 vssd1 vccd1 vccd1 loadstore_address[23] sky130_fd_sc_hd__xnor2_4
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11707_ _11610_/A _11610_/B _11613_/A vssd1 vssd1 vccd1 vccd1 _11709_/B sky130_fd_sc_hd__a21oi_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10093__B2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12687_ _12687_/A _12687_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[9] sky130_fd_sc_hd__xor2_4
XFILLER_0_21_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11638_ reg1_val[19] curr_PC[19] vssd1 vssd1 vccd1 vccd1 _11640_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11569_ _12336_/A _11569_/B vssd1 vssd1 vccd1 vccd1 _11573_/B sky130_fd_sc_hd__xnor2_1
X_13308_ _13309_/CLK hold187/X vssd1 vssd1 vccd1 vccd1 hold185/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07797__B1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13239_ _13239_/A _13239_/B vssd1 vssd1 vccd1 vccd1 _13239_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__11269__A _12471_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07800_ _07800_/A _07800_/B vssd1 vssd1 vccd1 vccd1 _07869_/B sky130_fd_sc_hd__xnor2_1
X_08780_ _08772_/B _08772_/C _08779_/X vssd1 vssd1 vccd1 vccd1 _08781_/C sky130_fd_sc_hd__a21o_1
X_07731_ _07731_/A _07731_/B vssd1 vssd1 vccd1 vccd1 _07750_/B sky130_fd_sc_hd__xor2_1
XANTENNA__12845__A1 _07983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08513__A2 _08576_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07662_ _07180_/Y _07242_/B _07243_/X vssd1 vssd1 vccd1 vccd1 _07667_/A sky130_fd_sc_hd__o21ai_4
X_06613_ instruction[1] instruction[2] instruction[25] pred_val vssd1 vssd1 vccd1
+ vccd1 _06613_/Y sky130_fd_sc_hd__o211ai_1
X_09401_ _09204_/X _09207_/X _09403_/S vssd1 vssd1 vccd1 vccd1 _09401_/X sky130_fd_sc_hd__mux2_1
X_07593_ _07340_/A _07339_/Y _07335_/Y vssd1 vssd1 vccd1 vccd1 _07599_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_47_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09332_ _09332_/A _09332_/B vssd1 vssd1 vccd1 vccd1 _09335_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12073__A2 _12422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10348__A _10748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09263_ _09139_/A _09139_/B _09140_/Y vssd1 vssd1 vccd1 vccd1 _09369_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09194_ _09192_/X _09193_/X _09419_/B vssd1 vssd1 vccd1 vccd1 _09194_/X sky130_fd_sc_hd__mux2_1
X_08214_ _08224_/A _08224_/B vssd1 vssd1 vccd1 vccd1 _08214_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08145_ _08454_/A _08145_/B vssd1 vssd1 vccd1 vccd1 _08150_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__12563__A _12719_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08076_ _08076_/A _08076_/B vssd1 vssd1 vccd1 vccd1 _08790_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11179__A _11179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10083__A _12224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07027_ _09672_/A _07029_/B vssd1 vssd1 vccd1 vccd1 _07031_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13089__A1 _09922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07392__A _09836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08978_ fanout68/X _09301_/A fanout56/X _07011_/Y vssd1 vssd1 vccd1 vccd1 _08979_/B
+ sky130_fd_sc_hd__o22a_2
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ _07969_/A _07929_/B vssd1 vssd1 vccd1 vccd1 _08003_/B sky130_fd_sc_hd__xnor2_1
X_10940_ _11779_/A _07171_/A fanout38/X _11764_/A vssd1 vssd1 vccd1 vccd1 _10941_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07712__B1 _10476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12610_ _12595_/B _12603_/B _12633_/A vssd1 vssd1 vccd1 vccd1 _12623_/B sky130_fd_sc_hd__o21ai_2
X_10871_ _10871_/A _12087_/B vssd1 vssd1 vccd1 vccd1 _10872_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_93_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06736__A _11134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12541_ reg1_val[12] curr_PC[12] _12638_/S vssd1 vssd1 vccd1 vccd1 _12543_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_54_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12472_ _12650_/B _12473_/B vssd1 vssd1 vccd1 vccd1 _12483_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_53_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11423_ _11424_/A _11424_/B vssd1 vssd1 vccd1 vccd1 _11520_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_124_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11575__B2 _07032_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11575__A1 _06998_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12473__A _12650_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_9 reg1_val[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11354_ _11354_/A _11354_/B vssd1 vssd1 vccd1 vccd1 _11354_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__08440__A1 _08540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08440__B2 _08515_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10305_ hold281/A _09425_/C _10569_/C _12416_/C1 vssd1 vssd1 vccd1 vccd1 _10305_/X
+ sky130_fd_sc_hd__a31o_1
X_11285_ _07192_/B fanout8/X _10092_/A vssd1 vssd1 vccd1 vccd1 _11285_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__08991__A2 _08877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13024_ hold162/X _13171_/B2 _13223_/A2 _13322_/Q vssd1 vssd1 vccd1 vccd1 hold163/A
+ sky130_fd_sc_hd__a22o_1
X_10236_ _10237_/A _10237_/B vssd1 vssd1 vccd1 vccd1 _10376_/B sky130_fd_sc_hd__nand2b_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09940__A1 _07221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10167_ _11538_/A _10300_/B hold211/A vssd1 vssd1 vccd1 vccd1 _10169_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__09940__B2 _09940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12827__A1 _07238_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10098_ _09942_/A _09942_/B _09939_/A vssd1 vssd1 vccd1 vccd1 _10100_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10302__A2 _11990_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13252__B2 _06577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12808_ _12808_/A _12820_/B vssd1 vssd1 vccd1 vccd1 _12808_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11271__B _11271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12739_ _12739_/A _12739_/B _12739_/C _12739_/D vssd1 vssd1 vccd1 vccd1 _12742_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07482__A2 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09759__A1 _12365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11015__B1 _12356_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11566__A1 _11752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07477__A _09341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09950_ fanout65/X fanout86/X fanout82/X fanout59/X vssd1 vssd1 vccd1 vccd1 _09951_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08901_ _07645_/A _07645_/B _07659_/B _07660_/B _07660_/A vssd1 vssd1 vccd1 vccd1
+ _08911_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_110_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12830__B _12862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09881_ _09167_/X _09175_/X _10295_/S vssd1 vssd1 vccd1 vccd1 _09881_/X sky130_fd_sc_hd__mux2_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06745__A1 _06927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ _08833_/A _08833_/B vssd1 vssd1 vccd1 vccd1 _08832_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10350__B fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08763_ _08362_/Y _08433_/B _08691_/B vssd1 vssd1 vccd1 vccd1 _08765_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07714_ _07191_/X _12823_/A1 _07282_/Y _07202_/Y vssd1 vssd1 vccd1 vccd1 _07715_/B
+ sky130_fd_sc_hd__a22o_1
X_08694_ _08281_/X _08363_/X _08761_/A _08693_/X _08277_/X vssd1 vssd1 vccd1 vccd1
+ _08776_/B sky130_fd_sc_hd__o221a_2
XFILLER_0_79_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07645_ _07645_/A _07645_/B vssd1 vssd1 vccd1 vccd1 _07659_/A sky130_fd_sc_hd__nand2_1
X_07576_ _10092_/A _07576_/B vssd1 vssd1 vccd1 vccd1 _07580_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10057__B2 _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10057__A1 _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09315_ _09315_/A _09315_/B vssd1 vssd1 vccd1 vccd1 _09316_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_90_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09246_ _09246_/A vssd1 vssd1 vccd1 vccd1 _09248_/A sky130_fd_sc_hd__inv_2
XFILLER_0_8_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09177_ reg1_val[13] reg1_val[18] _09180_/S vssd1 vssd1 vccd1 vccd1 _09177_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_50_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08128_ _08657_/B fanout76/X fanout72/X _08649_/A2 vssd1 vssd1 vccd1 vccd1 _08129_/B
+ sky130_fd_sc_hd__o22a_1
X_08059_ _08059_/A _08059_/B vssd1 vssd1 vccd1 vccd1 _08070_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11070_ _11070_/A _11070_/B vssd1 vssd1 vccd1 vccd1 _11088_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_113_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout96_A _09834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10021_ _11246_/S _10017_/X _10020_/Y _11029_/S vssd1 vssd1 vccd1 vccd1 _10021_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12740__B _12740_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11637__A _11637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11972_ _12113_/A _11972_/B vssd1 vssd1 vccd1 vccd1 _12049_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10923_ hold198/A _11990_/A1 _11032_/B _11648_/A vssd1 vssd1 vccd1 vccd1 _10923_/Y
+ sky130_fd_sc_hd__a31oi_1
X_10854_ _10854_/A _10854_/B vssd1 vssd1 vccd1 vccd1 _10858_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_109_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12524_ _12525_/A _12525_/B _12525_/C vssd1 vssd1 vccd1 vccd1 _12532_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_94_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10785_ _10703_/X _11050_/B _12356_/B1 vssd1 vssd1 vccd1 vccd1 _10785_/Y sky130_fd_sc_hd__o21ai_1
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12455_ _09152_/Y _09216_/X _12451_/Y _12454_/X vssd1 vssd1 vccd1 vccd1 _12455_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_50_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11406_ _11406_/A _12017_/A vssd1 vssd1 vccd1 vccd1 _11407_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_111_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12386_ _08859_/Y _12385_/X _12384_/Y vssd1 vssd1 vccd1 vccd1 _12434_/S sky130_fd_sc_hd__o21ai_1
XANTENNA__07297__A _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08413__A1 _10950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11337_ _10901_/X _11334_/X _11716_/A vssd1 vssd1 vccd1 vccd1 _11337_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_499 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11268_ curr_PC[15] _11268_/B vssd1 vssd1 vccd1 vccd1 _11375_/C sky130_fd_sc_hd__and2_1
XANTENNA__12650__B _12650_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11199_ _11199_/A _11199_/B vssd1 vssd1 vccd1 vccd1 _11201_/B sky130_fd_sc_hd__xnor2_1
X_13007_ _13019_/A hold205/X vssd1 vssd1 vccd1 vccd1 _13313_/D sky130_fd_sc_hd__and2_1
X_10219_ _10220_/A _10220_/B vssd1 vssd1 vccd1 vccd1 _10401_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_27_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12276__A2 _09880_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07430_ _07430_/A _07430_/B vssd1 vssd1 vccd1 vccd1 _07431_/B sky130_fd_sc_hd__nand2_1
X_07361_ _12224_/A _07361_/B vssd1 vssd1 vccd1 vccd1 _07361_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11236__B1 _10788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12984__B1 _13257_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09100_ _09330_/B _09100_/B vssd1 vssd1 vccd1 vccd1 _09101_/B sky130_fd_sc_hd__and2_2
XANTENNA__08101__B1 _09479_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07292_ _07292_/A _07292_/B _07374_/A vssd1 vssd1 vccd1 vccd1 _07293_/B sky130_fd_sc_hd__nor3_1
X_09031_ _09031_/A _09031_/B vssd1 vssd1 vccd1 vccd1 _09032_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_60_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06823__B _11138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold301 hold301/A vssd1 vssd1 vccd1 vccd1 hold301/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09601__B1 _12356_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07000__A _09672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08955__A2 _10245_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09933_ _09933_/A _09933_/B vssd1 vssd1 vccd1 vccd1 _09965_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_0_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09904__A1 _12379_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09864_ _09044_/A _09044_/B _09863_/X vssd1 vssd1 vccd1 vccd1 _09868_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08815_ _07599_/A _07599_/B _07602_/A vssd1 vssd1 vccd1 vccd1 _08826_/A sky130_fd_sc_hd__a21o_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09795_ _10245_/B2 _10476_/B _10476_/C _10245_/A1 fanout56/X vssd1 vssd1 vccd1 vccd1
+ _09796_/B sky130_fd_sc_hd__o32a_1
XANTENNA__07391__A1 _07121_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07391__B2 _07959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08746_ _08743_/A _08743_/B _08745_/X _08744_/A vssd1 vssd1 vccd1 vccd1 _08751_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11475__B1 _11591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ _08677_/A _08677_/B vssd1 vssd1 vccd1 vccd1 _08727_/B sky130_fd_sc_hd__xor2_2
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11192__A _11393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07694__A2 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08340__B1 _08457_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07628_ _07628_/A _07628_/B vssd1 vssd1 vccd1 vccd1 _07642_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07559_ _07559_/A _07559_/B vssd1 vssd1 vccd1 vccd1 _07681_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10570_ _09425_/C _10690_/B hold294/A vssd1 vssd1 vccd1 vccd1 _10570_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07446__A2 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09229_ _11637_/A _12420_/A0 _08663_/A vssd1 vssd1 vccd1 vccd1 _09229_/X sky130_fd_sc_hd__a21o_1
X_12240_ _12296_/B _12240_/B vssd1 vssd1 vccd1 vccd1 _12243_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_16_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12171_ _12172_/A _12172_/B vssd1 vssd1 vccd1 vccd1 _12243_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_32_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06957__A1 _12359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11122_ _11122_/A _11334_/A vssd1 vssd1 vccd1 vccd1 _11122_/X sky130_fd_sc_hd__and2_1
X_11053_ _10998_/A _10998_/B _10996_/Y vssd1 vssd1 vccd1 vccd1 _11115_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__10505__A2 _07171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10004_ _10004_/A _10137_/A _10137_/B _10331_/A vssd1 vssd1 vccd1 vccd1 _10004_/Y
+ sky130_fd_sc_hd__nor4_2
XANTENNA__07382__A1 fanout86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07382__B2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09659__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11955_ _11955_/A _11955_/B vssd1 vssd1 vccd1 vccd1 _11957_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10906_ _10824_/X _11050_/C _10905_/Y vssd1 vssd1 vccd1 vccd1 _10933_/A sky130_fd_sc_hd__o21a_1
XANTENNA__07685__A2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11886_ _11886_/A vssd1 vssd1 vccd1 vccd1 _11886_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_86_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10837_ _10838_/B _10838_/A vssd1 vssd1 vccd1 vccd1 _10837_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_13_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10768_ _10768_/A _10768_/B vssd1 vssd1 vccd1 vccd1 _10770_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12645__B _12645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12507_ _12675_/B _12508_/B vssd1 vssd1 vccd1 vccd1 _12518_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_81_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12438_ _12438_/A _12438_/B vssd1 vssd1 vccd1 vccd1 _12438_/Y sky130_fd_sc_hd__nor2_1
X_10699_ curr_PC[9] curr_PC[10] _10699_/C vssd1 vssd1 vccd1 vccd1 _10934_/C sky130_fd_sc_hd__and3_1
XFILLER_0_112_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10744__A2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12369_ _12412_/A _09562_/A _12368_/X _09242_/B vssd1 vssd1 vccd1 vccd1 _12369_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06930_ instruction[13] _06933_/B vssd1 vssd1 vccd1 vccd1 dest_idx[2] sky130_fd_sc_hd__and2_4
XANTENNA__11277__A _11584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06861_ reg1_val[22] _07014_/A vssd1 vssd1 vccd1 vccd1 _06861_/Y sky130_fd_sc_hd__nand2_1
X_08600_ _09670_/A _08600_/B vssd1 vssd1 vccd1 vccd1 _08609_/B sky130_fd_sc_hd__xnor2_1
X_06792_ _06815_/A _06817_/B1 _12665_/B _06791_/X vssd1 vssd1 vccd1 vccd1 _06792_/X
+ sky130_fd_sc_hd__a31o_1
X_09580_ _09578_/Y _09580_/B vssd1 vssd1 vccd1 vccd1 _09581_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_89_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11457__B1 _12421_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09114__A2 _11093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08531_ _09670_/A _08531_/B vssd1 vssd1 vccd1 vccd1 _08535_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08462_ _08462_/A _08462_/B vssd1 vssd1 vccd1 vccd1 _08469_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07413_ _07413_/A _07413_/B vssd1 vssd1 vccd1 vccd1 _07414_/B sky130_fd_sc_hd__and2_1
XFILLER_0_9_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08393_ _08393_/A _08393_/B vssd1 vssd1 vccd1 vccd1 _08436_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07344_ _07148_/Y fanout42/X _07173_/Y _07417_/B vssd1 vssd1 vccd1 vccd1 _07345_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06636__B1 _06783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10432__A1 _11029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07275_ fanout78/X fanout76/X fanout74/X fanout72/X vssd1 vssd1 vccd1 vccd1 _07276_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_103_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09014_ _09014_/A _09014_/B vssd1 vssd1 vccd1 vccd1 _09016_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12185__A1 _12050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08389__B1 _08576_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10735__A2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold142 hold142/A vssd1 vssd1 vccd1 vccd1 hold142/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 hold153/A vssd1 vssd1 vccd1 vccd1 hold153/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 hold131/A vssd1 vssd1 vccd1 vccd1 hold131/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 hold120/A vssd1 vssd1 vccd1 vccd1 hold120/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08928__A2 _07217_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold175 hold175/A vssd1 vssd1 vccd1 vccd1 hold175/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 hold164/A vssd1 vssd1 vccd1 vccd1 hold164/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 hold186/A vssd1 vssd1 vccd1 vccd1 hold186/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11187__A _11770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09916_ fanout47/X _11198_/A _11093_/A fanout45/X vssd1 vssd1 vccd1 vccd1 _09917_/B
+ sky130_fd_sc_hd__o22a_1
Xhold197 hold197/A vssd1 vssd1 vccd1 vccd1 hold197/X sky130_fd_sc_hd__dlygate4sd3_1
X_09847_ _09847_/A _09847_/B vssd1 vssd1 vccd1 vccd1 _09860_/A sky130_fd_sc_hd__xor2_4
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08561__B1 _08561_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09778_ _07417_/B _07232_/X _07238_/Y fanout42/X vssd1 vssd1 vccd1 vccd1 _09779_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout59_A _07033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08729_ _08678_/B _08678_/C _08678_/A vssd1 vssd1 vccd1 vccd1 _08730_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__09105__A2 _08877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11740_ _11650_/B _11822_/B hold274/A vssd1 vssd1 vccd1 vccd1 _11740_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11671_ _11671_/A _11946_/C vssd1 vssd1 vccd1 vccd1 _11672_/B sky130_fd_sc_hd__nand2_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10622_ _10476_/A fanout14/X fanout12/X _08411_/B vssd1 vssd1 vccd1 vccd1 _10623_/B
+ sky130_fd_sc_hd__o22a_1
X_13410_ instruction[4] vssd1 vssd1 vccd1 vccd1 sign_extend sky130_fd_sc_hd__buf_12
XFILLER_0_119_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10553_ _06768_/Y _10421_/X _06770_/B vssd1 vssd1 vccd1 vccd1 _10553_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_64_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13341_ _13360_/CLK hold84/X vssd1 vssd1 vccd1 vccd1 _13341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10484_ _10485_/A _10485_/B vssd1 vssd1 vccd1 vccd1 _10484_/Y sky130_fd_sc_hd__nand2_1
X_13272_ _13369_/CLK _13272_/D vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12223_ _12224_/A _12224_/B vssd1 vssd1 vccd1 vccd1 _12284_/A sky130_fd_sc_hd__or2_1
XANTENNA__10187__B1 _10049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12154_ _12103_/A _12103_/B _12102_/A vssd1 vssd1 vccd1 vccd1 _12175_/A sky130_fd_sc_hd__a21o_1
XANTENNA__11923__A1 _12631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07052__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11105_ _11106_/A _11106_/B vssd1 vssd1 vccd1 vccd1 _11105_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_75_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12085_ _12084_/B _12085_/B vssd1 vssd1 vccd1 vccd1 _12086_/B sky130_fd_sc_hd__nand2b_1
X_11036_ _11650_/B _11143_/B hold270/A vssd1 vssd1 vccd1 vccd1 _11036_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12987_ _13001_/A hold212/X vssd1 vssd1 vccd1 vccd1 _13303_/D sky130_fd_sc_hd__and2_1
XANTENNA__08304__B1 _09770_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11938_ _11939_/A _11939_/B vssd1 vssd1 vccd1 vccd1 _12030_/B sky130_fd_sc_hd__or2_1
X_11869_ _11870_/A _11870_/B vssd1 vssd1 vccd1 vccd1 _11952_/B sky130_fd_sc_hd__and2b_1
XANTENNA__06654__A _06723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09804__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09030__A _09031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07060_ _07102_/A _07102_/B vssd1 vssd1 vccd1 vccd1 _07104_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_125_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11914__A1 _12421_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07043__B1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07485__A _09834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11390__A2 _07157_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07594__A1 _12224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09701_ _09701_/A _09701_/B vssd1 vssd1 vccd1 vccd1 _09703_/B sky130_fd_sc_hd__xnor2_2
X_07962_ _07962_/A _07962_/B vssd1 vssd1 vccd1 vccd1 _08061_/B sky130_fd_sc_hd__xor2_1
X_06913_ reg1_idx[0] reg1_idx[1] reg1_idx[4] vssd1 vssd1 vccd1 vccd1 _06915_/C sky130_fd_sc_hd__and3_1
XANTENNA__11678__B1 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07893_ _07148_/Y _07959_/B fanout29/X _07959_/A vssd1 vssd1 vccd1 vccd1 _07894_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07346__A1 _09934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06844_ _11022_/A _06842_/X _06843_/X vssd1 vssd1 vccd1 vccd1 _06844_/Y sky130_fd_sc_hd__a21oi_1
X_09632_ _09836_/A _09632_/B vssd1 vssd1 vccd1 vccd1 _09633_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07346__B2 _07830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09563_ _09159_/X _09163_/X _09725_/S vssd1 vssd1 vccd1 vccd1 _09563_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06775_ _06773_/Y _06775_/B vssd1 vssd1 vccd1 vccd1 _10291_/A sky130_fd_sc_hd__nand2b_2
X_08514_ _10243_/A _08514_/B vssd1 vssd1 vccd1 vccd1 _08552_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09494_ _09494_/A _09494_/B vssd1 vssd1 vccd1 vccd1 _09495_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_38_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07649__A2 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08445_ _08598_/B _08561_/A2 _08561_/B1 _08538_/A1 vssd1 vssd1 vccd1 vccd1 _08446_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08376_ _08424_/A _08424_/B vssd1 vssd1 vccd1 vccd1 _08425_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_18_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07327_ _09944_/A _07327_/B vssd1 vssd1 vccd1 vccd1 _07387_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07258_ _07255_/A _07255_/B _10623_/A vssd1 vssd1 vccd1 vccd1 _07258_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09875__A _12404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09594__B _09596_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07189_ _09667_/A _07200_/C vssd1 vssd1 vccd1 vccd1 _07189_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_14_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09326__A2 _08877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07337__A1 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12910_ hold154/X hold245/X vssd1 vssd1 vccd1 vccd1 _12910_/X sky130_fd_sc_hd__and2b_1
XANTENNA__07337__B2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12841_ _07256_/Y _12863_/A2 hold37/X _13210_/A vssd1 vssd1 vccd1 vccd1 _13281_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09115__A _09341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _12780_/A _12772_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[26] sky130_fd_sc_hd__xnor2_4
XANTENNA__08837__B2 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08837__A1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11723_ _11723_/A _11723_/B vssd1 vssd1 vccd1 vccd1 _11723_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__11380__A _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11654_ _07078_/A _09257_/S _11653_/X vssd1 vssd1 vccd1 vccd1 _11654_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10605_ _10606_/A _10606_/B vssd1 vssd1 vccd1 vccd1 _10605_/X sky130_fd_sc_hd__and2_1
XFILLER_0_83_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout70 _09936_/A vssd1 vssd1 vccd1 vccd1 _12157_/A sky130_fd_sc_hd__buf_4
Xfanout92 _09779_/A vssd1 vssd1 vccd1 vccd1 _12224_/A sky130_fd_sc_hd__buf_8
Xfanout81 _07261_/Y vssd1 vssd1 vccd1 vccd1 _11198_/A sky130_fd_sc_hd__clkbuf_8
X_11585_ _11586_/A _11586_/B vssd1 vssd1 vccd1 vccd1 _11692_/B sky130_fd_sc_hd__or2_2
XFILLER_0_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13324_ _13392_/CLK hold226/X vssd1 vssd1 vccd1 vccd1 hold224/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10536_ _10536_/A _10536_/B vssd1 vssd1 vccd1 vccd1 _10538_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_51_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12149__A1 _12365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10724__A _11844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10467_ _10468_/A _10468_/B _10468_/C vssd1 vssd1 vccd1 vccd1 _10645_/A sky130_fd_sc_hd__a21oi_1
X_13255_ hold167/X hold140/X hold127/X vssd1 vssd1 vccd1 vccd1 hold306/A sky130_fd_sc_hd__a21o_1
X_12206_ _12206_/A _12206_/B vssd1 vssd1 vccd1 vccd1 _12211_/C sky130_fd_sc_hd__nor2_1
X_13186_ hold246/X _13223_/A2 _13185_/X _13223_/B2 vssd1 vssd1 vccd1 vccd1 hold247/A
+ sky130_fd_sc_hd__a22o_1
X_10398_ _10398_/A _10398_/B vssd1 vssd1 vccd1 vccd1 _10411_/A sky130_fd_sc_hd__xnor2_1
X_12137_ _12449_/B1 _12199_/B hold276/A vssd1 vssd1 vccd1 vccd1 _12139_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12068_ hold254/A _12068_/B vssd1 vssd1 vccd1 vccd1 _12136_/B sky130_fd_sc_hd__or2_1
XANTENNA__07328__A1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09317__A2 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11019_ _06897_/D _10909_/Y _10927_/S vssd1 vssd1 vccd1 vccd1 _11019_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__07328__B2 _09661_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08864__A _09947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08230_ _08230_/A _08230_/B vssd1 vssd1 vccd1 vccd1 _08231_/B sky130_fd_sc_hd__and2_1
XFILLER_0_27_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10938__A2 _07362_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09253__B2 _12379_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08161_ _08158_/A _08158_/B _08231_/A vssd1 vssd1 vccd1 vccd1 _08186_/A sky130_fd_sc_hd__a21oi_2
X_07112_ reg1_val[22] _07112_/B vssd1 vssd1 vccd1 vccd1 _07140_/C sky130_fd_sc_hd__or2_1
XFILLER_0_42_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08092_ _08575_/A _08092_/B vssd1 vssd1 vccd1 vccd1 _08122_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07043_ fanout65/X _08657_/B fanout59/X _08649_/A2 vssd1 vssd1 vccd1 vccd1 _07044_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09005__A1 _10725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09005__B2 _07232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout109_A _07237_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11899__B1 _09225_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08104__A _08334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10571__B1 _12416_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08994_ _09677_/A _07362_/B fanout16/X _07172_/Y vssd1 vssd1 vccd1 vccd1 _08995_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07945_ _08011_/B _08011_/A vssd1 vssd1 vccd1 vccd1 _07948_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__12863__A2 _12863_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11666__A3 _08974_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09615_ fanout42/X _10337_/A _07238_/Y _07417_/B vssd1 vssd1 vccd1 vccd1 _09616_/B
+ sky130_fd_sc_hd__a22o_1
X_07876_ _07876_/A _07876_/B vssd1 vssd1 vccd1 vccd1 _07877_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_92_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06827_ reg1_val[5] _06827_/B vssd1 vssd1 vccd1 vccd1 _06827_/Y sky130_fd_sc_hd__nand2_1
X_06758_ reg1_val[10] _07233_/A vssd1 vssd1 vccd1 vccd1 _10688_/S sky130_fd_sc_hd__and2_1
X_09546_ _09548_/A _09548_/B vssd1 vssd1 vccd1 vccd1 _09546_/X sky130_fd_sc_hd__or2_2
X_09477_ _09475_/X _09477_/B vssd1 vssd1 vccd1 vccd1 _09478_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_93_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06689_ reg2_val[20] _06810_/B _06724_/B1 _06688_/Y vssd1 vssd1 vccd1 vccd1 _07016_/A
+ sky130_fd_sc_hd__o2bb2a_4
X_08428_ _08438_/A _08438_/B _08414_/Y vssd1 vssd1 vccd1 vccd1 _08435_/B sky130_fd_sc_hd__o21a_1
XANTENNA__12379__A1 _09221_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12379__B2 _12379_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10929__A2 _12422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08359_ _08402_/A _08402_/B vssd1 vssd1 vccd1 vccd1 _08690_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09795__A2 _10476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11370_ _12365_/A _11344_/X _11345_/Y _11369_/X _11343_/Y vssd1 vssd1 vccd1 vccd1
+ _11370_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10321_ _10321_/A _10321_/B _10321_/C vssd1 vssd1 vccd1 vccd1 _10324_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_34_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06741__B _11038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13040_ hold119/X _13094_/A2 _13101_/A2 hold125/X _13039_/A vssd1 vssd1 vccd1 vccd1
+ hold126/A sky130_fd_sc_hd__o221a_1
X_10252_ _10383_/A _10251_/C _10097_/A vssd1 vssd1 vccd1 vccd1 _10253_/C sky130_fd_sc_hd__a21bo_1
X_10183_ _10149_/Y _10152_/X _10182_/Y _11752_/S vssd1 vssd1 vccd1 vccd1 _10183_/X
+ sky130_fd_sc_hd__a31o_1
Xfanout282 _13142_/A vssd1 vssd1 vccd1 vccd1 _13246_/A sky130_fd_sc_hd__buf_4
Xfanout271 _06606_/X vssd1 vssd1 vccd1 vccd1 _06927_/A sky130_fd_sc_hd__clkbuf_4
Xfanout260 hold191/X vssd1 vssd1 vccd1 vccd1 _13248_/A2 sky130_fd_sc_hd__buf_4
XANTENNA__08507__B1 _07282_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09180__A0 _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout293 reg1_val[0] vssd1 vssd1 vccd1 vccd1 _09218_/A sky130_fd_sc_hd__buf_4
XANTENNA__12067__B1 _11648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12824_ hold30/X _12826_/B vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__or2_1
XFILLER_0_84_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12755_ reg1_val[23] _12755_/B vssd1 vssd1 vccd1 vccd1 _12760_/D sky130_fd_sc_hd__xnor2_4
XFILLER_0_29_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11706_ _11797_/B _11706_/B vssd1 vssd1 vccd1 vccd1 _11709_/A sky130_fd_sc_hd__nand2_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10093__A2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12686_ _12691_/B _12693_/A vssd1 vssd1 vccd1 vccd1 _12687_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_25_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11637_ _11637_/A _11637_/B _11637_/C vssd1 vssd1 vccd1 vccd1 _11657_/D sky130_fd_sc_hd__or3_1
XANTENNA__09235__A1 _12365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11568_ fanout58/X fanout23/X fanout15/X _11868_/A vssd1 vssd1 vccd1 vccd1 _11569_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_64_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10519_ _10519_/A _10519_/B _10519_/C vssd1 vssd1 vccd1 vccd1 _10521_/A sky130_fd_sc_hd__and3_1
X_13307_ _13309_/CLK _13307_/D vssd1 vssd1 vccd1 vccd1 hold213/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07797__B2 _07148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07797__A1 _07173_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08994__B1 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11499_ _12096_/A _11499_/B vssd1 vssd1 vccd1 vccd1 _11500_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06651__B _06998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13238_ _13238_/A _13238_/B vssd1 vssd1 vccd1 vccd1 _13239_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_110_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13169_ _13169_/A _13169_/B vssd1 vssd1 vccd1 vccd1 _13169_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_383 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13098__A2 _06577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07730_ _07731_/A _07731_/B vssd1 vssd1 vccd1 vccd1 _07730_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12845__A2 _12863_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10305__B1 _12416_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07661_ _07370_/A _07369_/B _07367_/Y vssd1 vssd1 vccd1 vccd1 _07671_/A sky130_fd_sc_hd__a21o_1
X_06612_ instruction[1] instruction[2] instruction[25] pred_val vssd1 vssd1 vccd1
+ vccd1 _06612_/X sky130_fd_sc_hd__o211a_1
X_09400_ _09201_/X _09203_/X _09403_/S vssd1 vssd1 vccd1 vccd1 _09400_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12058__B1 _10788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07592_ _07592_/A _07592_/B vssd1 vssd1 vccd1 vccd1 _07660_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__12828__B _12870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09331_ _09331_/A _09331_/B vssd1 vssd1 vccd1 vccd1 _09332_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10629__A _11179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13005__A _13019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09262_ _09144_/A _09144_/B _09142_/X vssd1 vssd1 vccd1 vccd1 _09371_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__13022__A2 _13171_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09193_ reg1_val[2] reg1_val[29] _09211_/S vssd1 vssd1 vccd1 vccd1 _09193_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08213_ _08213_/A _08213_/B vssd1 vssd1 vccd1 vccd1 _08224_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_7_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08144_ _09770_/B2 _08484_/B _09479_/B1 _09940_/B2 vssd1 vssd1 vccd1 vccd1 _08145_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_70_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08075_ _08075_/A _08075_/B vssd1 vssd1 vccd1 vccd1 _08076_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_113_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07026_ _09672_/A _07029_/B vssd1 vssd1 vccd1 vccd1 _07030_/A sky130_fd_sc_hd__and2_1
XFILLER_0_87_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10544__B1 _10415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold13 hold75/X vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ _09672_/A _08977_/B vssd1 vssd1 vccd1 vccd1 _08981_/A sky130_fd_sc_hd__xnor2_4
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ _07924_/A _07924_/B _07972_/A vssd1 vssd1 vccd1 vccd1 _08003_/A sky130_fd_sc_hd__o21bai_2
X_07859_ _08334_/A _07859_/B vssd1 vssd1 vccd1 vccd1 _07883_/B sky130_fd_sc_hd__xnor2_1
X_10870_ _10737_/A _10737_/B _10733_/X vssd1 vssd1 vccd1 vccd1 _10872_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__07712__B2 _08457_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07712__A1 _10338_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout41_A fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09529_ _09529_/A _09529_/B vssd1 vssd1 vccd1 vccd1 _09530_/B sky130_fd_sc_hd__nor2_1
XANTENNA__06736__B _07270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10539__A _10539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12540_ _12546_/B _12540_/B vssd1 vssd1 vccd1 vccd1 new_PC[11] sky130_fd_sc_hd__and2_4
XFILLER_0_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07476__B1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12471_ reg1_val[2] curr_PC[2] _12471_/S vssd1 vssd1 vccd1 vccd1 _12473_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_47_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11422_ _11422_/A _11422_/B vssd1 vssd1 vccd1 vccd1 _11424_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12221__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11575__A2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08976__B1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11353_ _11351_/Y _11353_/B vssd1 vssd1 vccd1 vccd1 _11354_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_61_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08440__A2 _08576_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11284_ _11284_/A _11284_/B vssd1 vssd1 vccd1 vccd1 _11288_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10304_ _09425_/C _10569_/C hold281/A vssd1 vssd1 vccd1 vccd1 _10304_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13023_ _13249_/A hold207/X vssd1 vssd1 vccd1 vccd1 _13321_/D sky130_fd_sc_hd__and2_1
X_10235_ _12224_/A _10235_/B vssd1 vssd1 vccd1 vccd1 _10237_/B sky130_fd_sc_hd__xor2_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07583__A _09341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10166_ hold196/A hold300/A _10166_/C vssd1 vssd1 vccd1 vccd1 _10300_/B sky130_fd_sc_hd__or3_1
XANTENNA__09940__A2 _08877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12288__B1 _11844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12827__A2 _13101_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10097_ _10097_/A _10097_/B vssd1 vssd1 vccd1 vccd1 _10100_/A sky130_fd_sc_hd__and2_1
XFILLER_0_89_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07164__C1 _12438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12807_ _12428_/B _12871_/A2 hold10/X _13246_/A vssd1 vssd1 vccd1 vccd1 _13264_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__06927__A _06927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10999_ _11000_/A _11000_/B vssd1 vssd1 vccd1 vccd1 _11117_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13252__A2 _13254_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11263__B2 _12379_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12460__A0 _09218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12738_ reg1_val[20] _12755_/B vssd1 vssd1 vccd1 vccd1 _12760_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13004__A2 _13171_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12669_ reg1_val[6] _12670_/B vssd1 vssd1 vccd1 vccd1 _12671_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12212__B1 _11892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09880_ _11029_/S _09879_/Y _09251_/A vssd1 vssd1 vccd1 vccd1 _09880_/Y sky130_fd_sc_hd__a21boi_4
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08900_ _08900_/A _08900_/B vssd1 vssd1 vccd1 vccd1 _08912_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_57_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _07615_/A _07615_/B _07613_/X vssd1 vssd1 vccd1 vccd1 _08833_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__06745__A2 _06723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _11444_/B _11444_/C vssd1 vssd1 vccd1 vccd1 _11538_/B sky130_fd_sc_hd__nand2_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07713_ _10207_/A _07713_/B vssd1 vssd1 vccd1 vccd1 _07717_/A sky130_fd_sc_hd__xnor2_2
X_08693_ _08779_/B _08769_/A _08766_/A _08761_/B vssd1 vssd1 vccd1 vccd1 _08693_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA_fanout176_A _10159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07644_ _07644_/A _07644_/B vssd1 vssd1 vccd1 vccd1 _07645_/B sky130_fd_sc_hd__or2_1
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07575_ _10871_/A fanout33/X fanout72/X _08199_/B vssd1 vssd1 vccd1 vccd1 _07576_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_75_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10057__A2 fanout86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09314_ _09315_/A _09315_/B vssd1 vssd1 vccd1 vccd1 _09316_/A sky130_fd_sc_hd__or2_1
XFILLER_0_118_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09245_ _09728_/S _09250_/B _09244_/X vssd1 vssd1 vccd1 vccd1 _09246_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09176_ reg1_val[12] reg1_val[19] _09180_/S vssd1 vssd1 vccd1 vccd1 _09176_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10094__A _11582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08127_ _08664_/A _08127_/B vssd1 vssd1 vccd1 vccd1 _08198_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08058_ _08028_/X _08056_/B _08057_/Y vssd1 vssd1 vccd1 vccd1 _08070_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_31_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07009_ _07604_/A _07010_/B vssd1 vssd1 vccd1 vccd1 _07011_/A sky130_fd_sc_hd__or2_2
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout89_A _11284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12513__S _12520_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10020_ _11246_/S _10020_/B vssd1 vssd1 vccd1 vccd1 _10020_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12809__A2 _12820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11971_ _11622_/X _11967_/Y _11968_/Y _11232_/B _11970_/X vssd1 vssd1 vccd1 vccd1
+ _11972_/B sky130_fd_sc_hd__a221o_2
XFILLER_0_86_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10922_ _11990_/A1 _11032_/B hold198/A vssd1 vssd1 vccd1 vccd1 _10922_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_85_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10853_ _10854_/A _10854_/B vssd1 vssd1 vccd1 vccd1 _10980_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10784_ _11008_/A _10784_/B vssd1 vssd1 vccd1 vccd1 _11050_/B sky130_fd_sc_hd__xnor2_4
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07449__B1 _10974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12523_ _12532_/A _12523_/B vssd1 vssd1 vccd1 vccd1 _12525_/C sky130_fd_sc_hd__nand2_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07578__A _09836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12454_ _06963_/B _11829_/B _09252_/Y _09221_/Y _12453_/X vssd1 vssd1 vccd1 vccd1
+ _12454_/X sky130_fd_sc_hd__a221o_1
XANTENNA__08949__B1 _10240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11405_ _12336_/A _11405_/B vssd1 vssd1 vccd1 vccd1 _11407_/A sky130_fd_sc_hd__xnor2_1
X_12385_ fanout7/X _12385_/B vssd1 vssd1 vccd1 vccd1 _12385_/X sky130_fd_sc_hd__or2_1
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11336_ _11119_/X _11528_/A _11335_/X vssd1 vssd1 vccd1 vccd1 _11716_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__07621__B1 _10245_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10732__A _11770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13006_ hold182/X _13171_/B2 _13209_/A2 hold204/X vssd1 vssd1 vccd1 vccd1 hold205/A
+ sky130_fd_sc_hd__a22o_1
X_11267_ curr_PC[15] _11268_/B vssd1 vssd1 vccd1 vccd1 _11267_/X sky130_fd_sc_hd__or2_1
X_11198_ _11198_/A _12087_/B vssd1 vssd1 vccd1 vccd1 _11199_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11181__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10218_ _10218_/A _10218_/B vssd1 vssd1 vccd1 vccd1 _10220_/B sky130_fd_sc_hd__xor2_1
X_10149_ _10049_/Y _10147_/A _10148_/Y vssd1 vssd1 vccd1 vccd1 _10149_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10692__C1 _12376_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07360_ _12224_/A _07361_/B vssd1 vssd1 vccd1 vccd1 _07360_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_57_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08101__A1 _10221_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08101__B2 _09770_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07291_ _07292_/B _07374_/A _07292_/A vssd1 vssd1 vccd1 vccd1 _07663_/A sky130_fd_sc_hd__o21a_1
X_09030_ _09031_/A _09031_/B vssd1 vssd1 vccd1 vccd1 _09030_/X sky130_fd_sc_hd__and2_1
XFILLER_0_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold302 hold302/A vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09601__A1 _07172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09932_ _09930_/X _09932_/B vssd1 vssd1 vccd1 vccd1 _09933_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_7_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13161__B2 _13171_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09904__A2 _09880_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09863_ _09863_/A _10004_/A _10137_/A _10137_/B vssd1 vssd1 vccd1 vccd1 _09863_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__08112__A _09404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _09794_/A _09794_/B vssd1 vssd1 vccd1 vccd1 _09797_/A sky130_fd_sc_hd__xnor2_1
X_08814_ _07628_/A _07627_/Y _07625_/X vssd1 vssd1 vccd1 vccd1 _08827_/B sky130_fd_sc_hd__a21o_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08745_ _08745_/A _08745_/B vssd1 vssd1 vccd1 vccd1 _08745_/X sky130_fd_sc_hd__xor2_1
XANTENNA__07391__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11475__A1 _11476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08676_ _08677_/A _08677_/B _08727_/A vssd1 vssd1 vccd1 vccd1 _08678_/C sky130_fd_sc_hd__a21o_1
XANTENNA__08340__A1 _08657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07627_ _07628_/B vssd1 vssd1 vccd1 vccd1 _07627_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08340__B2 _08649_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07158__A_N _12224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07558_ _07558_/A _07741_/A vssd1 vssd1 vccd1 vccd1 _07681_/A sky130_fd_sc_hd__or2_1
XFILLER_0_119_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07489_ _09922_/A _07489_/B vssd1 vssd1 vccd1 vccd1 _07489_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_106_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09228_ _09239_/A _09228_/B vssd1 vssd1 vccd1 vccd1 _09228_/X sky130_fd_sc_hd__or2_4
XFILLER_0_51_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07851__B1 fanout72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09159_ _09157_/X _09158_/X _09383_/S vssd1 vssd1 vccd1 vccd1 _09159_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12170_ _12233_/D _12170_/B vssd1 vssd1 vccd1 vccd1 _12172_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07603__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11648__A _11648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11121_ _10899_/Y _11334_/A _11119_/X vssd1 vssd1 vccd1 vccd1 _11121_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_101_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11052_ _11893_/A _11052_/B vssd1 vssd1 vccd1 vccd1 _11052_/X sky130_fd_sc_hd__or2_1
X_10003_ _09709_/Y _10278_/A _10001_/Y vssd1 vssd1 vccd1 vccd1 _10003_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07382__A2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11383__A _11582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12479__A _12655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09659__A1 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09659__B2 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11954_ _11955_/A _11955_/B vssd1 vssd1 vccd1 vccd1 _12036_/B sky130_fd_sc_hd__nand2b_1
X_11885_ _11885_/A _12043_/A vssd1 vssd1 vccd1 vccd1 _11886_/A sky130_fd_sc_hd__and2_1
X_10905_ _10824_/X _11050_/C _09150_/X vssd1 vssd1 vccd1 vccd1 _10905_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10836_ _10836_/A _10836_/B vssd1 vssd1 vccd1 vccd1 _10838_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10767_ _10643_/A _10643_/B _10646_/A vssd1 vssd1 vccd1 vccd1 _10768_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_82_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06924__B _06926_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12506_ reg1_val[7] curr_PC[7] _12520_/S vssd1 vssd1 vccd1 vccd1 _12508_/B sky130_fd_sc_hd__mux2_1
X_10698_ _10665_/Y _10666_/X _10669_/Y _10788_/A _10697_/X vssd1 vssd1 vccd1 vccd1
+ _10698_/X sky130_fd_sc_hd__o221a_1
X_12437_ _12427_/X _12435_/Y _12436_/Y vssd1 vssd1 vccd1 vccd1 _12437_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10729__B1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12368_ _12444_/C _12367_/Y _12444_/B vssd1 vssd1 vccd1 vccd1 _12368_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_50_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11319_ _11319_/A _11319_/B vssd1 vssd1 vccd1 vccd1 _11320_/B sky130_fd_sc_hd__nor2_1
X_12299_ _12299_/A _12430_/A vssd1 vssd1 vccd1 vccd1 _12300_/C sky130_fd_sc_hd__or2_1
X_06860_ _06860_/A _06860_/B vssd1 vssd1 vccd1 vccd1 _06860_/X sky130_fd_sc_hd__or2_1
X_06791_ reg2_val[4] _06810_/B vssd1 vssd1 vccd1 vccd1 _06791_/X sky130_fd_sc_hd__and2_2
X_08530_ _08641_/B _08561_/B1 _08576_/A2 _08627_/A2 vssd1 vssd1 vccd1 vccd1 _08531_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08461_ _08485_/A _08485_/B _08497_/B _08460_/B _08460_/A vssd1 vssd1 vccd1 vccd1
+ _08469_/A sky130_fd_sc_hd__o32a_1
XANTENNA__11209__A1 _11093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07412_ _07433_/A _07433_/B vssd1 vssd1 vccd1 vccd1 _07428_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12836__B _12862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08392_ _08392_/A _08392_/B vssd1 vssd1 vccd1 vccd1 _08394_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_128_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07343_ _07343_/A _07343_/B vssd1 vssd1 vccd1 vccd1 _07356_/A sky130_fd_sc_hd__xnor2_2
X_07274_ _11038_/A _07274_/B vssd1 vssd1 vccd1 vccd1 _07274_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08107__A _10207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09013_ _09014_/B _09014_/A vssd1 vssd1 vccd1 vccd1 _09013_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_79_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold110 hold110/A vssd1 vssd1 vccd1 vccd1 hold110/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08389__A1 _08540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08389__B2 _08515_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold121 hold121/A vssd1 vssd1 vccd1 vccd1 hold121/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 hold143/A vssd1 vssd1 vccd1 vccd1 hold143/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 hold132/A vssd1 vssd1 vccd1 vccd1 hold132/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold176 hold176/A vssd1 vssd1 vccd1 vccd1 hold176/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 hold154/A vssd1 vssd1 vccd1 vccd1 hold154/X sky130_fd_sc_hd__buf_1
Xhold165 hold165/A vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 hold198/A vssd1 vssd1 vccd1 vccd1 hold198/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 hold187/A vssd1 vssd1 vccd1 vccd1 hold187/X sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ _12224_/A _09915_/B vssd1 vssd1 vccd1 vccd1 _09919_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_0_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09338__B1 _10599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11145__B1 _12376_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09889__A1 _12322_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09846_ _09844_/Y _09846_/B vssd1 vssd1 vccd1 vccd1 _09847_/B sky130_fd_sc_hd__and2b_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08561__A1 _08657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06989_ _06987_/A _06987_/B _07046_/C _07094_/B vssd1 vssd1 vccd1 vccd1 _06991_/B
+ sky130_fd_sc_hd__a31o_2
X_09777_ _09780_/A vssd1 vssd1 vccd1 vccd1 _09777_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08561__B2 _08649_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11448__A1 _11813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08728_ _10420_/B _10420_/C vssd1 vssd1 vccd1 vccd1 _10552_/B sky130_fd_sc_hd__and2_1
XFILLER_0_96_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _08661_/A _08659_/B vssd1 vssd1 vccd1 vccd1 _08666_/A sky130_fd_sc_hd__and2b_1
XANTENNA__11931__A _12093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _11868_/A fanout10/X fanout5/X fanout62/X vssd1 vssd1 vccd1 vccd1 _11764_/C
+ sky130_fd_sc_hd__o22a_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10959__B1 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10621_ _10504_/A _10503_/B _10503_/A vssd1 vssd1 vccd1 vccd1 _10636_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__06744__B _06810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08616__A2 _07166_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13340_ _13358_/CLK _13340_/D vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10552_ _11630_/A _10552_/B _10552_/C vssd1 vssd1 vccd1 vccd1 _10552_/X sky130_fd_sc_hd__or3_1
XFILLER_0_24_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13271_ _13369_/CLK _13271_/D vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10483_ _10366_/A _10366_/B _10363_/A vssd1 vssd1 vccd1 vccd1 _10485_/B sky130_fd_sc_hd__a21o_1
X_12222_ _12335_/B _12222_/B vssd1 vssd1 vccd1 vccd1 _12224_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12153_ _12151_/Y _12152_/X _12631_/S _12150_/X vssd1 vssd1 vccd1 vccd1 dest_val[25]
+ sky130_fd_sc_hd__a2bb2o_4
XANTENNA__07052__B2 _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07052__A1 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11104_ _10975_/A _10975_/B _10973_/A vssd1 vssd1 vccd1 vccd1 _11106_/B sky130_fd_sc_hd__a21o_1
X_12084_ _12085_/B _12084_/B vssd1 vssd1 vccd1 vccd1 _12086_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_20_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11035_ hold285/A _11035_/B vssd1 vssd1 vccd1 vccd1 _11143_/B sky130_fd_sc_hd__or2_1
XFILLER_0_99_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11439__A1 _10548_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12986_ hold196/X _13000_/A2 _13257_/A2 hold211/X vssd1 vssd1 vccd1 vccd1 hold212/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08304__B2 _08538_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08304__A1 _08598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11937_ _12030_/A _11937_/B vssd1 vssd1 vccd1 vccd1 _11939_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11841__A _11841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11868_ _11868_/A _12335_/B vssd1 vssd1 vccd1 vccd1 _11870_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_86_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10457__A _11179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11799_ _11799_/A _11884_/A vssd1 vssd1 vccd1 vccd1 _11966_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_55_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09804__A1 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10819_ curr_PC[11] _10934_/C vssd1 vssd1 vccd1 vccd1 _10819_/X sky130_fd_sc_hd__or2_1
XANTENNA__09311__A _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06654__B _12685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09804__B2 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07043__B2 _08649_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07043__A1 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07961_ _07962_/B _07962_/A vssd1 vssd1 vccd1 vccd1 _07966_/A sky130_fd_sc_hd__and2b_1
X_06912_ _06944_/B dest_pred_val _12218_/A vssd1 vssd1 vccd1 vccd1 take_branch sky130_fd_sc_hd__a21o_4
X_09700_ _09701_/B _09701_/A vssd1 vssd1 vccd1 vccd1 _09700_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__11678__A1 _12233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07892_ _10092_/A _07892_/B vssd1 vssd1 vccd1 vccd1 _07896_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07346__A2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06843_ _11038_/A reg1_val[13] vssd1 vssd1 vccd1 vccd1 _06843_/X sky130_fd_sc_hd__and2b_1
X_09631_ _07959_/B _07262_/X _07269_/Y fanout29/X vssd1 vssd1 vccd1 vccd1 _09632_/B
+ sky130_fd_sc_hd__a22o_1
X_09562_ _09562_/A vssd1 vssd1 vccd1 vccd1 _09562_/Y sky130_fd_sc_hd__inv_2
X_06774_ reg1_val[7] _07222_/A vssd1 vssd1 vccd1 vccd1 _06775_/B sky130_fd_sc_hd__nand2_1
X_08513_ _08598_/B _08576_/A2 _09472_/A _08538_/A1 vssd1 vssd1 vccd1 vccd1 _08514_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout256_A _13000_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09493_ _09494_/A _09494_/B vssd1 vssd1 vccd1 vccd1 _09495_/A sky130_fd_sc_hd__or2_1
XFILLER_0_77_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08444_ _08447_/A _08447_/B vssd1 vssd1 vccd1 vccd1 _08444_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09221__A _12359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08375_ _08375_/A _08375_/B vssd1 vssd1 vccd1 vccd1 _08424_/B sky130_fd_sc_hd__xnor2_2
X_07326_ fanout61/X _09943_/B2 fanout53/X _09650_/A vssd1 vssd1 vccd1 vccd1 _07327_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07257_ _07094_/A _07093_/X _07094_/Y _06979_/Y vssd1 vssd1 vccd1 vccd1 _07257_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07188_ reg1_val[16] _07188_/B vssd1 vssd1 vccd1 vccd1 _07200_/C sky130_fd_sc_hd__xnor2_2
XANTENNA__11198__A _11198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07034__A1 _07014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06793__B1 _06791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07337__A2 _10245_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09829_ _09830_/A _09830_/B vssd1 vssd1 vccd1 vccd1 _09829_/Y sky130_fd_sc_hd__nor2_1
X_12840_ hold36/X _12862_/B vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__or2_1
XANTENNA__06739__B _06810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _12790_/B _07357_/C _12780_/B vssd1 vssd1 vccd1 vccd1 _12772_/B sky130_fd_sc_hd__a21bo_2
XANTENNA__08837__A2 _09943_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08298__B1 _10338_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _11630_/B _11630_/C _11630_/A vssd1 vssd1 vccd1 vccd1 _11723_/B sky130_fd_sc_hd__a21o_1
X_11653_ _12421_/A1 _11652_/X _06707_/B vssd1 vssd1 vccd1 vccd1 _11653_/X sky130_fd_sc_hd__a21o_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10604_ _11284_/A _10604_/B vssd1 vssd1 vccd1 vccd1 _10606_/B sky130_fd_sc_hd__xnor2_1
Xfanout60 _07033_/X vssd1 vssd1 vccd1 vccd1 _12009_/A sky130_fd_sc_hd__buf_4
Xfanout82 _10476_/A vssd1 vssd1 vccd1 vccd1 fanout82/X sky130_fd_sc_hd__buf_8
Xfanout71 _07587_/Y vssd1 vssd1 vccd1 vccd1 _09936_/A sky130_fd_sc_hd__buf_6
XFILLER_0_36_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11584_ _11584_/A _11584_/B vssd1 vssd1 vccd1 vccd1 _11586_/B sky130_fd_sc_hd__xnor2_1
X_13323_ _13392_/CLK hold231/X vssd1 vssd1 vccd1 vccd1 hold229/A sky130_fd_sc_hd__dfxtp_1
Xfanout93 _09779_/A vssd1 vssd1 vccd1 vccd1 _12096_/A sky130_fd_sc_hd__buf_8
XFILLER_0_52_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10535_ _10536_/B _10536_/A vssd1 vssd1 vccd1 vccd1 _10655_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_52_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10466_ _10618_/B _10466_/B vssd1 vssd1 vccd1 vccd1 _10468_/C sky130_fd_sc_hd__nand2_1
X_13254_ hold127/X _13254_/A2 _12798_/Y _06577_/A vssd1 vssd1 vccd1 vccd1 _13256_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13185_ hold292/A _13184_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13185_/X sky130_fd_sc_hd__mux2_1
X_12205_ hold229/A _12447_/B1 _12266_/B _12205_/B1 vssd1 vssd1 vccd1 vccd1 _12206_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12136_ hold278/A _12136_/B vssd1 vssd1 vccd1 vccd1 _12199_/B sky130_fd_sc_hd__or2_1
X_10397_ _10397_/A _10397_/B vssd1 vssd1 vccd1 vccd1 _10398_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09970__B1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06784__B1 _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10580__A1 _12471_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12067_ hold206/A _12322_/A1 _12140_/B _11648_/A vssd1 vssd1 vccd1 vccd1 _12067_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11018_ _11809_/A _08744_/X _08745_/X _10788_/A vssd1 vssd1 vccd1 vccd1 _11018_/Y
+ sky130_fd_sc_hd__a31oi_1
XANTENNA__09306__A _09672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07328__A2 _10245_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12969_ _13238_/A _13239_/A _13238_/B vssd1 vssd1 vccd1 vccd1 _13243_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_75_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11571__A _12093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11832__B2 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11832__A1 _10159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08160_ _08230_/A _08230_/B vssd1 vssd1 vccd1 vccd1 _08231_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_83_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07111_ reg1_val[20] reg1_val[21] vssd1 vssd1 vccd1 vccd1 _07112_/B sky130_fd_sc_hd__or2_1
XANTENNA__09253__A2 _09221_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12606__S _12631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08091_ _08657_/B fanout80/X fanout76/X _08649_/A2 vssd1 vssd1 vccd1 vccd1 _08092_/B
+ sky130_fd_sc_hd__o22a_1
X_07042_ _07404_/A _07404_/B _07023_/X vssd1 vssd1 vccd1 vccd1 _07102_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_2_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09005__A2 _07959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08993_ _08867_/A _08867_/B _08865_/X vssd1 vssd1 vccd1 vccd1 _08997_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07944_ _07944_/A _07944_/B vssd1 vssd1 vccd1 vccd1 _08011_/B sky130_fd_sc_hd__xnor2_2
X_07875_ _07946_/A _07946_/B _07946_/C vssd1 vssd1 vccd1 vccd1 _07947_/A sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_4_2_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06826_ _06898_/C _06824_/X _06825_/X vssd1 vssd1 vccd1 vccd1 _06826_/Y sky130_fd_sc_hd__a21oi_1
X_09614_ _09614_/A _09614_/B vssd1 vssd1 vccd1 vccd1 _09618_/B sky130_fd_sc_hd__xor2_1
XANTENNA__12076__A1 _06946_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06757_ reg1_val[10] _07233_/A vssd1 vssd1 vccd1 vccd1 _06759_/A sky130_fd_sc_hd__nor2_1
X_09545_ _09545_/A _09545_/B vssd1 vssd1 vccd1 vccd1 _09548_/B sky130_fd_sc_hd__xnor2_4
X_06688_ _06703_/A _12665_/B vssd1 vssd1 vccd1 vccd1 _06688_/Y sky130_fd_sc_hd__nor2_1
X_09476_ _09476_/A _09476_/B _09476_/C vssd1 vssd1 vccd1 vccd1 _09477_/B sky130_fd_sc_hd__or3_1
XFILLER_0_19_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08427_ _08427_/A _08427_/B vssd1 vssd1 vccd1 vccd1 _08438_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08358_ _08358_/A _08358_/B vssd1 vssd1 vccd1 vccd1 _08402_/B sky130_fd_sc_hd__xor2_1
XANTENNA__08988__D1 _12795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09795__A3 _10476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08289_ _09404_/S _08289_/B vssd1 vssd1 vccd1 vccd1 _08290_/B sky130_fd_sc_hd__nor2_2
X_07309_ _07310_/A _07310_/B vssd1 vssd1 vccd1 vccd1 _07663_/B sky130_fd_sc_hd__and2_1
XFILLER_0_116_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10320_ _10821_/A _10317_/X _10318_/X _10319_/Y vssd1 vssd1 vccd1 vccd1 dest_val[7]
+ sky130_fd_sc_hd__a22o_4
XANTENNA__12000__A1 _09242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10251_ _10097_/A _10383_/A _10251_/C vssd1 vssd1 vccd1 vccd1 _10383_/B sky130_fd_sc_hd__nand3b_1
XANTENNA__08204__B1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10182_ _10155_/Y _10156_/X _10181_/X vssd1 vssd1 vccd1 vccd1 _10182_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09952__B1 _10240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout250 _06782_/X vssd1 vssd1 vccd1 vccd1 _12444_/B sky130_fd_sc_hd__clkbuf_8
Xfanout272 _06675_/B vssd1 vssd1 vccd1 vccd1 _06716_/B sky130_fd_sc_hd__clkbuf_8
Xfanout283 _06585_/Y vssd1 vssd1 vccd1 vccd1 _13142_/A sky130_fd_sc_hd__clkbuf_4
Xfanout261 _07248_/A vssd1 vssd1 vccd1 vccd1 _07585_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout294 _12359_/A vssd1 vssd1 vccd1 vccd1 _12438_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__10314__A1 _12064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12487__A _12660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12823_ _12823_/A1 _13101_/B2 hold47/X _13147_/A vssd1 vssd1 vccd1 vccd1 _13272_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11391__A _12096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10078__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12754_ _12760_/C _12753_/B _12751_/A vssd1 vssd1 vccd1 vccd1 _12756_/A sky130_fd_sc_hd__o21ai_4
X_11705_ _11705_/A _11705_/B _11705_/C vssd1 vssd1 vccd1 vccd1 _11706_/B sky130_fd_sc_hd__nand3_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13016__B1 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12685_ reg1_val[9] _12685_/B vssd1 vssd1 vccd1 vccd1 _12693_/A sky130_fd_sc_hd__nand2_1
X_11636_ _11636_/A _11636_/B _11636_/C vssd1 vssd1 vccd1 vccd1 _11637_/C sky130_fd_sc_hd__and3_1
XANTENNA__09235__A2 _11995_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09796__A _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11567_ _12050_/A _11567_/B _11567_/C _11567_/D vssd1 vssd1 vccd1 vccd1 _11567_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_4_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10518_ _10517_/A _10517_/B _10517_/C vssd1 vssd1 vccd1 vccd1 _10519_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13306_ _13309_/CLK hold210/X vssd1 vssd1 vccd1 vccd1 hold208/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07797__A2 _07959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08994__A1 _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08994__B2 _07172_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13237_ _13246_/A _13237_/B vssd1 vssd1 vccd1 vccd1 _13389_/D sky130_fd_sc_hd__and2_1
X_11498_ _07032_/Y fanout43/X fanout41/X _11946_/B vssd1 vssd1 vccd1 vccd1 _11499_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08205__A _08334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10449_ curr_PC[7] _10448_/C curr_PC[8] vssd1 vssd1 vccd1 vccd1 _10450_/C sky130_fd_sc_hd__a21oi_1
X_13168_ _13168_/A _13168_/B vssd1 vssd1 vccd1 vccd1 _13169_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09943__B1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12119_ _11440_/B _11802_/B _12115_/Y _12118_/Y vssd1 vssd1 vccd1 vccd1 _12120_/B
+ sky130_fd_sc_hd__a31o_1
X_13099_ _08874_/B _12820_/B hold7/X vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06772__A3 _12680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07660_ _07660_/A _07660_/B vssd1 vssd1 vccd1 vccd1 _07673_/A sky130_fd_sc_hd__xor2_4
X_06611_ instruction[25] _06675_/B vssd1 vssd1 vccd1 vccd1 _12642_/B sky130_fd_sc_hd__and2_4
XANTENNA__12058__A1 _10049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07591_ _07591_/A _07591_/B vssd1 vssd1 vccd1 vccd1 _07592_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_87_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09330_ _09330_/A _09330_/B _09330_/C vssd1 vssd1 vccd1 vccd1 _09331_/B sky130_fd_sc_hd__and3_1
XFILLER_0_62_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09261_ _10321_/A _10321_/B vssd1 vssd1 vccd1 vccd1 _09765_/A sky130_fd_sc_hd__or2_2
XFILLER_0_48_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08212_ _08235_/A _08235_/B _08201_/X vssd1 vssd1 vccd1 vccd1 _08224_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_62_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09192_ reg1_val[3] reg1_val[28] _09211_/S vssd1 vssd1 vccd1 vccd1 _09192_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12844__B _12862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout121_A _08334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08143_ _08125_/X _08216_/A _08153_/B vssd1 vssd1 vccd1 vccd1 _08143_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__13021__A _13162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10241__B1 _08454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08074_ _08179_/A _08179_/B _08017_/X vssd1 vssd1 vccd1 vccd1 _08076_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_113_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10792__A1 _12054_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07025_ reg1_val[2] _07025_/B vssd1 vssd1 vccd1 vccd1 _07029_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10349__B1_N _10479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10544__A1 _10276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11476__A _11476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11741__B1 _12376_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10544__B2 _10415_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ _06993_/Y fanout13/X fanout8/X _06993_/A vssd1 vssd1 vccd1 vccd1 _08977_/B
+ sky130_fd_sc_hd__o22a_2
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ _07971_/B _07927_/B vssd1 vssd1 vccd1 vccd1 _07972_/A sky130_fd_sc_hd__and2b_1
X_07858_ _09770_/B2 _08289_/B fanout75/X _09940_/B2 vssd1 vssd1 vccd1 vccd1 _07859_/B
+ sky130_fd_sc_hd__o22a_1
X_06809_ _06809_/A _06809_/B vssd1 vssd1 vccd1 vccd1 _06809_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__07712__A2 _08411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07789_ _07790_/A _07790_/B vssd1 vssd1 vccd1 vccd1 _07789_/Y sky130_fd_sc_hd__nor2_1
X_09528_ _09529_/A _09529_/B vssd1 vssd1 vccd1 vccd1 _09530_/A sky130_fd_sc_hd__and2_1
XFILLER_0_109_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout34_A _07201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09459_ _09624_/B _09459_/B vssd1 vssd1 vccd1 vccd1 _09461_/A sky130_fd_sc_hd__or2_2
XFILLER_0_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07476__B2 _07283_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07476__A1 _07221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10480__B1 _10479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12470_ _12476_/B _12470_/B vssd1 vssd1 vccd1 vccd1 new_PC[1] sky130_fd_sc_hd__and2_4
XFILLER_0_34_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11421_ _11422_/A _11422_/B vssd1 vssd1 vccd1 vccd1 _11520_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__12221__A1 _12335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12221__B2 _12286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11352_ reg1_val[16] curr_PC[16] vssd1 vssd1 vccd1 vccd1 _11353_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_62_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08976__B2 _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08976__A1 _06993_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10783__A1 _10283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10303_ hold260/A _10303_/B vssd1 vssd1 vccd1 vccd1 _10569_/C sky130_fd_sc_hd__or2_1
XFILLER_0_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11283_ fanout26/X fanout14/X fanout12/X fanout28/X vssd1 vssd1 vccd1 vccd1 _11284_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13022_ hold201/X _13171_/B2 _13209_/A2 hold162/X vssd1 vssd1 vccd1 vccd1 hold207/A
+ sky130_fd_sc_hd__a22o_1
X_10234_ fanout41/X _10234_/A2 _07274_/Y fanout43/X vssd1 vssd1 vccd1 vccd1 _10235_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10165_ _10162_/X _10164_/X _10165_/S vssd1 vssd1 vccd1 vccd1 _10165_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_100_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12288__A1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10096_ _10096_/A _10096_/B vssd1 vssd1 vccd1 vccd1 _10097_/B sky130_fd_sc_hd__or2_1
XANTENNA__07164__B1 _07147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12806_ hold9/X _12870_/B vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__or2_1
XFILLER_0_16_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12010__A _12084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10998_ _10998_/A _10998_/B vssd1 vssd1 vccd1 vccd1 _11000_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_123_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12737_ _12737_/A _12739_/D vssd1 vssd1 vccd1 vccd1 loadstore_address[19] sky130_fd_sc_hd__xnor2_4
XFILLER_0_127_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12668_ _12667_/A _12664_/Y _12666_/B vssd1 vssd1 vccd1 vccd1 _12672_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_25_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11619_ _11623_/B _11800_/A vssd1 vssd1 vccd1 vccd1 _11968_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11015__A2 _11050_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12664__B _12665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12599_ _12621_/A _12623_/A vssd1 vssd1 vccd1 vccd1 _12601_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_106_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmax_cap225 _06793_/Y vssd1 vssd1 vccd1 vccd1 _11029_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_122_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09916__B1 _11093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07774__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _07620_/A _07620_/B _07623_/Y vssd1 vssd1 vccd1 vccd1 _08834_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__06745__A3 _12708_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12279__B2 _12631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ _08761_/A _08761_/B vssd1 vssd1 vccd1 vccd1 _11444_/C sky130_fd_sc_hd__xnor2_2
X_07712_ _10338_/B2 _08411_/B _10476_/A _08457_/A2 vssd1 vssd1 vccd1 vccd1 _07713_/B
+ sky130_fd_sc_hd__o22a_1
X_08692_ _08761_/A _08766_/A _08761_/B _08363_/X vssd1 vssd1 vccd1 vccd1 _08769_/B
+ sky130_fd_sc_hd__o31ai_2
X_07643_ _07644_/A _07644_/B vssd1 vssd1 vccd1 vccd1 _07645_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_88_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout169_A _12805_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09313_ _11381_/A _09313_/B vssd1 vssd1 vccd1 vccd1 _09315_/B sky130_fd_sc_hd__xnor2_1
X_07574_ _07343_/A _07343_/B _07341_/Y vssd1 vssd1 vccd1 vccd1 _07592_/A sky130_fd_sc_hd__o21a_2
XANTENNA__07014__A _07014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08655__B1 _07173_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10462__B1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09244_ _09196_/X _09250_/B _09419_/B vssd1 vssd1 vccd1 vccd1 _09244_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09175_ _09171_/X _09174_/X _09727_/S vssd1 vssd1 vccd1 vccd1 _09175_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08126_ _06992_/A fanout84/X fanout80/X _08613_/A vssd1 vssd1 vccd1 vccd1 _08127_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09080__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06704__A2_N _06766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08057_ _08088_/A _08088_/B vssd1 vssd1 vccd1 vccd1 _08057_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_31_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07008_ reg1_val[4] _07008_/B vssd1 vssd1 vccd1 vccd1 _07010_/B sky130_fd_sc_hd__xor2_2
XANTENNA__07684__A _08454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08959_ _09066_/B _08959_/B vssd1 vssd1 vccd1 vccd1 _08984_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_98_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11970_ _11803_/Y _12114_/A _11969_/Y vssd1 vssd1 vccd1 vccd1 _11970_/X sky130_fd_sc_hd__a21o_1
X_10921_ hold185/A _10921_/B vssd1 vssd1 vccd1 vccd1 _11032_/B sky130_fd_sc_hd__or2_1
XFILLER_0_98_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06747__B _07195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10852_ _11770_/A _10852_/B vssd1 vssd1 vccd1 vccd1 _10854_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10783_ _10283_/B _10780_/X _10782_/X vssd1 vssd1 vccd1 vccd1 _10784_/B sky130_fd_sc_hd__a21o_2
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07449__A1 _10871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07449__B2 fanout86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12522_ _12685_/B _12522_/B vssd1 vssd1 vccd1 vccd1 _12523_/B sky130_fd_sc_hd__or2_1
XFILLER_0_94_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07859__A _08334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12453_ reg1_val[31] _07147_/B _11995_/B _12452_/X _12422_/A vssd1 vssd1 vccd1 vccd1
+ _12453_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08949__A1 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11404_ fanout62/X fanout23/X fanout15/X _11671_/A vssd1 vssd1 vccd1 vccd1 _11405_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_111_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12384_ _08876_/A fanout7/X _12335_/B vssd1 vssd1 vccd1 vccd1 _12384_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__08949__B2 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11335_ _11118_/A _11223_/Y _11225_/B vssd1 vssd1 vccd1 vccd1 _11335_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07621__B2 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07621__A1 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11266_ _12356_/B1 _11233_/X _11234_/Y _11236_/Y _11265_/X vssd1 vssd1 vccd1 vccd1
+ _11266_/X sky130_fd_sc_hd__a311o_1
X_13005_ _13019_/A hold183/X vssd1 vssd1 vccd1 vccd1 hold184/A sky130_fd_sc_hd__and2_1
X_10217_ _10218_/A _10218_/B vssd1 vssd1 vccd1 vccd1 _10401_/A sky130_fd_sc_hd__nor2_1
X_11197_ _11070_/A _11070_/B _11067_/A vssd1 vssd1 vccd1 vccd1 _11199_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__11181__B2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11181__A1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10148_ _10049_/Y _10147_/A _09150_/X vssd1 vssd1 vccd1 vccd1 _10148_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11844__A _11844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10079_ _12157_/A _10079_/B vssd1 vssd1 vccd1 vccd1 _10086_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__12659__B _12660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08885__B1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12984__A2 _13000_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08101__A2 _08484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07290_ _07373_/A _07373_/B vssd1 vssd1 vccd1 vccd1 _07374_/A sky130_fd_sc_hd__and2_1
XANTENNA__07769__A _09834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10195__A _11582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09601__A2 _12422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11944__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold303 hold303/A vssd1 vssd1 vccd1 vccd1 hold303/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09931_ _09931_/A _09931_/B _09816_/X vssd1 vssd1 vccd1 vccd1 _09932_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_111_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13161__A2 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09862_ _09862_/A _09862_/B vssd1 vssd1 vccd1 vccd1 _10331_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__08112__B _08112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ fanout59/X fanout86/X fanout82/X fanout57/X vssd1 vssd1 vccd1 vccd1 _09794_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07009__A _07604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08813_ _07669_/A _07669_/B _07670_/Y vssd1 vssd1 vccd1 vccd1 _08914_/A sky130_fd_sc_hd__o21ai_4
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08744_ _08744_/A _08744_/B vssd1 vssd1 vccd1 vccd1 _08744_/X sky130_fd_sc_hd__or2_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12121__B1 _11892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11473__B _12158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11475__A2 _12335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ _08624_/A _08725_/B _08624_/B vssd1 vssd1 vccd1 vccd1 _08727_/A sky130_fd_sc_hd__o21ba_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10683__B1 _12064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07626_ _07626_/A _07626_/B vssd1 vssd1 vccd1 vccd1 _07628_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08340__A2 _10338_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07557_ _07558_/A _07557_/B _07557_/C _07557_/D vssd1 vssd1 vccd1 vccd1 _07741_/A
+ sky130_fd_sc_hd__nor4_1
XANTENNA__13180__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07300__B1 _10240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07488_ _07148_/Y _07554_/B _07175_/A _07959_/A vssd1 vssd1 vccd1 vccd1 _07489_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09227_ _09239_/A _09228_/B vssd1 vssd1 vccd1 vccd1 _11829_/B sky130_fd_sc_hd__nor2_4
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07851__B2 _08540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07851__A1 _08515_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09158_ reg1_val[3] reg1_val[28] _09180_/S vssd1 vssd1 vccd1 vccd1 _09158_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11929__A _11929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08109_ _08156_/A _08156_/B vssd1 vssd1 vccd1 vccd1 _08157_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07603__B2 _09298_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07603__A1 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09089_ _09089_/A _09089_/B vssd1 vssd1 vccd1 vccd1 _09090_/B sky130_fd_sc_hd__nand2_1
X_11120_ _11120_/A _11227_/A vssd1 vssd1 vccd1 vccd1 _11334_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08303__A _08454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11051_ _11271_/A _11271_/C vssd1 vssd1 vccd1 vccd1 _11052_/B sky130_fd_sc_hd__nor2_1
X_10002_ _10137_/B _10331_/A vssd1 vssd1 vccd1 vccd1 _10278_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11664__A _11929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09659__A2 fanout86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11953_ _12036_/A _11953_/B vssd1 vssd1 vccd1 vccd1 _11955_/B sky130_fd_sc_hd__and2_1
X_11884_ _11884_/A _11965_/A vssd1 vssd1 vccd1 vccd1 _12043_/A sky130_fd_sc_hd__nor2_2
X_10904_ _11120_/A _10904_/B vssd1 vssd1 vccd1 vccd1 _11050_/C sky130_fd_sc_hd__xnor2_4
XFILLER_0_86_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10835_ _10835_/A vssd1 vssd1 vccd1 vccd1 _10836_/B sky130_fd_sc_hd__inv_2
XFILLER_0_94_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10766_ _10766_/A _10766_/B vssd1 vssd1 vccd1 vccd1 _10768_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12505_ _12511_/B _12505_/B vssd1 vssd1 vccd1 vccd1 new_PC[6] sky130_fd_sc_hd__and2_4
X_10697_ _10672_/Y _10673_/X _10684_/X _10696_/X vssd1 vssd1 vccd1 vccd1 _10697_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10729__A1 _12233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12436_ _12427_/X _12435_/Y _09149_/Y vssd1 vssd1 vccd1 vccd1 _12436_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11926__B1 _07608_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10729__B2 _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09595__A1 _11813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06940__B _06944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12367_ reg1_val[28] _12366_/C reg1_val[29] vssd1 vssd1 vccd1 vccd1 _12367_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11318_ _11318_/A _11318_/B _11318_/C vssd1 vssd1 vccd1 vccd1 _11319_/B sky130_fd_sc_hd__and3_1
X_12298_ _12298_/A _12298_/B vssd1 vssd1 vccd1 vccd1 _12430_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_38_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11249_ _11820_/A _11249_/B vssd1 vssd1 vccd1 vccd1 _11249_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06790_ _06790_/A _06790_/B vssd1 vssd1 vccd1 vccd1 _06898_/B sky130_fd_sc_hd__or2_1
XANTENNA__11457__A2 _12420_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_7_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10665__B1 _11050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08460_ _08460_/A _08460_/B vssd1 vssd1 vccd1 vccd1 _08497_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11209__A2 _12087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07411_ _09779_/A _07411_/B vssd1 vssd1 vccd1 vccd1 _07433_/B sky130_fd_sc_hd__xnor2_2
X_08391_ _08420_/A _08420_/B vssd1 vssd1 vccd1 vccd1 _08421_/A sky130_fd_sc_hd__or2_1
XFILLER_0_73_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10417__B1 _12356_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07342_ _07388_/A _07342_/B vssd1 vssd1 vccd1 vccd1 _07343_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_18_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07273_ _11038_/A _07274_/B vssd1 vssd1 vccd1 vccd1 _07273_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_73_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09012_ _09012_/A _09012_/B vssd1 vssd1 vccd1 vccd1 _09014_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12852__B _12862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold100 hold100/A vssd1 vssd1 vccd1 vccd1 hold100/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08389__A2 _08561_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold122 hold122/A vssd1 vssd1 vccd1 vccd1 hold122/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 hold133/A vssd1 vssd1 vccd1 vccd1 hold133/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 hold144/A vssd1 vssd1 vccd1 vccd1 hold144/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 hold111/A vssd1 vssd1 vccd1 vccd1 hold111/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout201_A _10243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07597__B1 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold177 hold177/A vssd1 vssd1 vccd1 vccd1 hold177/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 hold166/A vssd1 vssd1 vccd1 vccd1 hold166/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 hold155/A vssd1 vssd1 vccd1 vccd1 hold155/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 hold188/A vssd1 vssd1 vccd1 vccd1 hold188/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold199 hold199/A vssd1 vssd1 vccd1 vccd1 hold199/X sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ _07417_/B _10725_/A _07232_/X fanout42/X vssd1 vssd1 vccd1 vccd1 _09915_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09338__A1 _07830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09338__B2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09845_ _09845_/A _09845_/B vssd1 vssd1 vccd1 vccd1 _09846_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_0_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11484__A _11484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13175__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08561__A2 _08561_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06988_ _06998_/A _06995_/A vssd1 vssd1 vccd1 vccd1 _07046_/C sky130_fd_sc_hd__and2_1
X_09776_ _09776_/A _09776_/B vssd1 vssd1 vccd1 vccd1 _09780_/A sky130_fd_sc_hd__or2_1
X_08727_ _08727_/A _08727_/B vssd1 vssd1 vccd1 vccd1 _10420_/C sky130_fd_sc_hd__xnor2_2
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _08658_/A _08667_/S vssd1 vssd1 vccd1 vccd1 _08659_/B sky130_fd_sc_hd__xnor2_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_8_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13365_/CLK sky130_fd_sc_hd__clkbuf_8
X_07609_ _07983_/A _07316_/Y _07608_/Y _12642_/A vssd1 vssd1 vccd1 vccd1 _07610_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07521__B1 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08589_ _08568_/A _08568_/B _08568_/C vssd1 vssd1 vccd1 vccd1 _08589_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10959__A1 _12233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10620_ _10620_/A _10620_/B vssd1 vssd1 vccd1 vccd1 _10638_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10959__B2 _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10551_ _11630_/A _10552_/B _10552_/C vssd1 vssd1 vccd1 vccd1 _10551_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10482_ _10482_/A _10482_/B vssd1 vssd1 vccd1 vccd1 _10485_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13270_ _13365_/CLK _13270_/D vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12221_ _12335_/A _08877_/B fanout6/X _12286_/A vssd1 vssd1 vccd1 vccd1 _12222_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_121_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06760__B _06810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12152_ curr_PC[24] curr_PC[25] _12079_/B _12631_/S vssd1 vssd1 vccd1 vccd1 _12152_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08033__A _08334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07052__A2 _08613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11103_ _10956_/A _10956_/B _10976_/A vssd1 vssd1 vccd1 vccd1 _11106_/A sky130_fd_sc_hd__a21o_1
X_12083_ _12087_/B _12083_/B vssd1 vssd1 vccd1 vccd1 _12085_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12333__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11034_ _13310_/Q _11646_/B _11147_/B _11648_/A vssd1 vssd1 vccd1 vccd1 _11034_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__07760__B1 _09479_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12985_ _13001_/A hold197/X vssd1 vssd1 vccd1 vccd1 _13302_/D sky130_fd_sc_hd__and2_1
X_11936_ _11935_/B _11936_/B vssd1 vssd1 vccd1 vccd1 _11937_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08304__A2 _10221_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11867_ _11867_/A _11867_/B vssd1 vssd1 vccd1 vccd1 _11870_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11798_ _11798_/A _11798_/B vssd1 vssd1 vccd1 vccd1 _11965_/A sky130_fd_sc_hd__or2_4
XANTENNA__09804__A2 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13114__A _13147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10818_ _10818_/A _10818_/B _10818_/C _10817_/X vssd1 vssd1 vccd1 vccd1 _10818_/X
+ sky130_fd_sc_hd__or4b_1
XANTENNA__13061__A1 _10748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09265__B1 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10749_ _10749_/A _10749_/B vssd1 vssd1 vccd1 vccd1 _10751_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11569__A _12336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12419_ hold232/A _12447_/B1 _12417_/X _11648_/A vssd1 vssd1 vccd1 vccd1 _12419_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13399_ instruction[11] vssd1 vssd1 vccd1 vccd1 loadstore_dest[0] sky130_fd_sc_hd__buf_12
XANTENNA__11288__B _11288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07258__S _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07043__A2 _08657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07960_ _09836_/A _07960_/B vssd1 vssd1 vccd1 vccd1 _07962_/B sky130_fd_sc_hd__xnor2_2
X_06911_ instruction[2] _06911_/B _06911_/C vssd1 vssd1 vccd1 vccd1 _06911_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_65_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07891_ _09934_/A _08199_/B fanout33/X _09822_/A vssd1 vssd1 vccd1 vccd1 _07892_/B
+ sky130_fd_sc_hd__o22a_1
X_06842_ _06897_/D _06840_/X _06841_/X vssd1 vssd1 vccd1 vccd1 _06842_/X sky130_fd_sc_hd__a21o_1
X_09630_ _09630_/A _09630_/B vssd1 vssd1 vccd1 vccd1 _09633_/A sky130_fd_sc_hd__xor2_2
X_09561_ _10165_/S _09560_/A _09251_/A vssd1 vssd1 vccd1 vccd1 _09562_/A sky130_fd_sc_hd__o21ai_2
X_06773_ reg1_val[7] _07222_/A vssd1 vssd1 vccd1 vccd1 _06773_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_78_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11835__C1 _11834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08512_ _08518_/A _08518_/B vssd1 vssd1 vccd1 vccd1 _08512_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09492_ _11381_/A _09492_/B vssd1 vssd1 vccd1 vccd1 _09494_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout249_A _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06845__B _11134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08443_ _09670_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08447_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08374_ _08575_/A _08374_/B vssd1 vssd1 vccd1 vccd1 _08424_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__11063__B1 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07022__A _09947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07325_ _07325_/A _07325_/B vssd1 vssd1 vccd1 vccd1 _07343_/A sky130_fd_sc_hd__xnor2_2
X_07256_ _07094_/A _07093_/X _07094_/Y _06979_/Y vssd1 vssd1 vccd1 vccd1 _07256_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_0_61_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09559__A1 _11138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07187_ _11242_/A _07187_/B vssd1 vssd1 vccd1 vccd1 _07187_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11198__B _12087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07585__A3 _12779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09828_ _09828_/A _09828_/B vssd1 vssd1 vccd1 vccd1 _09830_/B sky130_fd_sc_hd__xnor2_2
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout64_A _07014_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09759_ _12365_/A _09716_/Y _09717_/X _09758_/X vssd1 vssd1 vccd1 vccd1 _09759_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_69_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08298__A1 _08657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12770_ _12770_/A _12770_/B vssd1 vssd1 vccd1 vccd1 _12780_/B sky130_fd_sc_hd__or2_1
XANTENNA__08298__B2 _08649_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06755__B _06766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11721_ _11720_/A _11720_/B _12356_/B1 vssd1 vssd1 vccd1 vccd1 _11721_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11652_ _09228_/X _09422_/B _11652_/S vssd1 vssd1 vccd1 vccd1 _11652_/X sky130_fd_sc_hd__mux2_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout50 _11484_/A vssd1 vssd1 vccd1 vccd1 _11770_/A sky130_fd_sc_hd__buf_12
X_10603_ _12009_/A fanout28/X fanout26/X fanout58/X vssd1 vssd1 vccd1 vccd1 _10604_/B
+ sky130_fd_sc_hd__o22a_1
Xfanout83 _07258_/X vssd1 vssd1 vccd1 vccd1 _10476_/A sky130_fd_sc_hd__buf_8
Xfanout61 _07019_/X vssd1 vssd1 vccd1 vccd1 fanout61/X sky130_fd_sc_hd__buf_6
Xfanout72 _10974_/A vssd1 vssd1 vccd1 vccd1 fanout72/X sky130_fd_sc_hd__buf_8
X_11583_ fanout30/X _08859_/Y _08974_/Y fanout32/X vssd1 vssd1 vccd1 vccd1 _11584_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13322_ _13392_/CLK hold164/X vssd1 vssd1 vccd1 vccd1 _13322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout94 _07146_/Y vssd1 vssd1 vccd1 vccd1 _09779_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_52_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10534_ _10534_/A _10534_/B vssd1 vssd1 vccd1 vccd1 _10536_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_51_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10465_ _10464_/B _10465_/B vssd1 vssd1 vccd1 vccd1 _10466_/B sky130_fd_sc_hd__nand2b_1
X_13253_ hold167/X hold140/X _13039_/A _13252_/X vssd1 vssd1 vccd1 vccd1 hold168/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_51_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13184_ _13184_/A _13184_/B vssd1 vssd1 vccd1 vccd1 _13184_/Y sky130_fd_sc_hd__xnor2_1
X_12204_ _12447_/B1 _12266_/B hold229/A vssd1 vssd1 vccd1 vccd1 _12206_/A sky130_fd_sc_hd__a21oi_1
X_10396_ _10394_/X _10396_/B vssd1 vssd1 vccd1 vccd1 _10397_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_60_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12135_ _10159_/B _12134_/Y _12444_/B vssd1 vssd1 vccd1 vccd1 _12135_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09970__A1 _07097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09970__B2 _07256_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12857__A1 _07032_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12066_ _12322_/A1 _12140_/B hold206/A vssd1 vssd1 vccd1 vccd1 _12066_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__13109__A _13147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ _11809_/A _08744_/X _08745_/X vssd1 vssd1 vccd1 vccd1 _11017_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07107__A _11134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12968_ hold28/X hold287/A vssd1 vssd1 vccd1 vccd1 _13238_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09486__B1 _10245_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06665__B _06675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11293__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11919_ _12446_/C1 _11906_/X _11918_/Y _11900_/Y vssd1 vssd1 vccd1 vccd1 _11919_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_75_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12899_ hold281/X hold30/X vssd1 vssd1 vccd1 vccd1 _13138_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_59_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07110_ _11134_/A _11242_/A _07141_/C _12740_/B _07248_/A vssd1 vssd1 vccd1 vccd1
+ _07210_/B sky130_fd_sc_hd__o41a_4
XFILLER_0_43_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08090_ _08664_/A _08090_/B vssd1 vssd1 vccd1 vccd1 _08122_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07041_ _07041_/A _07041_/B vssd1 vssd1 vccd1 vccd1 _07404_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_113_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08992_ _11497_/A _08992_/B vssd1 vssd1 vccd1 vccd1 _08998_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07943_ _07941_/A _07941_/B _07942_/X vssd1 vssd1 vccd1 vccd1 _08011_/A sky130_fd_sc_hd__a21o_2
XANTENNA__10859__B1 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13019__A _13019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11238__S _11813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07874_ _07874_/A _07874_/B vssd1 vssd1 vccd1 vccd1 _07946_/C sky130_fd_sc_hd__xor2_1
X_06825_ reg1_val[4] _11029_/S vssd1 vssd1 vccd1 vccd1 _06825_/X sky130_fd_sc_hd__and2_1
X_09613_ _09922_/A _09613_/B vssd1 vssd1 vccd1 vccd1 _09614_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06756_ _06927_/A _06723_/A _12696_/B _06755_/X vssd1 vssd1 vccd1 vccd1 _07233_/A
+ sky130_fd_sc_hd__a31o_4
X_09544_ _09544_/A _09544_/B vssd1 vssd1 vccd1 vccd1 _09545_/B sky130_fd_sc_hd__xor2_4
X_06687_ instruction[30] _06716_/B vssd1 vssd1 vccd1 vccd1 _12665_/B sky130_fd_sc_hd__and2_4
XFILLER_0_116_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09475_ _09476_/A _09476_/B _09476_/C vssd1 vssd1 vccd1 vccd1 _09475_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_38_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08426_ _08425_/A _08468_/A _08425_/B _08422_/X vssd1 vssd1 vccd1 vccd1 _08438_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_65_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08357_ _08357_/A _08357_/B vssd1 vssd1 vccd1 vccd1 _08402_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08288_ _10207_/A _08288_/B vssd1 vssd1 vccd1 vccd1 _08350_/A sky130_fd_sc_hd__xnor2_4
X_07308_ _07306_/A _07306_/B _07414_/A vssd1 vssd1 vccd1 vccd1 _07310_/B sky130_fd_sc_hd__o21bai_1
XFILLER_0_104_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07239_ _08112_/B _08457_/A2 fanout25/X _08501_/B1 vssd1 vssd1 vccd1 vccd1 _07240_/B
+ sky130_fd_sc_hd__o22a_2
X_10250_ _10249_/B _10249_/C _10249_/A vssd1 vssd1 vccd1 vccd1 _10251_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_14_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08204__A1 _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09952__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10547__C1 _10546_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08204__B2 _08649_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10181_ _09887_/X _10165_/X _10180_/X _10159_/Y vssd1 vssd1 vccd1 vccd1 _10181_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__09952__B2 _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07963__B1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12839__A1 _07262_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout273 _06588_/X vssd1 vssd1 vccd1 vccd1 _06675_/B sky130_fd_sc_hd__buf_4
Xfanout251 _06723_/A vssd1 vssd1 vccd1 vccd1 _06817_/B1 sky130_fd_sc_hd__buf_8
Xfanout262 _06964_/X vssd1 vssd1 vccd1 vccd1 _07248_/A sky130_fd_sc_hd__buf_4
XANTENNA__08507__A2 _12823_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout295 instruction[7] vssd1 vssd1 vccd1 vccd1 _12359_/A sky130_fd_sc_hd__buf_8
Xfanout284 _12054_/S vssd1 vssd1 vccd1 vccd1 _11813_/S sky130_fd_sc_hd__buf_6
XANTENNA__10314__A2 _12446_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12067__A2 _12322_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12822_ hold46/X _12826_/B vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__or2_1
XANTENNA__10078__B2 _10500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10078__A1 _10599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12753_ _12760_/C _12753_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[22] sky130_fd_sc_hd__xor2_4
X_11704_ _11705_/A _11705_/B _11705_/C vssd1 vssd1 vccd1 vccd1 _11797_/B sky130_fd_sc_hd__a21o_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12684_ reg1_val[9] _12685_/B vssd1 vssd1 vccd1 vccd1 _12691_/B sky130_fd_sc_hd__or2_1
X_11635_ _11636_/B _11636_/C _11636_/A vssd1 vssd1 vccd1 vccd1 _11637_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11566_ _11752_/S _11563_/X _11749_/C _11565_/Y vssd1 vssd1 vccd1 vccd1 dest_val[18]
+ sky130_fd_sc_hd__o22ai_4
XFILLER_0_24_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10517_ _10517_/A _10517_/B _10517_/C vssd1 vssd1 vccd1 vccd1 _10519_/B sky130_fd_sc_hd__or3_1
X_13305_ _13309_/CLK _13305_/D vssd1 vssd1 vccd1 vccd1 hold217/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08994__A2 _07362_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11497_ _11497_/A _11497_/B vssd1 vssd1 vccd1 vccd1 _11501_/B sky130_fd_sc_hd__xnor2_1
X_13236_ hold287/X _13248_/B1 _13235_/X _13248_/A2 vssd1 vssd1 vccd1 vccd1 _13237_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10448_ curr_PC[7] curr_PC[8] _10448_/C vssd1 vssd1 vccd1 vccd1 _10699_/C sky130_fd_sc_hd__and3_1
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13167_ _13249_/A hold271/X vssd1 vssd1 vccd1 vccd1 _13374_/D sky130_fd_sc_hd__and2_1
X_10379_ _10379_/A _10379_/B vssd1 vssd1 vccd1 vccd1 _10381_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09943__B2 _09943_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09943__A1 _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12118_ _11804_/Y _12115_/A _12117_/Y vssd1 vssd1 vccd1 vccd1 _12118_/Y sky130_fd_sc_hd__o21ai_1
X_13098_ hold6/X _06577_/A _13254_/A2 _06571_/Y rst vssd1 vssd1 vccd1 vccd1 hold7/A
+ sky130_fd_sc_hd__a221o_1
X_12049_ _12049_/A _12049_/B vssd1 vssd1 vccd1 vccd1 _12050_/C sky130_fd_sc_hd__and2_1
XANTENNA__11582__A _11582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07182__A1 _11134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06610_ instruction[1] instruction[2] instruction[0] pred_val vssd1 vssd1 vccd1 vccd1
+ _06610_/X sky130_fd_sc_hd__or4bb_4
XANTENNA__06676__A _06723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07590_ _07589_/A _07589_/C _07589_/B vssd1 vssd1 vccd1 vccd1 _07591_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__07271__S _11179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09052__A _09922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09260_ curr_PC[0] curr_PC[1] vssd1 vssd1 vccd1 vccd1 _09260_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_118_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11018__B1 _10788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08211_ _08211_/A _08211_/B vssd1 vssd1 vccd1 vccd1 _08235_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_90_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09191_ _09187_/X _09190_/X _09725_/S vssd1 vssd1 vccd1 vccd1 _09191_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09631__B1 _07269_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08142_ _08140_/A _08140_/B _08218_/A vssd1 vssd1 vccd1 vccd1 _08153_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08073_ _08073_/A _08073_/B vssd1 vssd1 vccd1 vccd1 _08179_/B sky130_fd_sc_hd__xor2_2
X_07024_ _12642_/A reg1_val[1] _07248_/A vssd1 vssd1 vccd1 vccd1 _07025_/B sky130_fd_sc_hd__o21a_1
XANTENNA_fanout114_A _07221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12860__B _12862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11757__A _12335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10544__A2 _10276_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11476__B _12335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ _12359_/A _08973_/X _06661_/X vssd1 vssd1 vccd1 vccd1 fanout8/A sky130_fd_sc_hd__a21o_2
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ _10246_/A _07926_/B vssd1 vssd1 vccd1 vccd1 _07971_/B sky130_fd_sc_hd__xnor2_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08370__B1 _09770_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07857_ _10207_/A _07857_/B vssd1 vssd1 vccd1 vccd1 _07883_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06808_ reg1_val[2] _07172_/A vssd1 vssd1 vccd1 vccd1 _06809_/B sky130_fd_sc_hd__or2_1
X_07788_ _11381_/A _07788_/B vssd1 vssd1 vccd1 vccd1 _07790_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11257__B1 _12376_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06739_ reg2_val[13] _06810_/B vssd1 vssd1 vccd1 vccd1 _06739_/X sky130_fd_sc_hd__and2_1
X_09527_ _09527_/A _09527_/B vssd1 vssd1 vccd1 vccd1 _09529_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09870__B1 _12356_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09458_ _09457_/B _09458_/B vssd1 vssd1 vccd1 vccd1 _09459_/B sky130_fd_sc_hd__and2b_1
XANTENNA_fanout27_A fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07476__A2 _08112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12527__S _12638_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09389_ _09177_/X _09179_/X _09403_/S vssd1 vssd1 vccd1 vccd1 _09389_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08409_ _09472_/A _08484_/B _09479_/B1 _08649_/B1 vssd1 vssd1 vccd1 vccd1 _08410_/B
+ sky130_fd_sc_hd__o22a_1
X_11420_ _11320_/A _11320_/B _11319_/A vssd1 vssd1 vccd1 vccd1 _11422_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12221__A2 _08877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11351_ reg1_val[16] curr_PC[16] vssd1 vssd1 vccd1 vccd1 _11351_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08976__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11980__A1 _11813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10302_ hold215/A _11990_/A1 _10434_/B _12205_/B1 vssd1 vssd1 vccd1 vccd1 _10302_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11282_ _11282_/A _11282_/B vssd1 vssd1 vccd1 vccd1 _11291_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11841__D_N _11807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08189__B1 _09770_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13021_ _13162_/A hold202/X vssd1 vssd1 vccd1 vccd1 hold203/A sky130_fd_sc_hd__and2_1
X_10233_ _10233_/A _10233_/B vssd1 vssd1 vccd1 vccd1 _10237_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_100_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10164_ _09436_/Y _11138_/B _11138_/A vssd1 vssd1 vccd1 vccd1 _10164_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12288__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10095_ _10096_/A _10096_/B vssd1 vssd1 vccd1 vccd1 _10097_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09571__S _10297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11496__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07164__A1 _07172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06927__C _12218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12805_ _12805_/A _12805_/B vssd1 vssd1 vccd1 vccd1 _12805_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_123_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10997_ _10997_/A _10997_/B vssd1 vssd1 vccd1 vccd1 _10998_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_96_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12996__B1 _13257_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08113__B1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ reg1_val[19] _12755_/B vssd1 vssd1 vccd1 vccd1 _12739_/D sky130_fd_sc_hd__xnor2_4
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12667_ _12667_/A _12667_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[5] sky130_fd_sc_hd__xor2_4
XFILLER_0_108_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11618_ _11618_/A _11711_/A vssd1 vssd1 vccd1 vccd1 _11800_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_53_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12598_ _12598_/A _12598_/B _12598_/C vssd1 vssd1 vccd1 vccd1 _12623_/A sky130_fd_sc_hd__and3_1
XFILLER_0_108_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11549_ hold246/A hold292/A _11549_/C vssd1 vssd1 vccd1 vccd1 _11649_/B sky130_fd_sc_hd__or3_1
XFILLER_0_52_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12680__B _12680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13219_ _13249_/A _13219_/B vssd1 vssd1 vccd1 vccd1 _13385_/D sky130_fd_sc_hd__and2_1
XANTENNA__09916__A1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09916__B2 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_10_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13360_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08760_ _11345_/C _11345_/D _11345_/B vssd1 vssd1 vccd1 vccd1 _11444_/B sky130_fd_sc_hd__a21oi_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08886__A _09341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07711_ _07731_/A _07731_/B vssd1 vssd1 vccd1 vccd1 _07711_/Y sky130_fd_sc_hd__nand2_1
X_08691_ _08691_/A _08691_/B vssd1 vssd1 vccd1 vccd1 _08761_/B sky130_fd_sc_hd__or2_2
X_07642_ _07642_/A _07642_/B vssd1 vssd1 vccd1 vccd1 _07644_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09312_ fanout98/X _08199_/B fanout33/X fanout84/X vssd1 vssd1 vccd1 vccd1 _09313_/B
+ sky130_fd_sc_hd__o22a_1
X_07573_ _07503_/A _07503_/B _07504_/Y vssd1 vssd1 vccd1 vccd1 _07674_/A sky130_fd_sc_hd__a21bo_2
XANTENNA__08655__B2 _09218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10462__A1 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10462__B2 _12009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09243_ _11029_/S _09250_/B vssd1 vssd1 vccd1 vccd1 _09251_/A sky130_fd_sc_hd__or2_4
XFILLER_0_35_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09174_ _09172_/X _09173_/X _09403_/S vssd1 vssd1 vccd1 vccd1 _09174_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08125_ _08131_/A _08131_/B vssd1 vssd1 vccd1 vccd1 _08125_/X sky130_fd_sc_hd__and2_1
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09080__A1 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09080__B2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08056_ _08056_/A _08056_/B vssd1 vssd1 vccd1 vccd1 _08088_/B sky130_fd_sc_hd__xnor2_2
X_07007_ reg1_val[3] _07007_/B vssd1 vssd1 vccd1 vccd1 _08658_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_12_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08958_ _08957_/B _08958_/B vssd1 vssd1 vccd1 vccd1 _08959_/B sky130_fd_sc_hd__and2b_1
X_07909_ _07910_/B _07910_/C _08656_/A vssd1 vssd1 vccd1 vccd1 _07913_/A sky130_fd_sc_hd__o21ai_1
X_08889_ _08890_/A _08890_/B vssd1 vssd1 vccd1 vccd1 _08946_/A sky130_fd_sc_hd__and2_2
XFILLER_0_98_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10920_ _10917_/X _10919_/Y _11820_/A _10914_/X vssd1 vssd1 vccd1 vccd1 _10920_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_85_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10851_ _07032_/Y fanout32/X fanout30/X _11946_/B vssd1 vssd1 vccd1 vccd1 _10852_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12978__B1 _13257_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10782_ _10545_/Y _11009_/A _10781_/Y vssd1 vssd1 vccd1 vccd1 _10782_/X sky130_fd_sc_hd__a21o_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07449__A2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12521_ _12685_/B _12522_/B vssd1 vssd1 vccd1 vccd1 _12532_/A sky130_fd_sc_hd__nand2_1
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12452_ reg1_val[31] _07147_/B _11554_/A vssd1 vssd1 vccd1 vccd1 _12452_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_124_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11403_ _12017_/A _11403_/B vssd1 vssd1 vccd1 vccd1 _11409_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08949__A2 _10473_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11402__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12383_ _12336_/A _12336_/B _12339_/A vssd1 vssd1 vccd1 vccd1 _12389_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_50_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11334_ _11334_/A _11528_/A vssd1 vssd1 vccd1 vccd1 _11334_/X sky130_fd_sc_hd__and2_1
XANTENNA__07621__A2 _10245_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11265_ _11265_/A _11265_/B _11265_/C vssd1 vssd1 vccd1 vccd1 _11265_/X sky130_fd_sc_hd__or3_1
X_13004_ hold193/A _13171_/B2 _13209_/A2 hold182/X vssd1 vssd1 vccd1 vccd1 hold183/A
+ sky130_fd_sc_hd__a22o_1
X_10216_ _10086_/A _10086_/B _10084_/Y vssd1 vssd1 vccd1 vccd1 _10218_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_30_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11196_ _11196_/A _11196_/B vssd1 vssd1 vccd1 vccd1 _11204_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__11181__A2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10147_ _10147_/A vssd1 vssd1 vccd1 vccd1 _10147_/Y sky130_fd_sc_hd__inv_2
X_10078_ _10599_/A fanout23/X fanout15/X _10500_/A vssd1 vssd1 vccd1 vccd1 _10079_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06938__B _06944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08885__B2 _07198_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08885__A1 _10871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12675__B _12675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12719_ reg1_val[15] _12719_/B vssd1 vssd1 vccd1 vccd1 _12721_/C sky130_fd_sc_hd__xnor2_2
XANTENNA__10476__A _10476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11944__A1 _12233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11944__B2 _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold304 hold304/A vssd1 vssd1 vccd1 vccd1 hold304/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09930_ _09931_/A _09931_/B _09816_/X vssd1 vssd1 vccd1 vccd1 _09930_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_0_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09861_ _09861_/A _09861_/B vssd1 vssd1 vccd1 vccd1 _09862_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_0_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _10749_/A _09792_/B vssd1 vssd1 vccd1 vccd1 _09799_/A sky130_fd_sc_hd__xnor2_1
X_08812_ _07674_/A _07674_/B _07672_/X vssd1 vssd1 vccd1 vccd1 _08917_/A sky130_fd_sc_hd__a21oi_4
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ _08743_/A _08743_/B vssd1 vssd1 vccd1 vccd1 _08744_/B sky130_fd_sc_hd__and2_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13027__A _13162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout279_A _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout181_A _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08674_ _08674_/A _08674_/B vssd1 vssd1 vccd1 vccd1 _08723_/B sky130_fd_sc_hd__or2_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07625_ _07626_/A _07626_/B vssd1 vssd1 vccd1 vccd1 _07625_/X sky130_fd_sc_hd__and2_1
XANTENNA__11770__A _11770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13082__C1 _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07556_ _07556_/A _07556_/B _07556_/C vssd1 vssd1 vccd1 vccd1 _07557_/D sky130_fd_sc_hd__nor3_1
XANTENNA__10435__A1 _11990_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09226_ _09232_/A _09226_/B vssd1 vssd1 vccd1 vccd1 _09226_/X sky130_fd_sc_hd__or2_1
XFILLER_0_63_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07300__A1 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07300__B2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07487_ _07682_/A _07682_/B _07486_/C vssd1 vssd1 vccd1 vccd1 _07490_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07851__A2 _10595_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10199__B1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09157_ reg1_val[2] reg1_val[29] _09180_/S vssd1 vssd1 vccd1 vccd1 _09157_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07695__A _09672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08108_ _08108_/A _08108_/B vssd1 vssd1 vccd1 vccd1 _08156_/B sky130_fd_sc_hd__xnor2_1
X_09088_ _09089_/A _09089_/B vssd1 vssd1 vccd1 vccd1 _09281_/B sky130_fd_sc_hd__or2_1
XANTENNA__07603__A2 _09298_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06811__B1 _06810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08039_ _06992_/A _09661_/B2 fanout98/X _08613_/A vssd1 vssd1 vccd1 vccd1 _08040_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12360__A1 _12359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11050_ _11050_/A _11050_/B _11050_/C _11050_/D vssd1 vssd1 vccd1 vccd1 _11271_/C
+ sky130_fd_sc_hd__or4_2
XANTENNA__11163__A2 _11124_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11945__A _12336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10001_ _09862_/A _09862_/B _10000_/X vssd1 vssd1 vccd1 vccd1 _10001_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__06758__B _07233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11952_ _11952_/A _11952_/B _11952_/C vssd1 vssd1 vccd1 vccd1 _11953_/B sky130_fd_sc_hd__or3_1
X_11883_ _11883_/A _11883_/B vssd1 vssd1 vccd1 vccd1 _12042_/A sky130_fd_sc_hd__nand2_4
X_10903_ _10416_/A _10902_/X _10901_/X vssd1 vssd1 vccd1 vccd1 _10904_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_58_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10834_ _10834_/A _10834_/B vssd1 vssd1 vccd1 vccd1 _10835_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10765_ _10765_/A _10765_/B vssd1 vssd1 vccd1 vccd1 _10766_/B sky130_fd_sc_hd__xnor2_1
X_12504_ _12504_/A _12504_/B _12504_/C vssd1 vssd1 vccd1 vccd1 _12505_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_81_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10696_ _09222_/Y _10682_/X _10695_/Y _10159_/A _10694_/X vssd1 vssd1 vccd1 vccd1
+ _10696_/X sky130_fd_sc_hd__o221a_1
X_12435_ _12435_/A _12435_/B vssd1 vssd1 vccd1 vccd1 _12435_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11926__B2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11926__A1 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10729__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12366_ reg1_val[28] reg1_val[29] _12366_/C vssd1 vssd1 vccd1 vccd1 _12444_/C sky130_fd_sc_hd__and3_1
X_11317_ _11318_/A _11318_/B _11318_/C vssd1 vssd1 vccd1 vccd1 _11319_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_105_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12297_ _12297_/A vssd1 vssd1 vccd1 vccd1 _12298_/B sky130_fd_sc_hd__inv_2
XANTENNA__11139__C1 _11029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11248_ _11029_/S _11246_/X _11247_/X vssd1 vssd1 vccd1 vccd1 _11249_/B sky130_fd_sc_hd__a21oi_2
X_11179_ _11179_/A _11179_/B vssd1 vssd1 vccd1 vccd1 _11180_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09325__A _09325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08307__B1 _09940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10114__B1 _11198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11590__A _11591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07410_ _07507_/A _07507_/B vssd1 vssd1 vccd1 vccd1 _07433_/A sky130_fd_sc_hd__or2_1
XFILLER_0_9_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08390_ _08564_/A _08390_/B vssd1 vssd1 vccd1 vccd1 _08420_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07341_ _07388_/A _07342_/B vssd1 vssd1 vccd1 vccd1 _07341_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_116_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06718__A2_N _06766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07272_ _07195_/A _07215_/B _07195_/B vssd1 vssd1 vccd1 vccd1 _07274_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_73_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12625__S _12638_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09011_ _09010_/A _08880_/B _09010_/Y vssd1 vssd1 vccd1 vccd1 _09012_/B sky130_fd_sc_hd__a21oi_2
Xhold101 hold101/A vssd1 vssd1 vccd1 vccd1 hold101/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold123 hold123/A vssd1 vssd1 vccd1 vccd1 hold123/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 hold134/A vssd1 vssd1 vccd1 vccd1 hold134/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 hold112/A vssd1 vssd1 vccd1 vccd1 hold112/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07597__B2 _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07597__A1 _09325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold167 hold298/A vssd1 vssd1 vccd1 vccd1 hold167/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold145 hold145/A vssd1 vssd1 vccd1 vccd1 hold145/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 hold156/A vssd1 vssd1 vccd1 vccd1 hold156/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold189 hold189/A vssd1 vssd1 vccd1 vccd1 hold189/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 hold178/A vssd1 vssd1 vccd1 vccd1 hold178/X sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ _09821_/A _09821_/B _09820_/A vssd1 vssd1 vccd1 vccd1 _09926_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_0_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09338__A2 _07198_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09844_ _09845_/A _09845_/B vssd1 vssd1 vccd1 vccd1 _09844_/Y sky130_fd_sc_hd__nor2_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06987_ _06987_/A _06987_/B vssd1 vssd1 vccd1 vccd1 _06987_/Y sky130_fd_sc_hd__nand2_1
X_09775_ _09774_/B _09775_/B vssd1 vssd1 vccd1 vccd1 _09776_/B sky130_fd_sc_hd__and2b_1
X_08726_ _10287_/B _10287_/C vssd1 vssd1 vccd1 vccd1 _10420_/B sky130_fd_sc_hd__and2_2
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ _12808_/A _08657_/B vssd1 vssd1 vccd1 vccd1 _08667_/S sky130_fd_sc_hd__nor2_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07608_ _07608_/A _07608_/B vssd1 vssd1 vccd1 vccd1 _07608_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__07521__A1 _08540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07521__B2 _08515_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08588_ _08592_/A _08592_/B vssd1 vssd1 vccd1 vccd1 _08588_/X sky130_fd_sc_hd__and2_1
XFILLER_0_119_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10959__A2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07539_ _07529_/A _07735_/A _07559_/B vssd1 vssd1 vccd1 vccd1 _07539_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_106_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10550_ _11538_/A _10549_/B _10581_/C vssd1 vssd1 vccd1 vccd1 _10550_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_17_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10481_ _10481_/A _10481_/B vssd1 vssd1 vccd1 vccd1 _10482_/B sky130_fd_sc_hd__nand2_1
X_09209_ _09207_/X _09208_/X _09403_/S vssd1 vssd1 vccd1 vccd1 _09209_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11908__A1 _12447_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12220_ curr_PC[27] _12220_/B vssd1 vssd1 vccd1 vccd1 _12220_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_32_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12151_ curr_PC[25] _12216_/C vssd1 vssd1 vccd1 vccd1 _12151_/Y sky130_fd_sc_hd__nor2_1
X_11102_ _11102_/A _11102_/B vssd1 vssd1 vccd1 vccd1 _11107_/A sky130_fd_sc_hd__or2_1
X_12082_ _12233_/B fanout10/X fanout5/X _12233_/A vssd1 vssd1 vccd1 vccd1 _12083_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12333__B2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11033_ _11646_/B _11147_/B _13310_/Q vssd1 vssd1 vccd1 vccd1 _11033_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12333__A1 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07760__A1 _10595_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12984_ hold300/X _13000_/A2 _13257_/A2 hold196/X vssd1 vssd1 vccd1 vccd1 hold197/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07760__B2 _10338_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11935_ _11936_/B _11935_/B vssd1 vssd1 vccd1 vccd1 _12030_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11866_ _11867_/A _11867_/B vssd1 vssd1 vccd1 vccd1 _11952_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_86_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11797_ _11797_/A _11797_/B _11797_/C vssd1 vssd1 vccd1 vccd1 _11798_/B sky130_fd_sc_hd__and3_1
XFILLER_0_95_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10817_ _09222_/Y _10803_/X _10804_/X _09242_/B _10816_/X vssd1 vssd1 vccd1 vccd1
+ _10817_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_55_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13061__A2 _13101_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09265__A1 _09934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09265__B2 _09822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10748_ _10748_/A _10749_/B vssd1 vssd1 vccd1 vccd1 _10874_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_55_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12418_ _12447_/B1 _12417_/X hold232/A vssd1 vssd1 vccd1 vccd1 _12418_/Y sky130_fd_sc_hd__a21oi_1
X_10679_ _10679_/A _10679_/B _10679_/C vssd1 vssd1 vccd1 vccd1 _10679_/X sky130_fd_sc_hd__and3_1
XFILLER_0_2_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13398_ _13398_/CLK hold161/X vssd1 vssd1 vccd1 vccd1 hold160/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10583__B1 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12349_ _12430_/A _12430_/B vssd1 vssd1 vccd1 vccd1 _12350_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06910_ instruction[2] _06911_/B _06911_/C vssd1 vssd1 vccd1 vccd1 _12218_/A sky130_fd_sc_hd__and3_4
XANTENNA__08528__B1 _09770_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10335__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07890_ _07889_/B _07889_/C _07889_/A vssd1 vssd1 vccd1 vccd1 _07932_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__09055__A _09779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06841_ _07195_/A reg1_val[12] vssd1 vssd1 vccd1 vccd1 _06841_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_65_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09560_ _09560_/A vssd1 vssd1 vccd1 vccd1 _09560_/Y sky130_fd_sc_hd__inv_2
X_06772_ _06815_/A _06817_/B1 _12680_/B _06771_/X vssd1 vssd1 vccd1 vccd1 _07222_/A
+ sky130_fd_sc_hd__a31o_4
XANTENNA__06642__A2_N _06766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09491_ _09661_/B2 _08199_/B fanout33/X fanout98/X vssd1 vssd1 vccd1 vccd1 _09492_/B
+ sky130_fd_sc_hd__o22a_1
X_08511_ _08511_/A _08511_/B vssd1 vssd1 vccd1 vccd1 _08518_/B sky130_fd_sc_hd__xnor2_2
X_08442_ _09669_/B2 _09770_/B2 _09940_/B2 _08627_/A2 vssd1 vssd1 vccd1 vccd1 _08443_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07303__A _09667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08373_ _08657_/B _08457_/A2 _08501_/B1 _08649_/A2 vssd1 vssd1 vccd1 vccd1 _08374_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_128_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11063__B2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11063__A1 _12233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07324_ _07325_/A _07325_/B vssd1 vssd1 vccd1 vccd1 _07601_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07255_ _07255_/A _07255_/B vssd1 vssd1 vccd1 vccd1 _07255_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_73_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06861__B _07014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10664__A _10900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07186_ _11134_/A _07141_/C _07585_/B1 vssd1 vssd1 vccd1 vccd1 _07187_/B sky130_fd_sc_hd__o21a_1
XANTENNA__11495__A _12336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09827_ _09827_/A _09827_/B vssd1 vssd1 vccd1 vccd1 _09828_/B sky130_fd_sc_hd__xor2_2
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09758_ _12446_/C1 _09732_/X _09738_/X _09757_/X vssd1 vssd1 vccd1 vccd1 _09758_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_69_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08709_ _08802_/A _08802_/B _08707_/X _07818_/X _07747_/Y vssd1 vssd1 vccd1 vccd1
+ _08710_/B sky130_fd_sc_hd__a32o_2
XANTENNA_fanout57_A _07035_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11720_ _11720_/A _11720_/B vssd1 vssd1 vccd1 vccd1 _11720_/Y sky130_fd_sc_hd__nand2_1
X_09689_ _09687_/Y _09689_/B vssd1 vssd1 vccd1 vccd1 _09690_/B sky130_fd_sc_hd__and2b_1
XANTENNA__08298__A2 _10595_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11651_ _11650_/B _11739_/B hold262/A vssd1 vssd1 vccd1 vccd1 _11651_/X sky130_fd_sc_hd__a21o_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout40 _07170_/Y vssd1 vssd1 vccd1 vccd1 _07171_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__13043__A2 _12820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11582_ _11582_/A _11582_/B vssd1 vssd1 vccd1 vccd1 _11586_/A sky130_fd_sc_hd__xnor2_1
X_10602_ _11393_/A _10602_/B vssd1 vssd1 vccd1 vccd1 _10606_/A sky130_fd_sc_hd__xnor2_1
Xfanout73 _07273_/X vssd1 vssd1 vccd1 vccd1 _10974_/A sky130_fd_sc_hd__buf_6
XANTENNA__12251__B1 _09150_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout62 _07019_/X vssd1 vssd1 vccd1 vccd1 fanout62/X sky130_fd_sc_hd__buf_4
Xfanout51 _07079_/X vssd1 vssd1 vccd1 vccd1 fanout51/X sky130_fd_sc_hd__buf_8
XFILLER_0_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13321_ _13373_/CLK _13321_/D vssd1 vssd1 vccd1 vccd1 hold206/A sky130_fd_sc_hd__dfxtp_1
X_10533_ _10534_/A _10534_/B vssd1 vssd1 vccd1 vccd1 _10655_/A sky130_fd_sc_hd__nand2_1
Xfanout95 _07116_/X vssd1 vssd1 vccd1 vccd1 _11929_/A sky130_fd_sc_hd__buf_8
XFILLER_0_52_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout84 _11309_/A vssd1 vssd1 vccd1 vccd1 fanout84/X sky130_fd_sc_hd__buf_6
XANTENNA__06771__B _06810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10464_ _10465_/B _10464_/B vssd1 vssd1 vccd1 vccd1 _10618_/B sky130_fd_sc_hd__nand2b_1
X_13252_ hold167/X _13254_/A2 _12797_/Y _06577_/A vssd1 vssd1 vccd1 vccd1 _13252_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13183_ _13183_/A _13183_/B vssd1 vssd1 vccd1 vccd1 _13184_/B sky130_fd_sc_hd__nand2_1
X_12203_ _13322_/Q _12203_/B vssd1 vssd1 vccd1 vccd1 _12266_/B sky130_fd_sc_hd__or2_1
X_10395_ _10395_/A _10395_/B _10395_/C vssd1 vssd1 vccd1 vccd1 _10396_/B sky130_fd_sc_hd__or3_1
XFILLER_0_32_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12134_ _12134_/A _12134_/B vssd1 vssd1 vccd1 vccd1 _12134_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__09970__A2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08979__A _09947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06784__A2 _06783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12857__A2 _12863_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12065_ hold201/A _12065_/B vssd1 vssd1 vccd1 vccd1 _12140_/B sky130_fd_sc_hd__or2_1
X_11016_ _10937_/X _11050_/D _11015_/Y vssd1 vssd1 vccd1 vccd1 _11016_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07107__B _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08930__B1 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12967_ _13234_/A _12966_/B _12876_/X vssd1 vssd1 vccd1 vccd1 _13239_/A sky130_fd_sc_hd__a21o_1
XANTENNA__10749__A _10749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09486__B2 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09486__A1 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11293__B2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11293__A1 _11671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11918_ _11908_/Y _11909_/X _11917_/X vssd1 vssd1 vccd1 vccd1 _11918_/Y sky130_fd_sc_hd__o21ai_1
X_12898_ hold252/X hold32/X vssd1 vssd1 vccd1 vccd1 _13143_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_59_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11849_ _11939_/A _11849_/B vssd1 vssd1 vccd1 vccd1 _11851_/A sky130_fd_sc_hd__nand2_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11045__A1 _09225_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06962__A _12404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07040_ _07604_/A _07040_/B vssd1 vssd1 vccd1 vccd1 _07404_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08991_ _09325_/A _08877_/B fanout6/X _12808_/A vssd1 vssd1 vccd1 vccd1 _08992_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_11_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07942_ _07953_/B _07953_/A vssd1 vssd1 vccd1 vccd1 _07942_/X sky130_fd_sc_hd__and2b_1
XANTENNA__10859__A1 _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10859__B2 _11198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07873_ _07880_/A _07880_/B vssd1 vssd1 vccd1 vccd1 _07946_/B sky130_fd_sc_hd__and2b_1
X_06824_ _09745_/B _06822_/X _06823_/X vssd1 vssd1 vccd1 vccd1 _06824_/X sky130_fd_sc_hd__a21o_1
X_09612_ _07554_/B _10725_/A _07232_/X _07175_/A vssd1 vssd1 vccd1 vccd1 _09613_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12858__B _12862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09543_ _09544_/A _09544_/B vssd1 vssd1 vccd1 vccd1 _09543_/X sky130_fd_sc_hd__and2_1
X_06755_ reg2_val[10] _06766_/B vssd1 vssd1 vccd1 vccd1 _06755_/X sky130_fd_sc_hd__and2_1
XANTENNA__11808__B1 _09150_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13035__A _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06686_ _11913_/S _06686_/B vssd1 vssd1 vccd1 vccd1 _06860_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_78_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09474_ _11946_/C _09474_/B vssd1 vssd1 vccd1 vccd1 _09476_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__08129__A _08575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07488__B1 _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09229__A1 _11637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08425_ _08425_/A _08425_/B vssd1 vssd1 vccd1 vccd1 _08468_/B sky130_fd_sc_hd__nor2_1
X_08356_ _08365_/B _08365_/A vssd1 vssd1 vccd1 vccd1 _08357_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_18_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08988__B1 _11844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07307_ _07413_/A _07413_/B vssd1 vssd1 vccd1 vccd1 _07414_/A sky130_fd_sc_hd__nor2_2
XANTENNA__06591__B _06944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08287_ _09472_/A _08411_/B _10476_/A _08649_/B1 vssd1 vssd1 vccd1 vccd1 _08288_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_18_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07238_ _07238_/A _07238_/B vssd1 vssd1 vccd1 vccd1 _07238_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_6_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07169_ _07168_/A _07168_/B _07168_/C vssd1 vssd1 vccd1 vccd1 _07170_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08204__A2 _08289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10180_ _06782_/X _12446_/C1 _10179_/Y _10174_/X _10169_/Y vssd1 vssd1 vccd1 vccd1
+ _10180_/X sky130_fd_sc_hd__a311o_1
XANTENNA__09952__A2 _08484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07963__A1 _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12839__A2 _12863_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout230 _06677_/B1 vssd1 vssd1 vccd1 vccd1 _06724_/B1 sky130_fd_sc_hd__buf_4
Xfanout241 _06960_/X vssd1 vssd1 vccd1 vccd1 _12422_/A sky130_fd_sc_hd__buf_4
XANTENNA__07963__B2 _08649_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout274 _13019_/A vssd1 vssd1 vccd1 vccd1 _13210_/A sky130_fd_sc_hd__buf_4
Xfanout263 _12639_/A vssd1 vssd1 vccd1 vccd1 _12633_/A sky130_fd_sc_hd__clkbuf_8
Xfanout252 _06703_/A vssd1 vssd1 vccd1 vccd1 _06723_/A sky130_fd_sc_hd__clkbuf_8
Xfanout285 _12404_/S vssd1 vssd1 vccd1 vccd1 _12054_/S sky130_fd_sc_hd__buf_4
X_12821_ _07282_/Y _13101_/B2 hold19/X _13147_/A vssd1 vssd1 vccd1 vccd1 _13271_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__06766__B _06766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10078__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12752_ _12744_/Y _12748_/B _12746_/B vssd1 vssd1 vccd1 vccd1 _12753_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_29_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11703_ _11703_/A _11703_/B vssd1 vssd1 vccd1 vccd1 _11705_/C sky130_fd_sc_hd__xnor2_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12683_ _12682_/A _12679_/Y _12681_/B vssd1 vssd1 vccd1 vccd1 _12687_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_127_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13016__A2 _13171_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11634_ _12359_/A _11634_/B vssd1 vssd1 vccd1 vccd1 _11636_/C sky130_fd_sc_hd__or2_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11565_ curr_PC[18] _11564_/B _11752_/S vssd1 vssd1 vccd1 vccd1 _11565_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11496_ _11671_/A fanout10/X fanout5/X fanout52/X vssd1 vssd1 vccd1 vccd1 _11497_/B
+ sky130_fd_sc_hd__o22a_1
X_10516_ _10516_/A _10516_/B vssd1 vssd1 vccd1 vccd1 _10517_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13304_ _13304_/CLK _13304_/D vssd1 vssd1 vccd1 vccd1 hold215/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13235_ hold282/X _13234_/Y fanout2/A vssd1 vssd1 vccd1 vccd1 _13235_/X sky130_fd_sc_hd__mux2_1
X_10447_ _10788_/A _10419_/X _10420_/Y _10446_/X _10418_/X vssd1 vssd1 vccd1 vccd1
+ _10447_/X sky130_fd_sc_hd__o311a_1
XFILLER_0_40_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13166_ hold270/X _13209_/A2 _13165_/X _13171_/B2 vssd1 vssd1 vccd1 vccd1 hold271/A
+ sky130_fd_sc_hd__a22o_1
X_10378_ _10379_/B _10379_/A vssd1 vssd1 vccd1 vccd1 _10525_/B sky130_fd_sc_hd__and2b_1
XANTENNA__09943__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08502__A _08502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12117_ _11969_/Y _12114_/B _12116_/Y vssd1 vssd1 vccd1 vccd1 _12117_/Y sky130_fd_sc_hd__a21oi_1
X_13097_ _09936_/A _12820_/B _13096_/X vssd1 vssd1 vccd1 vccd1 _13358_/D sky130_fd_sc_hd__a21oi_1
X_12048_ _12300_/A _12048_/B vssd1 vssd1 vccd1 vccd1 _12184_/A sky130_fd_sc_hd__xor2_2
XANTENNA__07182__A2 _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06676__B _12680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10479__A _10479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11266__A1 _12356_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08210_ _08208_/A _08208_/B _08270_/A vssd1 vssd1 vccd1 vccd1 _08235_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__07788__A _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09190_ _09188_/X _09189_/X _09383_/S vssd1 vssd1 vccd1 vccd1 _09190_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09631__B2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09631__A1 _07959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08141_ _08217_/A _08217_/B vssd1 vssd1 vccd1 vccd1 _08218_/A sky130_fd_sc_hd__or2_1
XFILLER_0_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08072_ _08072_/A _08072_/B vssd1 vssd1 vccd1 vccd1 _08179_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_125_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07023_ _07041_/A _07041_/B vssd1 vssd1 vccd1 vccd1 _07023_/X sky130_fd_sc_hd__or2_1
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13191__B2 _13223_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11476__C _11591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08974_ _12359_/A _08973_/X _06661_/X vssd1 vssd1 vccd1 vccd1 _08974_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__buf_1
XANTENNA__07028__A _09672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07925_ _08540_/B _10595_/A1 _10338_/B2 _08515_/A2 vssd1 vssd1 vccd1 vccd1 _07926_/B
+ sky130_fd_sc_hd__o22a_1
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08370__A1 _08641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07856_ _08501_/B1 _08411_/B _10476_/A _10221_/B2 vssd1 vssd1 vccd1 vccd1 _07857_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09243__A _11029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06807_ reg1_val[2] _07172_/A vssd1 vssd1 vccd1 vccd1 _09743_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08370__B2 _08627_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07787_ _09934_/A fanout33/X _07283_/X _08199_/B vssd1 vssd1 vccd1 vccd1 _07788_/B
+ sky130_fd_sc_hd__o22a_1
X_06738_ _06738_/A _11150_/S vssd1 vssd1 vccd1 vccd1 _11131_/A sky130_fd_sc_hd__nor2_1
X_09526_ _09527_/A _09527_/B vssd1 vssd1 vccd1 vccd1 _09694_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09457_ _09458_/B _09457_/B vssd1 vssd1 vccd1 vccd1 _09624_/B sky130_fd_sc_hd__and2b_1
X_06669_ _12207_/S vssd1 vssd1 vccd1 vccd1 _06669_/Y sky130_fd_sc_hd__inv_2
X_08408_ _08408_/A _08408_/B vssd1 vssd1 vccd1 vccd1 _08427_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_108_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09388_ _09386_/X _09387_/X _09727_/S vssd1 vssd1 vccd1 vccd1 _09388_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_117_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08339_ _08342_/A _08342_/B vssd1 vssd1 vccd1 vccd1 _08339_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11350_ _11243_/B _11245_/B _11243_/A vssd1 vssd1 vccd1 vccd1 _11354_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_61_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10301_ _11990_/A1 _10434_/B hold215/A vssd1 vssd1 vccd1 vccd1 _10301_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11281_ _11282_/A _11282_/B vssd1 vssd1 vccd1 vccd1 _11417_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10852__A _11770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13020_ hold219/A _13171_/B2 _13209_/A2 hold201/X vssd1 vssd1 vccd1 vccd1 hold202/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08189__A1 _08540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08189__B2 _08515_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10232_ _10233_/A _10233_/B vssd1 vssd1 vccd1 vccd1 _10376_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_30_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10163_ _09570_/X _09573_/X _10297_/S vssd1 vssd1 vccd1 vccd1 _11138_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10940__B1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11683__A _12096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10094_ _11582_/A _10094_/B vssd1 vssd1 vccd1 vccd1 _10096_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11496__A1 _11671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11496__B2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07164__A2 _07149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09153__A _12438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12804_ _12804_/A _12804_/B vssd1 vssd1 vccd1 vccd1 _12816_/B sky130_fd_sc_hd__nor2_2
XANTENNA__11248__A1 _11029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10996_ _10997_/A _10997_/B vssd1 vssd1 vccd1 vccd1 _10996_/Y sky130_fd_sc_hd__nand2_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09310__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08113__A1 _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08113__B2 _08649_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08992__A _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _12739_/C _12734_/B _12732_/A vssd1 vssd1 vccd1 vccd1 _12737_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_29_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _12664_/Y _12666_/B vssd1 vssd1 vccd1 vccd1 _12667_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_115_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12597_ _12597_/A _12597_/B _12597_/C vssd1 vssd1 vccd1 vccd1 _12621_/A sky130_fd_sc_hd__or3_1
X_11617_ _11617_/A _11617_/B vssd1 vssd1 vccd1 vccd1 _11799_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_53_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12019__A _12096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06678__A_N _07036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11548_ _11042_/Y _11547_/X _12064_/S vssd1 vssd1 vccd1 vccd1 _11548_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_80_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11479_ _11479_/A _11479_/B _11479_/C vssd1 vssd1 vccd1 vccd1 _11480_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_110_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13218_ hold278/X _13223_/A2 _13217_/X _13223_/B2 vssd1 vssd1 vccd1 vccd1 _13219_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11184__B1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09916__A2 _11198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13149_ _13149_/A _13149_/B vssd1 vssd1 vccd1 vccd1 _13149_/Y sky130_fd_sc_hd__xnor2_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07710_ _07805_/A _07805_/B _07707_/Y vssd1 vssd1 vccd1 vccd1 _07731_/B sky130_fd_sc_hd__a21o_1
X_08690_ _08690_/A _08690_/B _08690_/C vssd1 vssd1 vccd1 vccd1 _08691_/B sky130_fd_sc_hd__and3_1
XFILLER_0_73_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07641_ _07642_/A _07642_/B vssd1 vssd1 vccd1 vccd1 _07641_/X sky130_fd_sc_hd__and2b_1
XANTENNA__12436__B1 _09149_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07572_ _07677_/A _07677_/B _07506_/X vssd1 vssd1 vccd1 vccd1 _07676_/A sky130_fd_sc_hd__a21oi_4
X_09311_ _10623_/A _09311_/B vssd1 vssd1 vccd1 vccd1 _09315_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08655__A2 _07148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10462__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09242_ _12795_/A _09242_/B vssd1 vssd1 vccd1 vccd1 _09250_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_63_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09173_ reg1_val[11] reg1_val[20] _09180_/S vssd1 vssd1 vccd1 vccd1 _09173_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09604__A1 _11752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08124_ _10092_/A _08124_/B vssd1 vssd1 vccd1 vccd1 _08131_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09080__A2 fanout86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08055_ _08085_/A _08085_/B _08050_/Y vssd1 vssd1 vccd1 vccd1 _08088_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_113_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07006_ _12642_/A _12644_/A reg1_val[2] _07248_/A vssd1 vssd1 vccd1 vccd1 _07007_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_3_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08957_ _08958_/B _08957_/B vssd1 vssd1 vccd1 vccd1 _09066_/B sky130_fd_sc_hd__and2b_1
X_07908_ _07080_/A _07080_/B _08613_/A vssd1 vssd1 vccd1 vccd1 _07910_/C sky130_fd_sc_hd__a21oi_1
X_08888_ _09836_/A _08888_/B vssd1 vssd1 vccd1 vccd1 _08890_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07839_ _09298_/B2 fanout51/X _09661_/B2 _09298_/A1 vssd1 vssd1 vccd1 vccd1 _07840_/B
+ sky130_fd_sc_hd__o22a_1
X_10850_ _11182_/A _10850_/B vssd1 vssd1 vccd1 vccd1 _10854_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11008__A _11008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12427__B1 _11892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10847__A _12093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10781_ _10539_/A _10656_/A _10656_/B vssd1 vssd1 vccd1 vccd1 _10781_/Y sky130_fd_sc_hd__a21boi_1
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09509_ _09510_/A _09510_/B vssd1 vssd1 vccd1 vccd1 _09509_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_109_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ reg1_val[9] curr_PC[9] _12520_/S vssd1 vssd1 vccd1 vccd1 _12522_/B sky130_fd_sc_hd__mux2_1
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12451_ hold175/A _12449_/X _12450_/Y vssd1 vssd1 vccd1 vccd1 _12451_/Y sky130_fd_sc_hd__a21oi_1
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11402__A1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11402_ fanout52/X fanout10/X fanout5/X _11476_/A vssd1 vssd1 vccd1 vccd1 _11403_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11402__B2 _11476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12382_ _08973_/A _06961_/X _12357_/Y _12381_/X _12631_/S vssd1 vssd1 vccd1 vccd1
+ dest_val[29] sky130_fd_sc_hd__o221a_4
XFILLER_0_50_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11333_ _11333_/A _11433_/A vssd1 vssd1 vccd1 vccd1 _11528_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_50_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11264_ _11264_/A _11264_/B _11254_/X vssd1 vssd1 vccd1 vccd1 _11265_/C sky130_fd_sc_hd__or3b_1
XFILLER_0_120_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11166__B1 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13003_ _13019_/A hold194/X vssd1 vssd1 vccd1 vccd1 hold195/A sky130_fd_sc_hd__and2_1
X_10215_ _10215_/A _10215_/B vssd1 vssd1 vccd1 vccd1 _10218_/A sky130_fd_sc_hd__xnor2_1
X_11195_ _11195_/A _11195_/B vssd1 vssd1 vccd1 vccd1 _11196_/B sky130_fd_sc_hd__xnor2_2
X_10146_ _10146_/A _10146_/B vssd1 vssd1 vccd1 vccd1 _10147_/A sky130_fd_sc_hd__nand2_2
XANTENNA__11469__A1 _11637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10077_ _10077_/A _10077_/B vssd1 vssd1 vccd1 vccd1 _10088_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08885__A2 _08112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10979_ _10980_/A _10980_/B _10980_/C vssd1 vssd1 vccd1 vccd1 _11102_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12718_ _12721_/B _12718_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[14] sky130_fd_sc_hd__and2_4
XANTENNA__10476__B _10476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09598__B1 _09422_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12649_ reg1_val[2] _12650_/B vssd1 vssd1 vccd1 vccd1 _12649_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__06970__A _11138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11944__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold305 hold305/A vssd1 vssd1 vccd1 vccd1 hold305/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13146__B2 _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09860_ _09860_/A _09860_/B vssd1 vssd1 vccd1 vccd1 _09861_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_21_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ fanout68/X _10473_/B2 _10240_/A fanout65/X vssd1 vssd1 vccd1 vccd1 _09792_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09770__B1 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08811_ _08809_/A _08809_/B _12364_/B vssd1 vssd1 vccd1 vccd1 _09040_/B sky130_fd_sc_hd__o21a_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08742_ _08741_/A _08741_/C _08741_/B vssd1 vssd1 vccd1 vccd1 _08743_/B sky130_fd_sc_hd__a21o_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08673_ _08674_/B _08723_/A _08674_/A vssd1 vssd1 vccd1 vccd1 _08725_/B sky130_fd_sc_hd__o21ba_1
XANTENNA_fanout174_A _12870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07624_ _07624_/A _07624_/B vssd1 vssd1 vccd1 vccd1 _07626_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12866__B _12870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06843__A_N _11038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12409__B1 _10788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09521__A _11770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08089__B1 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07555_ _07959_/A _07554_/B _09922_/A vssd1 vssd1 vccd1 vccd1 _07557_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07486_ _07682_/A _07682_/B _07486_/C vssd1 vssd1 vccd1 vccd1 _07490_/A sky130_fd_sc_hd__and3_1
XFILLER_0_106_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09225_ _09232_/A _09226_/B vssd1 vssd1 vccd1 vccd1 _09225_/Y sky130_fd_sc_hd__nor2_8
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08137__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07300__A2 _10473_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10199__A1 _11592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10199__B2 _10944_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09156_ _09154_/X _09155_/X _12808_/A vssd1 vssd1 vccd1 vccd1 _09156_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08107_ _10207_/A _08107_/B vssd1 vssd1 vccd1 vccd1 _08156_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09087_ _09667_/A _09087_/B vssd1 vssd1 vccd1 vccd1 _09089_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08038_ _08036_/A _08036_/B _08082_/A vssd1 vssd1 vccd1 vccd1 _08056_/B sky130_fd_sc_hd__o21a_1
X_10000_ _09707_/A _09707_/B _09862_/A _09862_/B vssd1 vssd1 vccd1 vccd1 _10000_/X
+ sky130_fd_sc_hd__o22a_1
X_09989_ _09843_/A _09843_/B _09841_/X vssd1 vssd1 vccd1 vccd1 _09991_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__08600__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09513__B1 _11198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11951_ _11952_/A _11952_/B _11952_/C vssd1 vssd1 vccd1 vccd1 _12036_/A sky130_fd_sc_hd__o21ai_1
X_11882_ _11882_/A vssd1 vssd1 vccd1 vccd1 _11883_/B sky130_fd_sc_hd__inv_2
X_10902_ _10902_/A _11122_/A vssd1 vssd1 vccd1 vccd1 _10902_/X sky130_fd_sc_hd__and2_1
XFILLER_0_39_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10833_ _10833_/A _10834_/B vssd1 vssd1 vccd1 vccd1 _10972_/A sky130_fd_sc_hd__nor2_1
X_10764_ _10765_/A _10765_/B vssd1 vssd1 vccd1 vccd1 _10764_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_94_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12503_ _12504_/A _12504_/B _12504_/C vssd1 vssd1 vccd1 vccd1 _12511_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_13_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10695_ _10165_/S _10025_/Y _09251_/A vssd1 vssd1 vccd1 vccd1 _10695_/Y sky130_fd_sc_hd__o21ai_2
X_12434_ _12390_/A _12389_/A _12434_/S vssd1 vssd1 vccd1 vccd1 _12435_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11926__A2 _07316_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12365_ _12365_/A _12365_/B _12365_/C vssd1 vssd1 vccd1 vccd1 _12381_/B sky130_fd_sc_hd__and3_1
X_11316_ _11076_/A _11076_/B _11194_/B _11195_/B _11195_/A vssd1 vssd1 vccd1 vccd1
+ _11318_/C sky130_fd_sc_hd__a32oi_2
XFILLER_0_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12296_ _12296_/A _12296_/B _12296_/C vssd1 vssd1 vccd1 vccd1 _12297_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11247_ _11247_/A _11247_/B _11247_/C vssd1 vssd1 vccd1 vccd1 _11247_/X sky130_fd_sc_hd__and3_1
XANTENNA__07358__A2 _12779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ _11179_/A _11179_/B vssd1 vssd1 vccd1 vccd1 _11180_/A sky130_fd_sc_hd__and2_1
XFILLER_0_38_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11347__S _11813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10129_ _09992_/A _09992_/B _09990_/Y vssd1 vssd1 vccd1 vccd1 _10130_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__09325__B _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08307__B2 _08540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08307__A1 _08515_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10114__B2 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10114__A1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06965__A _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09341__A _09341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11082__S _11179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10417__A2 _10453_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07340_ _07340_/A _07340_/B vssd1 vssd1 vccd1 vccd1 _07342_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07271_ _11080_/A _11081_/A _11179_/A vssd1 vssd1 vccd1 vccd1 _07271_/X sky130_fd_sc_hd__mux2_1
X_09010_ _09010_/A _11946_/C vssd1 vssd1 vccd1 vccd1 _09010_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_26_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11378__B1 _07608_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07796__A _09341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08243__B1 _08457_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold124 hold124/A vssd1 vssd1 vccd1 vccd1 hold124/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 hold113/A vssd1 vssd1 vccd1 vccd1 hold113/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 hold102/A vssd1 vssd1 vccd1 vccd1 hold102/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 hold152/X vssd1 vssd1 vccd1 vccd1 hold135/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07597__A2 _07362_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold168 hold168/A vssd1 vssd1 vccd1 vccd1 hold168/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 hold146/A vssd1 vssd1 vccd1 vccd1 hold146/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 hold157/A vssd1 vssd1 vccd1 vccd1 hold157/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold179 hold179/A vssd1 vssd1 vccd1 vccd1 hold179/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10950__A _10950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09912_ _09856_/A _09856_/B _09857_/Y vssd1 vssd1 vccd1 vccd1 _09998_/A sky130_fd_sc_hd__o21ai_4
X_09843_ _09843_/A _09843_/B vssd1 vssd1 vccd1 vccd1 _09845_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09516__A _09834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07036__A _07036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06986_ _07036_/A _07014_/A _06986_/C vssd1 vssd1 vccd1 vccd1 _07048_/B sky130_fd_sc_hd__nand3_2
X_09774_ _09775_/B _09774_/B vssd1 vssd1 vccd1 vccd1 _09776_/A sky130_fd_sc_hd__and2b_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08725_ _08725_/A _08725_/B vssd1 vssd1 vccd1 vccd1 _10287_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08656_ _08656_/A _08656_/B vssd1 vssd1 vccd1 vccd1 _08661_/A sky130_fd_sc_hd__xnor2_2
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07607_ _07608_/A _07608_/B vssd1 vssd1 vccd1 vccd1 _12335_/A sky130_fd_sc_hd__and2_4
XFILLER_0_49_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08587_ _08587_/A _08587_/B vssd1 vssd1 vccd1 vccd1 _08592_/B sky130_fd_sc_hd__xor2_1
XANTENNA__07521__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07538_ _07537_/B _07537_/C _07537_/A vssd1 vssd1 vccd1 vccd1 _07559_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_76_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07469_ _07469_/A _07469_/B vssd1 vssd1 vccd1 vccd1 _07492_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10480_ _10479_/B _10479_/C _10479_/A vssd1 vssd1 vccd1 vccd1 _10481_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_63_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09208_ reg1_val[10] reg1_val[21] _09211_/S vssd1 vssd1 vccd1 vccd1 _09208_/X sky130_fd_sc_hd__mux2_1
X_09139_ _09139_/A _09139_/B vssd1 vssd1 vccd1 vccd1 _09141_/B sky130_fd_sc_hd__xnor2_2
X_12150_ _09149_/Y _12122_/Y _12123_/X _12127_/X _12149_/X vssd1 vssd1 vccd1 vccd1
+ _12150_/X sky130_fd_sc_hd__a311o_1
X_11101_ _10984_/B _10984_/C _10984_/A vssd1 vssd1 vccd1 vccd1 _11111_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_102_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10860__A _12157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12081_ _12631_/S _12077_/X _12078_/X _12080_/Y vssd1 vssd1 vccd1 vccd1 dest_val[24]
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12333__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11032_ hold198/A _11032_/B vssd1 vssd1 vccd1 vccd1 _11147_/B sky130_fd_sc_hd__or2_1
XANTENNA__09145__B _09146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07760__A2 _08484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12983_ _13001_/A hold240/X vssd1 vssd1 vccd1 vccd1 _13301_/D sky130_fd_sc_hd__and2_1
X_11934_ _12012_/B _11934_/B vssd1 vssd1 vccd1 vccd1 _11936_/B sky130_fd_sc_hd__or2_1
XFILLER_0_99_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13046__B1 _13254_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11865_ _12335_/B _11865_/B vssd1 vssd1 vccd1 vccd1 _11867_/B sky130_fd_sc_hd__xnor2_1
X_11796_ _11797_/A _11797_/B _11797_/C vssd1 vssd1 vccd1 vccd1 _11796_/X sky130_fd_sc_hd__a21o_1
X_10816_ _10806_/Y _10807_/X _11733_/B _10159_/A _10814_/X vssd1 vssd1 vccd1 vccd1
+ _10816_/X sky130_fd_sc_hd__o221a_1
XANTENNA__09265__A2 _07362_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10747_ _11179_/A _10747_/B vssd1 vssd1 vccd1 vccd1 _10749_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10678_ _10679_/A _10679_/B _10679_/C vssd1 vssd1 vccd1 vccd1 _10678_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_4_11_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12417_ hold241/A _12417_/B vssd1 vssd1 vccd1 vccd1 _12417_/X sky130_fd_sc_hd__or2_1
XFILLER_0_70_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13397_ _13398_/CLK hold4/X vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10032__B1 _09257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10583__B2 _10974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10583__A1 _11093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12348_ _12348_/A _12348_/B vssd1 vssd1 vccd1 vccd1 _12429_/A sky130_fd_sc_hd__or2_2
X_12279_ _12252_/X _12256_/X _12278_/X _12220_/X _12631_/S vssd1 vssd1 vccd1 vccd1
+ dest_val[27] sky130_fd_sc_hd__o32a_4
XANTENNA__08528__A1 _06992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08528__B2 _08613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06679__B _07036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10335__A1 _10599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10335__B2 _10500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06840_ _06754_/X _06838_/Y _06839_/X vssd1 vssd1 vccd1 vccd1 _06840_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06771_ reg2_val[7] _06810_/B vssd1 vssd1 vccd1 vccd1 _06771_/X sky130_fd_sc_hd__and2_2
XANTENNA__11835__B2 _10788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09490_ _10623_/A _09490_/B vssd1 vssd1 vccd1 vccd1 _09494_/A sky130_fd_sc_hd__xnor2_1
X_08510_ _08527_/A _08509_/Y _08505_/X vssd1 vssd1 vccd1 vccd1 _08518_/A sky130_fd_sc_hd__o21a_1
XANTENNA__09071__A _09944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08441_ _08564_/A _08441_/B vssd1 vssd1 vccd1 vccd1 _08447_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08372_ _08375_/A _08375_/B vssd1 vssd1 vccd1 vccd1 _08372_/X sky130_fd_sc_hd__or2_1
XANTENNA__10945__A _12224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11063__A2 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07323_ _07323_/A _07323_/B vssd1 vssd1 vccd1 vccd1 _07325_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11540__S _11813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07254_ _10749_/A _07254_/B vssd1 vssd1 vccd1 vccd1 _07255_/B sky130_fd_sc_hd__or2_1
XANTENNA_fanout137_A _10207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07185_ reg1_val[11] reg1_val[12] reg1_val[13] _07248_/B _07585_/B1 vssd1 vssd1 vccd1
+ vccd1 _07265_/B sky130_fd_sc_hd__o41a_1
XFILLER_0_41_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11771__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06793__A3 _12665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09826_ _09827_/A _09827_/B vssd1 vssd1 vccd1 vccd1 _09826_/Y sky130_fd_sc_hd__nor2_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06969_ _12438_/A _07147_/B vssd1 vssd1 vccd1 vccd1 _06969_/Y sky130_fd_sc_hd__nand2_2
X_09757_ _09221_/Y _09732_/B _12319_/B _12379_/B2 _09756_/X vssd1 vssd1 vccd1 vccd1
+ _09757_/X sky130_fd_sc_hd__a221o_1
X_08708_ _08708_/A _08708_/B vssd1 vssd1 vccd1 vccd1 _08920_/B sky130_fd_sc_hd__xnor2_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _09688_/A _09688_/B vssd1 vssd1 vccd1 vccd1 _09689_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13028__B1 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _08638_/B _08646_/A _08638_/A vssd1 vssd1 vccd1 vccd1 _08674_/B sky130_fd_sc_hd__a21oi_1
X_11650_ hold262/A _11650_/B _11739_/B vssd1 vssd1 vccd1 vccd1 _11650_/Y sky130_fd_sc_hd__nand3_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout30 _07218_/X vssd1 vssd1 vccd1 vccd1 fanout30/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_49_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11581_ _11582_/A _11582_/B vssd1 vssd1 vccd1 vccd1 _11692_/A sky130_fd_sc_hd__or2_1
X_10601_ _11671_/A fanout47/X fanout45/X fanout52/X vssd1 vssd1 vccd1 vccd1 _10602_/B
+ sky130_fd_sc_hd__o22a_1
Xfanout74 fanout75/X vssd1 vssd1 vccd1 vccd1 fanout74/X sky130_fd_sc_hd__buf_6
Xfanout63 _07014_/Y vssd1 vssd1 vccd1 vccd1 fanout63/X sky130_fd_sc_hd__buf_6
Xfanout41 fanout42/X vssd1 vssd1 vccd1 vccd1 fanout41/X sky130_fd_sc_hd__clkbuf_8
Xfanout52 _07079_/X vssd1 vssd1 vccd1 vccd1 fanout52/X sky130_fd_sc_hd__buf_4
XANTENNA__08455__B1 _09770_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13320_ _13373_/CLK hold203/X vssd1 vssd1 vccd1 vccd1 hold201/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10532_ _10532_/A _10532_/B vssd1 vssd1 vccd1 vccd1 _10534_/B sky130_fd_sc_hd__xnor2_2
Xfanout96 _09834_/A vssd1 vssd1 vccd1 vccd1 _11393_/A sky130_fd_sc_hd__buf_4
XFILLER_0_52_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout85 _07257_/X vssd1 vssd1 vccd1 vccd1 _11309_/A sky130_fd_sc_hd__buf_6
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10463_ _11182_/A _10463_/B vssd1 vssd1 vccd1 vccd1 _10464_/B sky130_fd_sc_hd__xnor2_1
X_13251_ hold140/X _12804_/A _13039_/A hold141/X vssd1 vssd1 vccd1 vccd1 hold142/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12202_ _12202_/A _12202_/B vssd1 vssd1 vccd1 vccd1 _12211_/B sky130_fd_sc_hd__nor2_1
X_13182_ _13210_/A _13182_/B vssd1 vssd1 vccd1 vccd1 _13377_/D sky130_fd_sc_hd__and2_1
XFILLER_0_103_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10394_ _10395_/A _10395_/B _10395_/C vssd1 vssd1 vccd1 vccd1 _10394_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10590__A _12096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12133_ _12131_/Y _12133_/B vssd1 vssd1 vccd1 vccd1 _12134_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_20_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12064_ _10293_/X _12063_/Y _12064_/S vssd1 vssd1 vccd1 vccd1 _12064_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11015_ _10937_/X _11050_/D _12356_/B1 vssd1 vssd1 vccd1 vccd1 _11015_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10317__A1 _12365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08995__A _11844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08930__B2 _07134_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08930__A1 _07121_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_max_cap102_A _07983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12966_ _12876_/X _12966_/B vssd1 vssd1 vccd1 vccd1 _13234_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09486__A2 _10245_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11293__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11917_ _11911_/Y _11912_/X _11916_/X vssd1 vssd1 vccd1 vccd1 _11917_/X sky130_fd_sc_hd__o21ba_1
X_12897_ hold294/A hold22/X vssd1 vssd1 vccd1 vccd1 _13148_/A sky130_fd_sc_hd__nand2b_1
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ _11848_/A _11848_/B vssd1 vssd1 vccd1 vccd1 _11849_/B sky130_fd_sc_hd__or2_1
XFILLER_0_74_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11779_ _11779_/A _12428_/B vssd1 vssd1 vccd1 vccd1 _11781_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08990_ _08876_/A _11946_/C _12385_/B vssd1 vssd1 vccd1 vccd1 _08990_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07941_ _07941_/A _07941_/B vssd1 vssd1 vccd1 vccd1 _07953_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__10859__A2 _07362_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07872_ _07872_/A _07872_/B vssd1 vssd1 vccd1 vccd1 _07880_/B sky130_fd_sc_hd__xnor2_2
X_06823_ reg1_val[3] _11138_/A vssd1 vssd1 vccd1 vccd1 _06823_/X sky130_fd_sc_hd__and2_1
X_09611_ _09614_/A vssd1 vssd1 vccd1 vccd1 _09611_/Y sky130_fd_sc_hd__inv_2
X_06754_ _10808_/S _06754_/B vssd1 vssd1 vccd1 vccd1 _06754_/X sky130_fd_sc_hd__or2_1
X_09542_ _09542_/A _09542_/B vssd1 vssd1 vccd1 vccd1 _09544_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_78_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10659__B _10779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06685_ reg1_val[22] _07014_/A vssd1 vssd1 vccd1 vccd1 _06686_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09473_ _09822_/A _08877_/B fanout6/X _09677_/A vssd1 vssd1 vccd1 vccd1 _09474_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07488__A1 _07148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07488__B2 _07959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10492__B1 _07269_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09229__A2 _12420_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08424_ _08424_/A _08424_/B vssd1 vssd1 vccd1 vccd1 _08425_/B sky130_fd_sc_hd__and2_1
XFILLER_0_19_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08355_ _08355_/A _08355_/B vssd1 vssd1 vccd1 vccd1 _08365_/B sky130_fd_sc_hd__xor2_2
XANTENNA__10244__B1 _10243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08988__A1 _12438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07306_ _07306_/A _07306_/B vssd1 vssd1 vccd1 vccd1 _07413_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08145__A _08454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06999__B1 _06993_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08286_ _08286_/A _08286_/B vssd1 vssd1 vccd1 vccd1 _08320_/A sky130_fd_sc_hd__xnor2_1
X_07237_ _07237_/A _07238_/B vssd1 vssd1 vccd1 vccd1 _07237_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_33_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07168_ _07168_/A _07168_/B _07168_/C vssd1 vssd1 vccd1 vccd1 _07170_/A sky130_fd_sc_hd__and3_1
XFILLER_0_42_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07963__A2 _08112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07099_ _09661_/B2 _10245_/B2 fanout98/X _10245_/A1 vssd1 vssd1 vccd1 vccd1 _07100_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout231 _06617_/Y vssd1 vssd1 vccd1 vccd1 _06677_/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout220 _07172_/A vssd1 vssd1 vccd1 vccd1 _10294_/S sky130_fd_sc_hd__clkbuf_4
Xfanout264 _12796_/A vssd1 vssd1 vccd1 vccd1 _12639_/A sky130_fd_sc_hd__clkbuf_8
Xfanout253 _06577_/Y vssd1 vssd1 vccd1 vccd1 _13094_/A2 sky130_fd_sc_hd__buf_4
Xfanout242 _12471_/S vssd1 vssd1 vccd1 vccd1 _10821_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__07176__B1 _07173_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout275 _13162_/A vssd1 vssd1 vccd1 vccd1 _13019_/A sky130_fd_sc_hd__buf_2
Xfanout286 _06584_/Y vssd1 vssd1 vccd1 vccd1 _12404_/S sky130_fd_sc_hd__clkbuf_8
X_09809_ _11182_/A _09809_/B vssd1 vssd1 vccd1 vccd1 _09811_/B sky130_fd_sc_hd__xnor2_1
X_12820_ hold18/X _12820_/B vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__or2_1
XANTENNA__09423__B _12359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07224__A _09836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12751_ _12751_/A _12751_/B vssd1 vssd1 vccd1 vccd1 _12760_/C sky130_fd_sc_hd__nand2_4
X_11702_ _11703_/A _11703_/B vssd1 vssd1 vccd1 vccd1 _11797_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_96_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12682_ _12682_/A _12682_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[8] sky130_fd_sc_hd__xor2_4
X_11633_ _11541_/A _11539_/Y _11553_/S vssd1 vssd1 vccd1 vccd1 _11634_/B sky130_fd_sc_hd__o21ba_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11564_ curr_PC[18] _11564_/B vssd1 vssd1 vccd1 vccd1 _11749_/C sky130_fd_sc_hd__and2_2
XFILLER_0_37_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11495_ _12336_/A _11495_/B vssd1 vssd1 vccd1 vccd1 _11503_/A sky130_fd_sc_hd__xnor2_2
X_10515_ _10515_/A _10515_/B vssd1 vssd1 vccd1 vccd1 _10516_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_80_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13303_ _13304_/CLK _13303_/D vssd1 vssd1 vccd1 vccd1 hold211/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13234_ _13234_/A _13234_/B vssd1 vssd1 vccd1 vccd1 _13234_/Y sky130_fd_sc_hd__xnor2_1
X_10446_ _09242_/B _10433_/X _10445_/X _10424_/X vssd1 vssd1 vccd1 vccd1 _10446_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07894__A _09836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13165_ hold285/A _13164_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13165_/X sky130_fd_sc_hd__mux2_1
X_10377_ _10525_/A _10377_/B vssd1 vssd1 vccd1 vccd1 _10379_/B sky130_fd_sc_hd__or2_1
X_12116_ _11964_/A _12039_/Y _12041_/B vssd1 vssd1 vccd1 vccd1 _12116_/Y sky130_fd_sc_hd__a21oi_1
X_13096_ hold57/X _06577_/A _13254_/A2 hold6/X rst vssd1 vssd1 vccd1 vccd1 _13096_/X
+ sky130_fd_sc_hd__a221o_1
X_12047_ _11340_/B _11713_/Y _12043_/A _12043_/B _12046_/X vssd1 vssd1 vccd1 vccd1
+ _12048_/B sky130_fd_sc_hd__a41o_1
XANTENNA__11355__S _12064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12949_ _13198_/A _12948_/B _12886_/X vssd1 vssd1 vccd1 vccd1 _13203_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_87_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12975__A _13001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08667__A0 _08658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06692__B _07016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08140_ _08140_/A _08140_/B vssd1 vssd1 vccd1 vccd1 _08217_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09631__A2 _07262_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11974__B1 _09150_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08071_ _08170_/A _08170_/B vssd1 vssd1 vccd1 vccd1 _08072_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_70_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07022_ _09947_/A _07022_/B vssd1 vssd1 vccd1 vccd1 _07041_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13191__A2 _13223_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06602__C1 _06675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08973_ _08973_/A _08973_/B _08973_/C _08973_/D vssd1 vssd1 vccd1 vccd1 _08973_/X
+ sky130_fd_sc_hd__or4_2
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07924_ _07924_/A _07924_/B vssd1 vssd1 vccd1 vccd1 _07927_/B sky130_fd_sc_hd__xor2_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08370__A2 _10221_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07855_ _07861_/B _07861_/A vssd1 vssd1 vccd1 vccd1 _07855_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_127_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06806_ reg1_val[2] _07172_/A vssd1 vssd1 vccd1 vccd1 _06809_/A sky130_fd_sc_hd__nand2_1
X_07786_ _10207_/A _07786_/B vssd1 vssd1 vccd1 vccd1 _07790_/A sky130_fd_sc_hd__xnor2_1
X_06737_ _11134_/A _07270_/A vssd1 vssd1 vccd1 vccd1 _11150_/S sky130_fd_sc_hd__and2_1
XANTENNA__12454__B2 _09221_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09525_ _09525_/A _09525_/B vssd1 vssd1 vccd1 vccd1 _09527_/B sky130_fd_sc_hd__xor2_1
XANTENNA__07044__A _07604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06668_ _07046_/B reg1_val[26] vssd1 vssd1 vccd1 vccd1 _12207_/S sky130_fd_sc_hd__and2b_1
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09456_ _09779_/A _09456_/B vssd1 vssd1 vccd1 vccd1 _09457_/B sky130_fd_sc_hd__xor2_1
X_08407_ _08407_/A _08407_/B vssd1 vssd1 vccd1 vccd1 _08435_/A sky130_fd_sc_hd__xor2_1
X_06599_ instruction[19] _06944_/B vssd1 vssd1 vccd1 vccd1 _06599_/X sky130_fd_sc_hd__or2_1
X_09387_ _09173_/X _09176_/X _09403_/S vssd1 vssd1 vccd1 vccd1 _09387_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08338_ _09670_/A _08338_/B vssd1 vssd1 vccd1 vccd1 _08342_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08269_ _08269_/A _08269_/B vssd1 vssd1 vccd1 vccd1 _08270_/B sky130_fd_sc_hd__nand2_1
X_11280_ _11389_/A _11280_/B vssd1 vssd1 vccd1 vccd1 _11282_/B sky130_fd_sc_hd__nand2_1
X_10300_ hold211/A _10300_/B vssd1 vssd1 vccd1 vccd1 _10434_/B sky130_fd_sc_hd__or2_1
XFILLER_0_61_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10231_ _11398_/A _10231_/B vssd1 vssd1 vccd1 vccd1 _10233_/B sky130_fd_sc_hd__xor2_1
XANTENNA__08189__A2 _10221_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10162_ _10160_/X _10161_/X _11246_/S vssd1 vssd1 vccd1 vccd1 _10162_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10940__B2 _11764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10940__A1 _11779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10093_ _11671_/A fanout28/X fanout26/X fanout52/X vssd1 vssd1 vccd1 vccd1 _10094_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12142__B1 _12205_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12779__B _12779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11496__A2 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07164__A3 _07959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12803_ rst _12803_/B _12803_/C vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__nor3_1
XANTENNA__12795__A _12795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08649__B1 _08649_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10995_ _10995_/A _10995_/B vssd1 vssd1 vccd1 vccd1 _10997_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10456__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12996__A2 _13000_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12734_ _12739_/C _12734_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[18] sky130_fd_sc_hd__xor2_4
XANTENNA__09310__B2 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08113__A2 _08199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09310__A1 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ reg1_val[5] _12665_/B vssd1 vssd1 vccd1 vccd1 _12666_/B sky130_fd_sc_hd__nand2_1
X_11616_ _11616_/A _11616_/B _11616_/C vssd1 vssd1 vccd1 vccd1 _11617_/B sky130_fd_sc_hd__nand3_1
X_12596_ _12596_/A _12596_/B vssd1 vssd1 vccd1 vccd1 _12611_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_108_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10208__B1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11547_ _11547_/A _11547_/B vssd1 vssd1 vccd1 vccd1 _11547_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_4_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11478_ _11479_/A _11479_/B _11479_/C vssd1 vssd1 vccd1 vccd1 _11600_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_52_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09377__A1 _10049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13217_ hold254/X _13216_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13217_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11184__A1 _11946_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10429_ _10429_/A _10429_/B vssd1 vssd1 vccd1 vccd1 _10429_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__11184__B2 _07013_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13148_ _13148_/A _13148_/B vssd1 vssd1 vccd1 vccd1 _13149_/B sky130_fd_sc_hd__nand2_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10931__B2 _12379_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ _07212_/C _13089_/A2 hold104/X vssd1 vssd1 vccd1 vccd1 hold105/A sky130_fd_sc_hd__o21a_1
XANTENNA__06968__A _12438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12689__B _12689_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07640_ _08893_/B _07640_/B vssd1 vssd1 vccd1 vccd1 _07642_/B sky130_fd_sc_hd__and2_1
X_07571_ _07571_/A _07571_/B vssd1 vssd1 vccd1 vccd1 _07677_/B sky130_fd_sc_hd__xor2_4
XANTENNA__11813__S _11813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09310_ fanout61/X fanout86/X fanout82/X fanout53/X vssd1 vssd1 vccd1 vccd1 _09311_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11644__C1 _09242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09241_ _09241_/A _09241_/B vssd1 vssd1 vccd1 vccd1 _09241_/X sky130_fd_sc_hd__or2_1
XFILLER_0_113_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09172_ reg1_val[10] reg1_val[21] _09180_/S vssd1 vssd1 vccd1 vccd1 _09172_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08123_ _08649_/B1 _08199_/B fanout33/X _09404_/S vssd1 vssd1 vccd1 vccd1 _08124_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08054_ _08054_/A vssd1 vssd1 vccd1 vccd1 _08085_/B sky130_fd_sc_hd__inv_2
XFILLER_0_113_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07005_ _09947_/A vssd1 vssd1 vccd1 vccd1 _09302_/A sky130_fd_sc_hd__inv_6
XFILLER_0_31_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10164__S _11138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12372__B1 _11648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10922__A1 _11990_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ _10479_/A _08956_/B vssd1 vssd1 vccd1 vccd1 _08958_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06597__B _06944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07907_ _12642_/A _07907_/B _07907_/C vssd1 vssd1 vccd1 vccd1 _07910_/B sky130_fd_sc_hd__and3_1
X_08887_ _07959_/B _07232_/X _07238_/Y fanout29/X vssd1 vssd1 vccd1 vccd1 _08888_/B
+ sky130_fd_sc_hd__a22o_1
X_07838_ _07837_/A _07837_/B _07837_/C vssd1 vssd1 vccd1 vccd1 _07841_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12978__A2 _13000_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09508_ _09508_/A _09508_/B vssd1 vssd1 vccd1 vccd1 _09510_/B sky130_fd_sc_hd__xnor2_1
X_07769_ _09834_/A _07769_/B vssd1 vssd1 vccd1 vccd1 _07781_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10780_ _10780_/A _11009_/A vssd1 vssd1 vccd1 vccd1 _10780_/X sky130_fd_sc_hd__and2_1
XFILLER_0_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout32_A _07213_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _10159_/A _12412_/B _09433_/Y _09429_/X vssd1 vssd1 vccd1 vccd1 _09439_/X
+ sky130_fd_sc_hd__o211a_1
X_12450_ hold175/A _12449_/X _09238_/Y vssd1 vssd1 vccd1 vccd1 _12450_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11401_ _11401_/A _11401_/B vssd1 vssd1 vccd1 vccd1 _11410_/B sky130_fd_sc_hd__or2_1
XFILLER_0_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11402__A2 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12381_ _12381_/A _12381_/B _12381_/C _12369_/X vssd1 vssd1 vccd1 vccd1 _12381_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_104_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11332_ _11330_/Y _11332_/B vssd1 vssd1 vccd1 vccd1 _11526_/A sky130_fd_sc_hd__nand2b_2
XANTENNA__08333__A _08564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11166__A1 _11779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11263_ _09222_/Y _11249_/B _11262_/X _12379_/B2 vssd1 vssd1 vccd1 vccd1 _11264_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_120_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11194_ _11194_/A _11194_/B vssd1 vssd1 vccd1 vccd1 _11195_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11166__B2 _11764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13002_ _13310_/Q _13171_/B2 _13209_/A2 hold193/X vssd1 vssd1 vccd1 vccd1 hold194/A
+ sky130_fd_sc_hd__a22o_1
X_10214_ _11179_/A _10214_/B vssd1 vssd1 vccd1 vccd1 _10215_/B sky130_fd_sc_hd__xnor2_1
X_10145_ _09554_/B _10138_/C _10143_/Y _10661_/A vssd1 vssd1 vccd1 vccd1 _10146_/B
+ sky130_fd_sc_hd__o211ai_2
X_10076_ _10224_/A _10076_/B vssd1 vssd1 vccd1 vccd1 _10077_/B sky130_fd_sc_hd__or2_1
XANTENNA__12418__A1 _12447_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10978_ _10848_/A _10848_/B _10845_/A vssd1 vssd1 vccd1 vccd1 _10983_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08508__A _08658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12717_ _12717_/A _12717_/B _12717_/C vssd1 vssd1 vccd1 vccd1 _12718_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_128_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10476__C _10476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12648_ _12647_/A _12647_/B _12646_/B vssd1 vssd1 vccd1 vccd1 _12652_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_115_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12579_ _12633_/A _12580_/B vssd1 vssd1 vccd1 vccd1 _12598_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_108_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12464__S _12471_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06970__B _10297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10601__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold306 hold306/A vssd1 vssd1 vccd1 vccd1 hold306/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09339__A _09834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13146__A2 _12803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09770__A1 _07217_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08810_ _09040_/A _08810_/B vssd1 vssd1 vccd1 vccd1 _08810_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _09790_/A _09790_/B vssd1 vssd1 vccd1 vccd1 _09831_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09770__B2 _09770_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08741_ _08741_/A _08741_/B _08741_/C vssd1 vssd1 vccd1 vccd1 _08743_/A sky130_fd_sc_hd__nand3_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08672_ _08645_/X _08721_/A _08671_/B vssd1 vssd1 vccd1 vccd1 _08723_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09802__A _11582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07623_ _07624_/B _07624_/A vssd1 vssd1 vccd1 vccd1 _07623_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_17_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08089__B2 _08613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08089__A1 _06992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07554_ _07959_/A _07554_/B _07706_/B vssd1 vssd1 vccd1 vccd1 _07557_/B sky130_fd_sc_hd__and3_1
XANTENNA__08418__A _08575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07485_ _09834_/A _07485_/B vssd1 vssd1 vccd1 vccd1 _07486_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09224_ _09237_/B _09228_/B vssd1 vssd1 vccd1 vccd1 _09224_/X sky130_fd_sc_hd__or2_1
XANTENNA__11779__A _11779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10199__A2 _07213_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09155_ _09218_/A reg1_val[31] _09180_/S vssd1 vssd1 vccd1 vccd1 _09155_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09249__A _11138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08106_ _08561_/A2 _10476_/A _09940_/B2 _08411_/B vssd1 vssd1 vccd1 vccd1 _08107_/B
+ sky130_fd_sc_hd__o22a_1
X_09086_ _09661_/B2 fanout78/X fanout74/X fanout98/X vssd1 vssd1 vccd1 vccd1 _09087_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08037_ _08081_/A _08081_/B vssd1 vssd1 vccd1 vccd1 _08082_/A sky130_fd_sc_hd__or2_1
XFILLER_0_101_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09988_ _09831_/A _09831_/B _09829_/Y vssd1 vssd1 vccd1 vccd1 _09991_/A sky130_fd_sc_hd__a21oi_4
X_08939_ _08939_/A _08939_/B vssd1 vssd1 vccd1 vccd1 _08941_/B sky130_fd_sc_hd__xnor2_1
X_11950_ _11950_/A _11950_/B vssd1 vssd1 vccd1 vccd1 _11952_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09513__B2 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09513__A1 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10901_ _10658_/X _11122_/A _10899_/Y vssd1 vssd1 vccd1 vccd1 _10901_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07524__B1 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11881_ _11881_/A _11881_/B _11881_/C vssd1 vssd1 vccd1 vccd1 _11882_/A sky130_fd_sc_hd__and3_1
XFILLER_0_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10832_ _10950_/A _07255_/B fanout8/A _10831_/Y vssd1 vssd1 vccd1 vccd1 _10834_/B
+ sky130_fd_sc_hd__o31ai_2
XANTENNA__13073__A1 _11182_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10763_ _10616_/A _10707_/A _10619_/A vssd1 vssd1 vccd1 vccd1 _10765_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07232__A _07233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10831__B1 _10950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12502_ _12511_/A _12502_/B vssd1 vssd1 vccd1 vccd1 _12504_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_82_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10694_ _10686_/Y _10687_/X _10692_/X _10693_/Y vssd1 vssd1 vccd1 vccd1 _10694_/X
+ sky130_fd_sc_hd__o211a_1
X_12433_ _12433_/A _12433_/B vssd1 vssd1 vccd1 vccd1 _12435_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12364_ _12364_/A _12364_/B _08810_/Y vssd1 vssd1 vccd1 vccd1 _12365_/C sky130_fd_sc_hd__or3b_1
XFILLER_0_1_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11315_ _11199_/A _11199_/B _11202_/A vssd1 vssd1 vccd1 vccd1 _11320_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_50_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12295_ _12296_/A _12296_/B _12296_/C vssd1 vssd1 vccd1 vccd1 _12298_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__09201__A0 _11134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11246_ _10295_/X _10297_/X _11246_/S vssd1 vssd1 vccd1 vccd1 _11246_/X sky130_fd_sc_hd__mux2_1
X_11177_ _11582_/A _11177_/B vssd1 vssd1 vccd1 vccd1 _11179_/B sky130_fd_sc_hd__xnor2_1
X_10128_ _10128_/A _10128_/B vssd1 vssd1 vccd1 vccd1 _10130_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__07407__A _09672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10059_ _07298_/Y _10476_/B _10476_/C _10240_/A _12233_/B vssd1 vssd1 vccd1 vccd1
+ _10060_/B sky130_fd_sc_hd__o32a_1
XANTENNA__09504__A1 _09673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08307__A2 _08561_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10114__A2 _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12272__C1 _12376_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12811__A1 _07148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07270_ _07270_/A _07270_/B vssd1 vssd1 vccd1 vccd1 _07270_/X sky130_fd_sc_hd__xor2_4
XANTENNA__12983__A _13001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06981__A _07078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11378__A1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11378__B2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08243__A1 _08641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08243__B2 _08627_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold103 hold103/A vssd1 vssd1 vccd1 vccd1 hold103/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 hold114/A vssd1 vssd1 vccd1 vccd1 hold114/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 hold125/A vssd1 vssd1 vccd1 vccd1 hold125/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12327__B1 _12421_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold136 hold136/A vssd1 vssd1 vccd1 vccd1 hold136/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 hold158/A vssd1 vssd1 vccd1 vccd1 hold158/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 hold147/A vssd1 vssd1 vccd1 vccd1 hold147/X sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _09861_/A _09861_/B _09859_/X vssd1 vssd1 vccd1 vccd1 _09999_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_1_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold169 hold198/X vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12223__A _12224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09842_ _09842_/A _09842_/B vssd1 vssd1 vccd1 vccd1 _09843_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09773_ _09922_/A _09773_/B vssd1 vssd1 vccd1 vccd1 _09774_/B sky130_fd_sc_hd__xor2_1
XANTENNA__07317__A _10476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06985_ _07036_/A _07014_/A _06986_/C vssd1 vssd1 vccd1 vccd1 _06987_/B sky130_fd_sc_hd__and3_1
XANTENNA_fanout284_A _12054_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08724_ _10151_/B _10151_/C vssd1 vssd1 vccd1 vccd1 _10287_/B sky130_fd_sc_hd__and2_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ _07983_/A _07148_/Y _07173_/Y _09218_/A vssd1 vssd1 vccd1 vccd1 _08656_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07606_ _07094_/B _07315_/A _07315_/B _08973_/A vssd1 vssd1 vccd1 vccd1 _07608_/B
+ sky130_fd_sc_hd__o211ai_4
X_08586_ _08584_/Y _08605_/B _08571_/Y vssd1 vssd1 vccd1 vccd1 _08592_/A sky130_fd_sc_hd__o21ai_1
X_07537_ _07537_/A _07537_/B _07537_/C vssd1 vssd1 vccd1 vccd1 _07737_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_64_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07987__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07468_ _07468_/A _07468_/B vssd1 vssd1 vccd1 vccd1 _07469_/B sky130_fd_sc_hd__and2_1
XFILLER_0_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11369__A1 _09225_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09207_ reg1_val[11] reg1_val[20] _09211_/S vssd1 vssd1 vccd1 vccd1 _09207_/X sky130_fd_sc_hd__mux2_1
X_07399_ _07400_/B _07435_/A _07400_/A vssd1 vssd1 vccd1 vccd1 _07401_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_72_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09138_ _09025_/A _09025_/B _09023_/Y vssd1 vssd1 vccd1 vccd1 _09139_/B sky130_fd_sc_hd__a21oi_4
X_11100_ _11100_/A _11100_/B vssd1 vssd1 vccd1 vccd1 _11113_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_32_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09069_ _09069_/A _09069_/B vssd1 vssd1 vccd1 vccd1 _09112_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__12869__A1 _08859_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12080_ _12631_/S _12216_/C vssd1 vssd1 vccd1 vccd1 _12080_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09707__A _09707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11031_ _12412_/A _11027_/X _11030_/Y _12446_/C1 vssd1 vssd1 vccd1 vccd1 _11031_/X
+ sky130_fd_sc_hd__o211a_1
X_12982_ hold221/X _13000_/A2 _13257_/A2 hold239/X vssd1 vssd1 vccd1 vccd1 hold240/A
+ sky130_fd_sc_hd__a22o_1
X_11933_ _11932_/B _11933_/B vssd1 vssd1 vccd1 vccd1 _11934_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_99_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11864_ _12009_/A fanout10/X fanout5/X fanout58/X vssd1 vssd1 vccd1 vccd1 _11865_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11057__B1 _11058_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10815_ _11247_/A _09885_/X _09251_/A vssd1 vssd1 vccd1 vccd1 _11733_/B sky130_fd_sc_hd__o21ai_2
X_11795_ _11797_/A _11797_/B _11797_/C vssd1 vssd1 vccd1 vccd1 _11798_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10746_ fanout75/X fanout17/X fanout14/X _08289_/B vssd1 vssd1 vccd1 vccd1 _10747_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_54_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10677_ _10561_/A _10558_/Y _10560_/B vssd1 vssd1 vccd1 vccd1 _10679_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__10280__A1 _10136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12416_ hold297/A _12449_/B1 _12414_/X _12415_/Y _12416_/C1 vssd1 vssd1 vccd1 vccd1
+ _12416_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_70_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13396_ _13396_/CLK hold129/X vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10032__A1 _12416_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10583__A2 _07362_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12347_ _12346_/A _12346_/B _12346_/C vssd1 vssd1 vccd1 vccd1 _12348_/B sky130_fd_sc_hd__o21a_1
XANTENNA__07984__B1 _08664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12278_ _12365_/A _12257_/Y _12258_/X _12277_/X vssd1 vssd1 vccd1 vccd1 _12278_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11229_ _11229_/A _11434_/A vssd1 vssd1 vccd1 vccd1 _11229_/X sky130_fd_sc_hd__and2_1
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08528__A2 _10221_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11532__A1 max_cap3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10335__A2 _08877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06770_ _06768_/Y _06770_/B vssd1 vssd1 vccd1 vccd1 _10423_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__09489__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11296__B1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12189__S _12404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08440_ _08540_/B _08576_/A2 _09472_/A _08515_/A2 vssd1 vssd1 vccd1 vccd1 _08441_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_86_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08371_ _09670_/A _08371_/B vssd1 vssd1 vccd1 vccd1 _08375_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_18_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09661__B1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07322_ _07323_/A _07323_/B vssd1 vssd1 vccd1 vccd1 _07601_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_116_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07253_ _10749_/A _07254_/B vssd1 vssd1 vccd1 vccd1 _07255_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_73_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12218__A _12218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07184_ reg1_val[17] _07184_/B vssd1 vssd1 vccd1 vccd1 _10209_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__10023__A1 _10297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11771__A1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11771__B2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09825_ _11497_/A _09825_/B vssd1 vssd1 vccd1 vccd1 _09827_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_39_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06968_ _12438_/A _07147_/B vssd1 vssd1 vccd1 vccd1 _07314_/B sky130_fd_sc_hd__and2_2
X_09756_ _09225_/Y _09745_/Y _09746_/Y _09755_/Y vssd1 vssd1 vccd1 vccd1 _09756_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_69_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09687_ _09688_/A _09688_/B vssd1 vssd1 vccd1 vccd1 _09687_/Y sky130_fd_sc_hd__nor2_1
X_08707_ _08708_/A _08708_/B vssd1 vssd1 vccd1 vccd1 _08707_/X sky130_fd_sc_hd__xor2_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06899_ _08663_/A _06894_/Y _10423_/A _06809_/Y _09418_/A vssd1 vssd1 vccd1 vccd1
+ _06900_/C sky130_fd_sc_hd__o2111a_1
X_08638_ _08638_/A _08638_/B _08646_/A vssd1 vssd1 vccd1 vccd1 _08674_/A sky130_fd_sc_hd__and3_1
XFILLER_0_84_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11039__A0 _12420_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout20 _11497_/A vssd1 vssd1 vccd1 vccd1 _12017_/A sky130_fd_sc_hd__buf_4
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout31 fanout32/X vssd1 vssd1 vccd1 vccd1 _07959_/B sky130_fd_sc_hd__clkbuf_8
X_08569_ _08569_/A _08569_/B vssd1 vssd1 vccd1 vccd1 _08585_/A sky130_fd_sc_hd__xnor2_2
X_11580_ _11929_/A _11580_/B vssd1 vssd1 vccd1 vccd1 _11582_/B sky130_fd_sc_hd__xor2_1
Xfanout64 _07014_/Y vssd1 vssd1 vccd1 vccd1 _11868_/A sky130_fd_sc_hd__buf_4
X_10600_ _10600_/A _10600_/B vssd1 vssd1 vccd1 vccd1 _10611_/A sky130_fd_sc_hd__xnor2_2
Xfanout42 _07159_/X vssd1 vssd1 vccd1 vccd1 fanout42/X sky130_fd_sc_hd__buf_6
Xfanout53 _07072_/Y vssd1 vssd1 vccd1 vccd1 fanout53/X sky130_fd_sc_hd__buf_6
XFILLER_0_49_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08455__B2 _08649_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08455__A1 _08657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout75 _07271_/X vssd1 vssd1 vccd1 vccd1 fanout75/X sky130_fd_sc_hd__buf_8
X_10531_ _10532_/B _10532_/A vssd1 vssd1 vccd1 vccd1 _10531_/Y sky130_fd_sc_hd__nand2b_1
Xfanout86 _08411_/B vssd1 vssd1 vccd1 vccd1 fanout86/X sky130_fd_sc_hd__buf_8
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout97 _07116_/X vssd1 vssd1 vccd1 vccd1 _09834_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_52_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13250_ hold140/X _13250_/B vssd1 vssd1 vccd1 vccd1 hold141/A sky130_fd_sc_hd__nand2_1
XFILLER_0_45_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13200__B2 _13223_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12201_ hold284/A _12449_/B1 _12270_/B _12376_/C1 vssd1 vssd1 vccd1 vccd1 _12202_/B
+ sky130_fd_sc_hd__a31o_1
X_10462_ fanout65/X fanout36/X fanout34/X _12009_/A vssd1 vssd1 vccd1 vccd1 _10463_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13181_ hold292/X _13223_/A2 _13180_/X _13223_/B2 vssd1 vssd1 vccd1 vccd1 _13182_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10871__A _10871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10393_ _10393_/A _10393_/B vssd1 vssd1 vccd1 vccd1 _10395_/C sky130_fd_sc_hd__xor2_1
XANTENNA__12562__S _12638_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12132_ reg1_val[25] curr_PC[25] vssd1 vssd1 vccd1 vccd1 _12133_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08341__A _08575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12063_ _12063_/A _12063_/B vssd1 vssd1 vccd1 vccd1 _12063_/Y sky130_fd_sc_hd__xnor2_1
X_11014_ _11227_/A _11014_/B vssd1 vssd1 vccd1 vccd1 _11050_/D sky130_fd_sc_hd__xor2_4
XANTENNA__07718__B1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11906__S _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08930__A2 _07417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12965_ hold282/X hold58/X vssd1 vssd1 vccd1 vccd1 _12966_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_35_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11916_ _09152_/Y _10563_/X _10575_/X _09221_/Y _11915_/Y vssd1 vssd1 vccd1 vccd1
+ _11916_/X sky130_fd_sc_hd__a221o_1
X_12896_ hold279/X hold85/X vssd1 vssd1 vccd1 vccd1 _13153_/A sky130_fd_sc_hd__nand2b_1
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ _11848_/A _11848_/B vssd1 vssd1 vccd1 vccd1 _11939_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_68_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ _11778_/A _11778_/B vssd1 vssd1 vccd1 vccd1 _11781_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10729_ _12233_/B fanout36/X fanout34/X _12233_/A vssd1 vssd1 vccd1 vccd1 _10730_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_43_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08516__A _08564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13379_ _13379_/CLK _13379_/D vssd1 vssd1 vccd1 vccd1 hold264/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_7_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13390_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_62_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07957__B1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07940_ _07938_/A _07938_/B _08015_/A vssd1 vssd1 vccd1 vccd1 _07953_/A sky130_fd_sc_hd__a21bo_2
XANTENNA__10308__A2 _12420_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07871_ _07868_/A _07868_/B _07952_/A vssd1 vssd1 vccd1 vccd1 _07880_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_92_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12501__A _12670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06822_ _06809_/Y _06820_/X _06821_/X vssd1 vssd1 vccd1 vccd1 _06822_/X sky130_fd_sc_hd__a21o_1
X_09610_ _09936_/A _09610_/B vssd1 vssd1 vccd1 vccd1 _09614_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08921__A2 _08799_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06753_ _10808_/S _06754_/B vssd1 vssd1 vccd1 vccd1 _06753_/Y sky130_fd_sc_hd__nor2_1
X_09541_ _09542_/B _09542_/A vssd1 vssd1 vccd1 vccd1 _09541_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__11808__A2 _11807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08134__B1 _08501_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06684_ _07014_/A reg1_val[22] vssd1 vssd1 vccd1 vccd1 _11913_/S sky130_fd_sc_hd__and2b_1
XFILLER_0_92_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09472_ _09472_/A _11497_/A vssd1 vssd1 vccd1 vccd1 _09478_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_25_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07488__A2 _07554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10492__B2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06696__B1 _06766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10492__A1 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08423_ _08423_/A _08423_/B vssd1 vssd1 vccd1 vccd1 _08468_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_25_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08354_ _08351_/A _08351_/B _08353_/X vssd1 vssd1 vccd1 vccd1 _08365_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_128_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07305_ _10623_/A _07305_/B vssd1 vssd1 vccd1 vccd1 _07413_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06999__B2 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06999__A1 _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08285_ _08323_/A _08323_/B vssd1 vssd1 vccd1 vccd1 _08285_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_27_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07236_ _07215_/A _07133_/A _06974_/B _07215_/B vssd1 vssd1 vccd1 vccd1 _07238_/B
+ sky130_fd_sc_hd__o31a_4
X_07167_ reg1_val[24] _07167_/B vssd1 vssd1 vccd1 vccd1 _07168_/C sky130_fd_sc_hd__xor2_2
XFILLER_0_42_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11744__A1 _07016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08799__C _08799_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07098_ _07092_/B _10350_/A _10479_/A vssd1 vssd1 vccd1 vccd1 _07098_/X sky130_fd_sc_hd__mux2_2
Xfanout232 _12271_/A1 vssd1 vssd1 vccd1 vccd1 _11650_/B sky130_fd_sc_hd__buf_4
Xfanout210 _06946_/X vssd1 vssd1 vccd1 vccd1 _12446_/C1 sky130_fd_sc_hd__clkbuf_8
Xfanout221 _06805_/X vssd1 vssd1 vccd1 vccd1 _07172_/A sky130_fd_sc_hd__buf_4
Xfanout254 _06577_/Y vssd1 vssd1 vccd1 vccd1 _12805_/A sky130_fd_sc_hd__buf_4
Xfanout243 _12520_/S vssd1 vssd1 vccd1 vccd1 _12471_/S sky130_fd_sc_hd__clkbuf_4
Xfanout265 _12796_/A vssd1 vssd1 vccd1 vccd1 _12755_/B sky130_fd_sc_hd__buf_12
XANTENNA__07176__A1 _07166_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout276 _13162_/A vssd1 vssd1 vccd1 vccd1 _13249_/A sky130_fd_sc_hd__buf_4
X_09808_ fanout53/X _08199_/B fanout34/X fanout51/X vssd1 vssd1 vccd1 vccd1 _09809_/B
+ sky130_fd_sc_hd__o22a_1
Xfanout287 _06581_/Y vssd1 vssd1 vccd1 vccd1 _06992_/A sky130_fd_sc_hd__buf_6
XANTENNA__08373__B1 _08501_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07176__B2 _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout62_A _07019_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09739_ _10295_/S _09198_/X _09248_/B vssd1 vssd1 vccd1 vccd1 _09739_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_69_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09873__B1 _10788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12750_ reg1_val[22] _12755_/B vssd1 vssd1 vccd1 vccd1 _12751_/B sky130_fd_sc_hd__or2_1
X_11701_ _11701_/A _11701_/B vssd1 vssd1 vccd1 vccd1 _11703_/B sky130_fd_sc_hd__xnor2_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _12679_/Y _12681_/B vssd1 vssd1 vccd1 vccd1 _12682_/B sky130_fd_sc_hd__nand2b_2
X_11632_ _11813_/S _11632_/B vssd1 vssd1 vccd1 vccd1 _11636_/B sky130_fd_sc_hd__or2_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09625__B1 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07240__A _09341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13302_ _13304_/CLK _13302_/D vssd1 vssd1 vccd1 vccd1 hold196/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10786__A2 _11050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11563_ _10788_/A _11537_/Y _11538_/X _11562_/Y _11536_/Y vssd1 vssd1 vccd1 vccd1
+ _11563_/X sky130_fd_sc_hd__o311a_1
XFILLER_0_24_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11494_ _11868_/A fanout23/X fanout15/X fanout62/X vssd1 vssd1 vccd1 vccd1 _11495_/B
+ sky130_fd_sc_hd__o22a_1
X_10514_ _10514_/A _10514_/B vssd1 vssd1 vccd1 vccd1 _10515_/B sky130_fd_sc_hd__xor2_1
X_13233_ _13246_/A hold283/X vssd1 vssd1 vccd1 vccd1 _13388_/D sky130_fd_sc_hd__and2_1
XFILLER_0_107_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10445_ _09222_/Y _10432_/Y _10444_/Y _10159_/A _10443_/X vssd1 vssd1 vccd1 vccd1
+ _10445_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_122_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13164_ _13164_/A _13164_/B vssd1 vssd1 vccd1 vccd1 _13164_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12115_ _12115_/A vssd1 vssd1 vccd1 vccd1 _12115_/Y sky130_fd_sc_hd__inv_2
X_10376_ _10376_/A _10376_/B _10376_/C vssd1 vssd1 vccd1 vccd1 _10377_/B sky130_fd_sc_hd__and3_1
X_13095_ _07361_/B _13101_/B2 hold144/X vssd1 vssd1 vccd1 vccd1 _13357_/D sky130_fd_sc_hd__o21a_1
X_12046_ _11715_/X _12043_/A _12043_/B _12302_/A vssd1 vssd1 vccd1 vccd1 _12046_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_99_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12948_ _12886_/X _12948_/B vssd1 vssd1 vccd1 vccd1 _13198_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12879_ hold276/X hold44/X vssd1 vssd1 vccd1 vccd1 _12880_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_87_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10226__A1 _10225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12991__A _13001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08070_ _08070_/A _08070_/B vssd1 vssd1 vccd1 vccd1 _08170_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07021_ _09669_/B2 fanout63/X _09301_/A fanout61/X vssd1 vssd1 vccd1 vccd1 _07022_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09077__A _10479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10661__D _10779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08972_ _09673_/A _08972_/B vssd1 vssd1 vccd1 vccd1 _08982_/A sky130_fd_sc_hd__xnor2_4
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09805__A _11179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
X_07923_ _08454_/A _07923_/B vssd1 vssd1 vccd1 vccd1 _07924_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout197_A _09228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07854_ _07850_/A _07850_/B _07888_/A vssd1 vssd1 vccd1 vccd1 _07861_/B sky130_fd_sc_hd__o21ba_1
X_06805_ _06815_/A _06817_/B1 _12655_/B _06803_/X vssd1 vssd1 vccd1 vccd1 _06805_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_127_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07785_ _08457_/A2 fanout86/X fanout82/X _08501_/B1 vssd1 vssd1 vccd1 vccd1 _07786_/B
+ sky130_fd_sc_hd__o22a_1
X_06736_ _11134_/A _07270_/A vssd1 vssd1 vccd1 vccd1 _06738_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_78_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12454__A2 _11829_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09524_ _09525_/A _09525_/B vssd1 vssd1 vccd1 vccd1 _09694_/A sky130_fd_sc_hd__nor2_1
X_06667_ reg2_val[26] _06766_/B _06677_/B1 _06666_/Y vssd1 vssd1 vccd1 vccd1 _07046_/B
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_66_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09455_ _07417_/B _10337_/A _12823_/A1 fanout42/X vssd1 vssd1 vccd1 vccd1 _09456_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08406_ _08406_/A _08406_/B vssd1 vssd1 vccd1 vccd1 _08407_/B sky130_fd_sc_hd__xor2_2
X_06598_ instruction[11] _06590_/X _06597_/X _06716_/B vssd1 vssd1 vccd1 vccd1 reg1_idx[0]
+ sky130_fd_sc_hd__o211a_4
XFILLER_0_74_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09386_ _09170_/X _09172_/X _09403_/S vssd1 vssd1 vccd1 vccd1 _09386_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08337_ _08627_/A2 _10221_/B2 _08501_/B1 _08641_/B vssd1 vssd1 vccd1 vccd1 _08338_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_62_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08268_ _08268_/A _08268_/B vssd1 vssd1 vccd1 vccd1 _08327_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_22_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07219_ _06827_/B _06793_/Y _06970_/X _06969_/Y vssd1 vssd1 vccd1 vccd1 _07283_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_6_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10230_ _07171_/A _07262_/X _07269_/Y fanout38/X vssd1 vssd1 vccd1 vccd1 _10231_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08199_ _09404_/S _08199_/B vssd1 vssd1 vccd1 vccd1 _08265_/B sky130_fd_sc_hd__nor2_1
X_10161_ _09567_/X _09572_/X _10295_/S vssd1 vssd1 vccd1 vccd1 _10161_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10940__A2 _07171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10092_ _10092_/A _10092_/B vssd1 vssd1 vccd1 vccd1 _10096_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10994_ _10995_/B _10995_/A vssd1 vssd1 vccd1 vccd1 _11108_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_97_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12802_ _12805_/A hold68/X vssd1 vssd1 vccd1 vccd1 _12803_/C sky130_fd_sc_hd__nor2_1
XANTENNA__08649__A1 _09404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08649__B2 _08657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10456__B2 _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10456__A1 _12233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ _12755_/B _07109_/C _12739_/A _12739_/B vssd1 vssd1 vccd1 vccd1 _12734_/B
+ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__09310__A2 fanout86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10596__A _12087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10208__A1 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12664_ reg1_val[5] _12665_/B vssd1 vssd1 vccd1 vccd1 _12664_/Y sky130_fd_sc_hd__nor2_1
X_12595_ _12633_/A _12595_/B vssd1 vssd1 vccd1 vccd1 _12596_/B sky130_fd_sc_hd__or2_1
X_11615_ _11617_/A vssd1 vssd1 vccd1 vccd1 _11615_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10208__B2 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11546_ _11454_/A _11451_/Y _11453_/B vssd1 vssd1 vccd1 vccd1 _11547_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11477_ _11477_/A _11600_/A vssd1 vssd1 vccd1 vccd1 _11479_/C sky130_fd_sc_hd__nor2_1
X_13216_ _13216_/A _13216_/B vssd1 vssd1 vccd1 vccd1 _13216_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__11184__A2 _07171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10428_ _10426_/Y _10428_/B vssd1 vssd1 vccd1 vccd1 _10429_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10359_ fanout43/X _07269_/Y _07274_/Y fanout41/X vssd1 vssd1 vccd1 vccd1 _10360_/B
+ sky130_fd_sc_hd__a22o_1
X_13147_ _13147_/A _13147_/B vssd1 vssd1 vccd1 vccd1 _13370_/D sky130_fd_sc_hd__and2_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13078_ hold113/A _12805_/A _13250_/B hold103/X _13259_/A vssd1 vssd1 vccd1 vccd1
+ hold104/A sky130_fd_sc_hd__o221a_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12029_ _12030_/A _12030_/B _12030_/C vssd1 vssd1 vccd1 vccd1 _12108_/B sky130_fd_sc_hd__a21o_1
XANTENNA__13147__A _13147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06968__B _07147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08337__B1 _08501_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06984__A _07016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07570_ _07568_/A _07568_/B _07569_/Y vssd1 vssd1 vccd1 vccd1 _07677_/A sky130_fd_sc_hd__a21bo_2
XFILLER_0_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10447__A1 _10788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09240_ hold293/A _09236_/Y _09238_/Y hold245/A _09235_/X vssd1 vssd1 vccd1 vccd1
+ _09241_/B sky130_fd_sc_hd__a221o_1
XFILLER_0_118_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09171_ _09169_/X _09170_/X _09383_/S vssd1 vssd1 vccd1 vccd1 _09171_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11947__A1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08122_ _08122_/A _08122_/B vssd1 vssd1 vccd1 vccd1 _08131_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_126_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08053_ _09341_/A _08053_/B vssd1 vssd1 vccd1 vccd1 _08054_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout112_A _07233_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07004_ reg1_val[5] _07004_/B vssd1 vssd1 vccd1 vccd1 _07004_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_113_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08576__B1 _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08955_ fanout57/X _10245_/B2 _10245_/A1 fanout63/X vssd1 vssd1 vccd1 vccd1 _08956_/B
+ sky130_fd_sc_hd__o22a_1
X_07906_ _07968_/A _07968_/B vssd1 vssd1 vccd1 vccd1 _07969_/A sky130_fd_sc_hd__nor2_1
X_08886_ _09341_/A _08886_/B vssd1 vssd1 vccd1 vccd1 _08890_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10686__A1 _11990_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07837_ _07837_/A _07837_/B _07837_/C vssd1 vssd1 vccd1 vccd1 _07842_/A sky130_fd_sc_hd__or3_1
XANTENNA__07055__A _09947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07768_ _12808_/A fanout46/X _09325_/A _07830_/B vssd1 vssd1 vccd1 vccd1 _07769_/B
+ sky130_fd_sc_hd__o22a_1
X_06719_ _07097_/A reg1_val[17] vssd1 vssd1 vccd1 vccd1 _06719_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_78_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06894__A _09218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09507_ _09507_/A _09507_/B vssd1 vssd1 vccd1 vccd1 _09508_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_78_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07699_ fanout61/X _09298_/B2 _09298_/A1 fanout53/X vssd1 vssd1 vccd1 vccd1 _07700_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_94_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _10165_/S _09437_/Y _09251_/A vssd1 vssd1 vccd1 vccd1 _12412_/B sky130_fd_sc_hd__o21ai_2
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout25_A _07235_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06655__A2_N _06783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09369_ _09369_/A _09369_/B vssd1 vssd1 vccd1 vccd1 _09371_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11400_ _11401_/A _11401_/B vssd1 vssd1 vccd1 vccd1 _11410_/A sky130_fd_sc_hd__nand2_1
X_12380_ _12380_/A _12380_/B _12376_/X vssd1 vssd1 vccd1 vccd1 _12381_/C sky130_fd_sc_hd__or3b_1
X_11331_ _11331_/A _11331_/B _11331_/C vssd1 vssd1 vccd1 vccd1 _11332_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_62_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11262_ _11247_/A _09215_/X _09251_/A vssd1 vssd1 vccd1 vccd1 _11262_/X sky130_fd_sc_hd__o21a_1
XANTENNA__11166__A2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11193_ _11193_/A _11193_/B vssd1 vssd1 vccd1 vccd1 _11194_/B sky130_fd_sc_hd__xor2_2
X_13001_ _13001_/A hold170/X vssd1 vssd1 vccd1 vccd1 hold171/A sky130_fd_sc_hd__and2_1
X_10213_ fanout65/X fanout78/X fanout74/X fanout59/X vssd1 vssd1 vccd1 vccd1 _10214_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12363__A1 _10049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10144_ _10138_/X _10139_/X _10143_/Y _10661_/A vssd1 vssd1 vccd1 vccd1 _10146_/A
+ sky130_fd_sc_hd__a31o_1
X_10075_ _10075_/A _10075_/B vssd1 vssd1 vccd1 vccd1 _10076_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_69_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10977_ _10976_/A _10976_/B _10976_/C vssd1 vssd1 vccd1 vccd1 _10984_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__13091__A2 _13101_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12823__C1 _13147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08508__B _08508_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12716_ _12717_/A _12717_/B _12717_/C vssd1 vssd1 vccd1 vccd1 _12721_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_128_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12647_ _12647_/A _12647_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[1] sky130_fd_sc_hd__xor2_4
XFILLER_0_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09598__A2 _12144_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10601__A1 _11671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12578_ reg1_val[18] curr_PC[18] _12638_/S vssd1 vssd1 vccd1 vccd1 _12580_/B sky130_fd_sc_hd__mux2_1
XANTENNA__06970__C _09728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06805__B1 _06803_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10601__B2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11529_ _11330_/Y _11430_/Y _11432_/B vssd1 vssd1 vccd1 vccd1 _11529_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_80_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold307 hold307/A vssd1 vssd1 vccd1 vccd1 hold307/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09770__A2 _07362_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08740_ _08733_/A _08733_/B _08733_/C _08739_/Y vssd1 vssd1 vccd1 vccd1 _08741_/C
+ sky130_fd_sc_hd__a31o_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08671_ _08671_/A _08671_/B vssd1 vssd1 vccd1 vccd1 _08721_/B sky130_fd_sc_hd__nor2_1
X_07622_ _10479_/A _07622_/B vssd1 vssd1 vccd1 vccd1 _07624_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_88_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08089__A2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07553_ _09834_/A _07553_/B vssd1 vssd1 vccd1 vccd1 _07706_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07484_ _07830_/B _09677_/A _07172_/Y fanout46/X vssd1 vssd1 vccd1 vccd1 _07485_/B
+ sky130_fd_sc_hd__o22a_1
X_09223_ _09237_/B _09228_/B vssd1 vssd1 vccd1 vccd1 _11554_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_118_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09154_ _12644_/A reg1_val[30] _09180_/S vssd1 vssd1 vccd1 vccd1 _09154_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11779__B _12428_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10053__C1 _11946_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08105_ _08108_/A _08108_/B vssd1 vssd1 vccd1 vccd1 _08110_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_114_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09085_ _09085_/A _09085_/B vssd1 vssd1 vccd1 vccd1 _09089_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_102_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06811__A3 _12650_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08036_ _08036_/A _08036_/B vssd1 vssd1 vccd1 vccd1 _08081_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09987_ _09784_/A _09784_/B _09783_/A vssd1 vssd1 vccd1 vccd1 _09992_/A sky130_fd_sc_hd__a21o_2
X_08938_ _08834_/A _08834_/B _08832_/Y vssd1 vssd1 vccd1 vccd1 _08939_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_99_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09513__A2 _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08869_ _08869_/A _08869_/B vssd1 vssd1 vccd1 vccd1 _08882_/A sky130_fd_sc_hd__xnor2_1
X_10900_ _10900_/A _11008_/A vssd1 vssd1 vccd1 vccd1 _11122_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07524__A1 _09943_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07524__B2 _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11880_ _11881_/A _11881_/B _11881_/C vssd1 vssd1 vccd1 vccd1 _11883_/A sky130_fd_sc_hd__a21o_1
X_10831_ _07255_/A fanout7/X _10950_/A vssd1 vssd1 vccd1 vccd1 _10831_/Y sky130_fd_sc_hd__o21ai_1
X_10762_ _10612_/A _10612_/B _10610_/Y vssd1 vssd1 vccd1 vccd1 _10765_/A sky130_fd_sc_hd__o21a_1
XANTENNA__12281__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07288__B1 _10500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12501_ _12670_/B _12501_/B vssd1 vssd1 vccd1 vccd1 _12502_/B sky130_fd_sc_hd__or2_1
X_12432_ _12351_/X _12430_/C _12430_/X _12249_/B _12431_/Y vssd1 vssd1 vccd1 vccd1
+ _12433_/B sky130_fd_sc_hd__o221a_1
X_10693_ _07233_/A _12422_/A _10689_/Y vssd1 vssd1 vccd1 vccd1 _10693_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10595__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12363_ _10049_/A _08810_/Y _12364_/B vssd1 vssd1 vccd1 vccd1 _12365_/B sky130_fd_sc_hd__a21bo_1
X_11314_ _11196_/A _11196_/B _11203_/Y vssd1 vssd1 vccd1 vccd1 _11324_/A sky130_fd_sc_hd__o21ai_2
X_12294_ _12346_/B _12294_/B vssd1 vssd1 vccd1 vccd1 _12296_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_22_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11245_ _11245_/A _11245_/B vssd1 vssd1 vccd1 vccd1 _11245_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10347__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11176_ fanout26/X fanout17/X fanout14/X fanout28/X vssd1 vssd1 vccd1 vccd1 _11177_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10127_ _10127_/A _10127_/B vssd1 vssd1 vccd1 vccd1 _10128_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__08960__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10058_ _10950_/A _10058_/B vssd1 vssd1 vccd1 vccd1 _10066_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06965__C _12359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07423__A _09922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12811__A2 _13101_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10784__A _11008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11378__A2 _07316_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08254__A _08580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08243__A2 _10338_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold104 hold104/A vssd1 vssd1 vccd1 vccd1 hold104/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 hold115/A vssd1 vssd1 vccd1 vccd1 hold115/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 hold126/A vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold137 hold137/A vssd1 vssd1 vccd1 vccd1 hold137/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 hold159/A vssd1 vssd1 vccd1 vccd1 hold159/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 hold148/A vssd1 vssd1 vccd1 vccd1 hold148/X sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ _10049_/A _09910_/B vssd1 vssd1 vccd1 vccd1 _09910_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10338__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09841_ _09960_/A _09841_/B _09842_/B vssd1 vssd1 vccd1 vccd1 _09841_/X sky130_fd_sc_hd__and3_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07203__B1 _10725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06984_ _07016_/A _06984_/B vssd1 vssd1 vccd1 vccd1 _06986_/C sky130_fd_sc_hd__and2_2
XANTENNA__10024__A _11138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09772_ _07554_/B _10234_/A2 _10725_/A _07175_/A vssd1 vssd1 vccd1 vccd1 _09773_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09427__A2_N _11554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07317__B _10476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08951__B1 _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09813__A _09944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08723_ _08723_/A _08723_/B vssd1 vssd1 vccd1 vccd1 _10151_/C sky130_fd_sc_hd__xor2_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout277_A _13001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08654_ _08654_/A _08654_/B vssd1 vssd1 vccd1 vccd1 _08719_/A sky130_fd_sc_hd__xnor2_2
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07605_ _06867_/B _07315_/A _07094_/B _08973_/A vssd1 vssd1 vccd1 vccd1 _07608_/A
+ sky130_fd_sc_hd__a211o_4
XANTENNA__13055__A2 _12820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09259__A1 _11752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08585_ _08585_/A _08585_/B vssd1 vssd1 vccd1 vccd1 _08605_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_119_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12263__B1 _12064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07536_ _07533_/A _07533_/C _07533_/B vssd1 vssd1 vccd1 vccd1 _07537_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_119_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09206_ _09202_/X _09205_/X _09727_/S vssd1 vssd1 vccd1 vccd1 _09206_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07467_ _07466_/A _07466_/B _07495_/A vssd1 vssd1 vccd1 vccd1 _07467_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_29_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07398_ _07434_/A _07434_/B vssd1 vssd1 vccd1 vccd1 _07435_/A sky130_fd_sc_hd__and2_1
XFILLER_0_8_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09137_ _09137_/A _09137_/B vssd1 vssd1 vccd1 vccd1 _09139_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10041__A2 _10026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09068_ _09069_/A _09069_/B vssd1 vssd1 vccd1 vccd1 _09278_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_114_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08019_ _08580_/A _08019_/B vssd1 vssd1 vccd1 vccd1 _08094_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout92_A _09779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09195__A0 _12644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09707__B _09707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11030_ _12412_/A _11030_/B vssd1 vssd1 vccd1 vccd1 _11030_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_99_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12981_ _13001_/A hold222/X vssd1 vssd1 vccd1 vccd1 hold223/A sky130_fd_sc_hd__and2_1
X_11932_ _11933_/B _11932_/B vssd1 vssd1 vccd1 vccd1 _12012_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_99_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08339__A _08342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11863_ _11770_/A _11770_/B _11775_/A vssd1 vssd1 vccd1 vccd1 _11867_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__13046__A2 _06577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10814_ _10811_/Y _10812_/X _10813_/Y _10809_/X vssd1 vssd1 vccd1 vccd1 _10814_/X
+ sky130_fd_sc_hd__o211a_1
X_11794_ _11881_/B _11794_/B vssd1 vssd1 vccd1 vccd1 _11797_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_94_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10804__A1 _12064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10745_ _10950_/A _10745_/B vssd1 vssd1 vccd1 vccd1 _10751_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12006__B1 _12093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10676_ reg1_val[10] curr_PC[10] vssd1 vssd1 vccd1 vccd1 _10679_/B sky130_fd_sc_hd__or2_1
XFILLER_0_70_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10280__A2 _10136_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12415_ _12449_/B1 _12414_/X hold297/A vssd1 vssd1 vccd1 vccd1 _12415_/Y sky130_fd_sc_hd__a21oi_1
X_13395_ _13396_/CLK hold307/X vssd1 vssd1 vccd1 vccd1 hold200/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12346_ _12346_/A _12346_/B _12346_/C vssd1 vssd1 vccd1 vccd1 _12348_/A sky130_fd_sc_hd__nor3_1
XANTENNA__10568__B1 _11554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12277_ _12277_/A _12277_/B _12277_/C _12272_/X vssd1 vssd1 vccd1 vccd1 _12277_/X
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_10_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11228_ _11010_/Y _11434_/A _11226_/X vssd1 vssd1 vccd1 vccd1 _11623_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07418__A _09779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11159_ curr_PC[13] curr_PC[14] _11159_/C vssd1 vssd1 vccd1 vccd1 _11268_/B sky130_fd_sc_hd__and3_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10779__A _10779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06976__B _07233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09489__A1 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09489__B2 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11296__B2 _11946_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11296__A1 _07032_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08370_ _08641_/B _10221_/B2 _09770_/B2 _08627_/A2 vssd1 vssd1 vccd1 vccd1 _08371_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_58_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06992__A _06992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07321_ _09947_/A _07321_/B vssd1 vssd1 vccd1 vccd1 _07323_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_105_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09661__A1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09661__B2 _09661_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11403__A _12017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07252_ reg1_val[12] _07252_/B vssd1 vssd1 vccd1 vccd1 _07254_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07183_ reg1_val[17] _07184_/B vssd1 vssd1 vccd1 vccd1 _07183_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_5_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11771__A2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12234__A _12335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09824_ _07283_/X _08877_/B fanout6/X _09934_/A vssd1 vssd1 vccd1 vccd1 _09825_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_10_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10731__B1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09755_ _09748_/Y _09749_/X _09754_/X vssd1 vssd1 vccd1 vccd1 _09755_/Y sky130_fd_sc_hd__o21ai_1
X_06967_ _12644_/A _06967_/B vssd1 vssd1 vccd1 vccd1 _08502_/A sky130_fd_sc_hd__xnor2_4
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06898_ _10155_/A _06898_/B _06898_/C _09745_/B vssd1 vssd1 vccd1 vccd1 _06901_/C
+ sky130_fd_sc_hd__and4b_1
X_09686_ _09686_/A _09686_/B vssd1 vssd1 vccd1 vccd1 _09688_/B sky130_fd_sc_hd__xnor2_1
X_08706_ _08706_/A _08706_/B vssd1 vssd1 vccd1 vccd1 _08805_/B sky130_fd_sc_hd__xnor2_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ _08637_/A _08637_/B _08637_/C vssd1 vssd1 vccd1 vccd1 _08646_/A sky130_fd_sc_hd__or3_2
XANTENNA__13028__A2 _13223_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11039__A1 _09422_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout10 _08877_/B vssd1 vssd1 vccd1 vccd1 fanout10/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout21 _12009_/B vssd1 vssd1 vccd1 vccd1 _11497_/A sky130_fd_sc_hd__buf_12
X_08568_ _08568_/A _08568_/B _08568_/C vssd1 vssd1 vccd1 vccd1 _08681_/B sky130_fd_sc_hd__nand3_2
Xfanout54 _07072_/Y vssd1 vssd1 vccd1 vccd1 _11671_/A sky130_fd_sc_hd__buf_4
XFILLER_0_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout65 _06997_/Y vssd1 vssd1 vccd1 vccd1 fanout65/X sky130_fd_sc_hd__buf_6
XFILLER_0_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout43 _07417_/B vssd1 vssd1 vccd1 vccd1 fanout43/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout32 _07213_/Y vssd1 vssd1 vccd1 vccd1 fanout32/X sky130_fd_sc_hd__clkbuf_8
X_08499_ _08500_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08521_/B sky130_fd_sc_hd__or2_1
X_07519_ _09669_/B2 fanout53/X fanout51/X _09301_/A vssd1 vssd1 vccd1 vccd1 _07520_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08455__A2 _10221_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout87 _07255_/Y vssd1 vssd1 vccd1 vccd1 _08411_/B sky130_fd_sc_hd__buf_8
X_10530_ _10530_/A _10530_/B vssd1 vssd1 vccd1 vccd1 _10532_/B sky130_fd_sc_hd__xnor2_1
Xfanout98 _07096_/Y vssd1 vssd1 vccd1 vccd1 fanout98/X sky130_fd_sc_hd__buf_6
Xfanout76 _11093_/A vssd1 vssd1 vccd1 vccd1 fanout76/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10461_ _10461_/A _10461_/B vssd1 vssd1 vccd1 vccd1 _10465_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_52_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13200__A2 _13223_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12200_ _12449_/B1 _12270_/B hold284/A vssd1 vssd1 vccd1 vccd1 _12202_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13180_ hold275/X _13179_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13180_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10871__B _12087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10392_ _11284_/A _10392_/B vssd1 vssd1 vccd1 vccd1 _10393_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07415__B1 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12131_ reg1_val[25] curr_PC[25] vssd1 vssd1 vccd1 vccd1 _12131_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_60_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12062_ _12060_/Y _12062_/B vssd1 vssd1 vccd1 vccd1 _12063_/B sky130_fd_sc_hd__and2b_1
X_11013_ _10006_/B _10542_/X _11009_/Y _11012_/Y vssd1 vssd1 vccd1 vccd1 _11014_/B
+ sky130_fd_sc_hd__o31a_2
XANTENNA__07718__B2 _10221_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07718__A1 _08501_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10599__A _10599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12964_ _13229_/A _13230_/A _13229_/B vssd1 vssd1 vccd1 vccd1 _13234_/A sky130_fd_sc_hd__a21bo_1
X_11915_ _07014_/A _09257_/S _11914_/X vssd1 vssd1 vccd1 vccd1 _11915_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09340__B1 _11093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12895_ hold288/A hold94/X vssd1 vssd1 vccd1 vccd1 _13158_/A sky130_fd_sc_hd__nand2b_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _12096_/A _11846_/B vssd1 vssd1 vccd1 vccd1 _11848_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _11687_/A _11687_/B _11675_/A vssd1 vssd1 vccd1 vccd1 _11788_/A sky130_fd_sc_hd__o21a_1
XANTENNA__12319__A _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10728_ _10728_/A _10728_/B vssd1 vssd1 vccd1 vccd1 _10739_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10659_ _10661_/C _10779_/A vssd1 vssd1 vccd1 vccd1 _10902_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13378_ _13379_/CLK _13378_/D vssd1 vssd1 vccd1 vccd1 hold246/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09628__A _09834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07406__B1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07957__A1 _08561_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12329_ _12379_/B2 _09732_/B _12319_/B _09221_/Y _12328_/X vssd1 vssd1 vccd1 vccd1
+ _12329_/Y sky130_fd_sc_hd__a221oi_2
XFILLER_0_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07957__B2 _08576_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07148__A _09728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12989__A _13001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10713__B1 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07870_ _07951_/A _07951_/B vssd1 vssd1 vccd1 vccd1 _07952_/A sky130_fd_sc_hd__nor2_1
X_06821_ reg1_val[2] _10297_/S vssd1 vssd1 vccd1 vccd1 _06821_/X sky130_fd_sc_hd__and2_1
X_06752_ reg1_val[11] _10813_/A vssd1 vssd1 vccd1 vccd1 _06754_/B sky130_fd_sc_hd__nor2_1
X_09540_ _09540_/A _09540_/B vssd1 vssd1 vccd1 vccd1 _09542_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_92_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09471_ _09471_/A _09471_/B vssd1 vssd1 vccd1 vccd1 _09511_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08134__A1 _08515_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08134__B2 _08540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06683_ reg2_val[22] _06810_/B _06724_/B1 _06682_/Y vssd1 vssd1 vccd1 vccd1 _07014_/A
+ sky130_fd_sc_hd__o2bb2a_4
X_08422_ _08423_/A _08423_/B vssd1 vssd1 vccd1 vccd1 _08422_/X sky130_fd_sc_hd__or2_1
XFILLER_0_25_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10492__A2 _07262_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07893__B1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08353_ _08405_/A _08405_/B vssd1 vssd1 vccd1 vccd1 _08353_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_18_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11133__A _11134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07304_ fanout86/X fanout80/X fanout76/X fanout82/X vssd1 vssd1 vccd1 vccd1 _07305_/B
+ sky130_fd_sc_hd__o22a_1
X_08284_ _08284_/A _08284_/B vssd1 vssd1 vccd1 vccd1 _08323_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07235_ _11582_/A _11473_/A _07234_/Y vssd1 vssd1 vccd1 vccd1 _07235_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_41_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06999__A2 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07166_ _07166_/A _07166_/B vssd1 vssd1 vccd1 vccd1 _07166_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_42_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11744__A2 _09257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07097_ _07097_/A _07097_/B vssd1 vssd1 vccd1 vccd1 _07097_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_41_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout222 _11028_/S vssd1 vssd1 vccd1 vccd1 _11246_/S sky130_fd_sc_hd__buf_4
Xfanout211 _09383_/S vssd1 vssd1 vccd1 vccd1 _09403_/S sky130_fd_sc_hd__clkbuf_8
Xfanout200 _09149_/Y vssd1 vssd1 vccd1 vccd1 _12356_/B1 sky130_fd_sc_hd__buf_4
Xfanout233 _12271_/A1 vssd1 vssd1 vccd1 vccd1 _12449_/B1 sky130_fd_sc_hd__buf_4
Xfanout255 _12804_/A vssd1 vssd1 vccd1 vccd1 _06577_/A sky130_fd_sc_hd__buf_4
Xfanout244 _06958_/A vssd1 vssd1 vccd1 vccd1 _12520_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__08373__A1 _08657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07176__A2 _07554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout277 _13001_/A vssd1 vssd1 vccd1 vccd1 _13162_/A sky130_fd_sc_hd__buf_2
XANTENNA__10180__A1 _06782_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09807_ _09807_/A _09807_/B vssd1 vssd1 vccd1 vccd1 _09811_/A sky130_fd_sc_hd__xnor2_1
Xfanout266 _12796_/A vssd1 vssd1 vccd1 vccd1 _12790_/B sky130_fd_sc_hd__clkbuf_8
X_07999_ _07889_/A _07889_/B _07889_/C vssd1 vssd1 vccd1 vccd1 _08001_/B sky130_fd_sc_hd__o21ai_1
Xfanout288 _06581_/Y vssd1 vssd1 vccd1 vccd1 _06993_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__08373__B2 _08649_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09273__A _09779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09738_ _09733_/X _09736_/X _09737_/Y vssd1 vssd1 vccd1 vccd1 _09738_/X sky130_fd_sc_hd__a21o_1
XANTENNA_fanout55_A fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09669_ _09301_/A fanout13/X fanout8/X _09669_/B2 vssd1 vssd1 vccd1 vccd1 _09670_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09873__A1 _10049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11700_ _11701_/A _11701_/B vssd1 vssd1 vccd1 vccd1 _11793_/B sky130_fd_sc_hd__and2b_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08617__A _09673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12680_ reg1_val[8] _12680_/B vssd1 vssd1 vccd1 vccd1 _12681_/B sky130_fd_sc_hd__nand2_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09625__A1 _11406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11631_ _11631_/A _11631_/B vssd1 vssd1 vccd1 vccd1 _11631_/Y sky130_fd_sc_hd__nand2_1
X_11562_ _11541_/Y _11542_/X _11561_/Y vssd1 vssd1 vccd1 vccd1 _11562_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09625__B2 _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07636__B1 _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10513_ _11929_/A _10513_/B vssd1 vssd1 vccd1 vccd1 _10514_/B sky130_fd_sc_hd__xnor2_1
X_13301_ _13304_/CLK _13301_/D vssd1 vssd1 vccd1 vccd1 hold300/A sky130_fd_sc_hd__dfxtp_1
X_11493_ _11493_/A _11493_/B vssd1 vssd1 vccd1 vccd1 _11504_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13232_ hold282/X _13248_/B1 _13231_/X _13248_/A2 vssd1 vssd1 vccd1 vccd1 hold283/A
+ sky130_fd_sc_hd__a22o_1
X_10444_ _11247_/A _10298_/X _09251_/A vssd1 vssd1 vccd1 vccd1 _10444_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13163_ _13163_/A _13163_/B vssd1 vssd1 vccd1 vccd1 _13164_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_110_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10375_ _10376_/A _10376_/B _10376_/C vssd1 vssd1 vccd1 vccd1 _10525_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12114_ _12114_/A _12114_/B vssd1 vssd1 vccd1 vccd1 _12115_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13094_ hold116/X _13094_/A2 _13101_/A2 hold56/X _13039_/A vssd1 vssd1 vccd1 vccd1
+ hold144/A sky130_fd_sc_hd__o221a_1
X_12045_ _11887_/Y _12043_/B _12044_/Y vssd1 vssd1 vccd1 vccd1 _12302_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_46_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12947_ hold262/X hold52/X vssd1 vssd1 vccd1 vccd1 _12948_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12878_ hold44/X hold276/X vssd1 vssd1 vccd1 vccd1 _12878_/X sky130_fd_sc_hd__and2b_1
X_11829_ _11829_/A _11829_/B vssd1 vssd1 vccd1 vccd1 _11829_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_56_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12049__A _12049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10226__A2 _11946_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11974__A2 _12049_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13176__B2 _13223_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07020_ _07020_/A _07020_/B vssd1 vssd1 vccd1 vccd1 _11779_/A sky130_fd_sc_hd__nand2_8
XANTENNA__08052__B1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ _09298_/A1 fanout17/X fanout14/X _09298_/B2 vssd1 vssd1 vccd1 vccd1 _08972_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_11_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_07922_ _08457_/A2 _08484_/B _09479_/B1 _08501_/B1 vssd1 vssd1 vccd1 vccd1 _07923_/B
+ sky130_fd_sc_hd__o22a_1
X_07853_ _07887_/B _07853_/B vssd1 vssd1 vccd1 vccd1 _07888_/A sky130_fd_sc_hd__and2b_1
X_06804_ _06815_/A _06817_/B1 _12655_/B _06803_/X vssd1 vssd1 vccd1 vccd1 _10297_/S
+ sky130_fd_sc_hd__a31oi_4
XANTENNA__09304__B1 _09672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07784_ _07784_/A _07784_/B vssd1 vssd1 vccd1 vccd1 _07800_/A sky130_fd_sc_hd__xor2_1
X_06735_ _06815_/A _06723_/A _12719_/B _06734_/X vssd1 vssd1 vccd1 vccd1 _07270_/A
+ sky130_fd_sc_hd__a31o_4
X_09523_ _09325_/A _11497_/A _09331_/B _09329_/X vssd1 vssd1 vccd1 vccd1 _09525_/B
+ sky130_fd_sc_hd__o31a_1
X_06666_ _06723_/A _12696_/B vssd1 vssd1 vccd1 vccd1 _06666_/Y sky130_fd_sc_hd__nor2_1
X_09454_ _09624_/A _09454_/B vssd1 vssd1 vccd1 vccd1 _09458_/B sky130_fd_sc_hd__or2_1
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09385_ _09381_/X _09384_/X _10294_/S vssd1 vssd1 vccd1 vccd1 _09385_/X sky130_fd_sc_hd__mux2_1
X_08405_ _08405_/A _08405_/B vssd1 vssd1 vccd1 vccd1 _08407_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_19_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06597_ instruction[18] _06944_/B vssd1 vssd1 vccd1 vccd1 _06597_/X sky130_fd_sc_hd__or2_1
XFILLER_0_47_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08336_ _08656_/A _08336_/B vssd1 vssd1 vccd1 vccd1 _08342_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__07618__B1 _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08267_ _08266_/B _08267_/B vssd1 vssd1 vccd1 vccd1 _08268_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_116_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07218_ _07213_/B _07213_/A _11584_/A vssd1 vssd1 vccd1 vccd1 _07218_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_6_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08198_ _08198_/A _08198_/B vssd1 vssd1 vccd1 vccd1 _08265_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_21_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09268__A _09922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07149_ _07149_/A _07149_/B vssd1 vssd1 vccd1 vccd1 _07149_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10207__A _10207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10160_ _09564_/X _09566_/X _10295_/S vssd1 vssd1 vccd1 vccd1 _10160_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09791__B1 _10240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12422__A _12422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10091_ _11868_/A fanout36/X fanout33/X fanout61/X vssd1 vssd1 vccd1 vccd1 _10092_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12142__A2 _12447_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11038__A _11038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10993_ _10993_/A _10993_/B vssd1 vssd1 vccd1 vccd1 _10995_/B sky130_fd_sc_hd__xor2_1
X_12801_ hold3/X hold67/X vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__nand2_1
XANTENNA__08649__A2 _08649_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10456__A2 _08289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11653__A1 _12421_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _12732_/A _12732_/B vssd1 vssd1 vccd1 vccd1 _12739_/C sky130_fd_sc_hd__nand2_4
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _12662_/A _12659_/Y _12661_/B vssd1 vssd1 vccd1 vccd1 _12667_/A sky130_fd_sc_hd__o21a_2
X_11614_ _11616_/A _11616_/B _11616_/C vssd1 vssd1 vccd1 vccd1 _11617_/A sky130_fd_sc_hd__a21o_1
X_12594_ _12633_/A _12595_/B vssd1 vssd1 vccd1 vccd1 _12596_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_108_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10208__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07609__B1 _07608_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11545_ _11545_/A _11545_/B vssd1 vssd1 vccd1 vccd1 _11547_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11476_ _11476_/A _12335_/B _11591_/A vssd1 vssd1 vccd1 vccd1 _11600_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_107_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13215_ _13249_/A hold255/X vssd1 vssd1 vccd1 vccd1 _13384_/D sky130_fd_sc_hd__and2_1
XANTENNA__06719__A_N _07097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10427_ reg1_val[8] curr_PC[8] vssd1 vssd1 vccd1 vccd1 _10428_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08034__B1 _10476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10358_ _11393_/A _10358_/B vssd1 vssd1 vccd1 vccd1 _10362_/A sky130_fd_sc_hd__xnor2_1
X_13146_ hold294/X _12803_/B _13145_/X _12804_/A vssd1 vssd1 vccd1 vccd1 _13147_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13077_ _11582_/A _13101_/B2 hold114/X vssd1 vssd1 vccd1 vccd1 hold115/A sky130_fd_sc_hd__o21a_1
X_10289_ _06830_/Y _10288_/Y _12054_/S vssd1 vssd1 vccd1 vccd1 _10291_/B sky130_fd_sc_hd__mux2_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12028_ _12108_/A _12028_/B vssd1 vssd1 vccd1 vccd1 _12030_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08337__B2 _08641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08337__A1 _08627_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12478__S _12520_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06984__B _06984_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11644__A1 _12064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07848__B1 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08257__A _08564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07161__A _09779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09170_ reg1_val[9] reg1_val[22] _09180_/S vssd1 vssd1 vccd1 vccd1 _09170_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11947__A2 _12009_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08121_ _08121_/A _08121_/B vssd1 vssd1 vccd1 vccd1 _08162_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_16_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12507__A _12675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08052_ _08649_/B1 _08112_/B fanout25/X _09404_/S vssd1 vssd1 vccd1 vccd1 _08053_/B
+ sky130_fd_sc_hd__o22a_1
X_07003_ reg1_val[4] _07083_/C _07248_/A vssd1 vssd1 vccd1 vccd1 _07004_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_3_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08576__A1 _08641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12372__A2 _12447_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08576__B2 _08627_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08954_ _08954_/A _08954_/B vssd1 vssd1 vccd1 vccd1 _08957_/B sky130_fd_sc_hd__xor2_1
X_07905_ _08334_/A _07905_/B vssd1 vssd1 vccd1 vccd1 _07968_/B sky130_fd_sc_hd__xnor2_2
X_08885_ _10871_/A _08112_/B fanout25/X _07198_/Y vssd1 vssd1 vccd1 vccd1 _08886_/B
+ sky130_fd_sc_hd__o22a_1
X_07836_ _09947_/A _07836_/B vssd1 vssd1 vccd1 vccd1 _07837_/C sky130_fd_sc_hd__xnor2_1
X_07767_ _07824_/A _07766_/Y _07762_/Y vssd1 vssd1 vccd1 vccd1 _07781_/A sky130_fd_sc_hd__a21oi_2
X_06718_ reg2_val[17] _06766_/B _06724_/B1 _06717_/Y vssd1 vssd1 vccd1 vccd1 _07097_/A
+ sky130_fd_sc_hd__o2bb2a_4
X_09506_ _09507_/A _09507_/B vssd1 vssd1 vccd1 vccd1 _09506_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07839__B1 _09661_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07071__A _07907_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07698_ _07701_/A _07701_/B vssd1 vssd1 vccd1 vccd1 _07698_/X sky130_fd_sc_hd__or2_1
XFILLER_0_109_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06649_ reg2_val[25] _06766_/B _06677_/B1 _06648_/Y vssd1 vssd1 vccd1 vccd1 _06998_/A
+ sky130_fd_sc_hd__o2bb2a_4
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09437_ _11138_/A _09436_/A _09249_/Y vssd1 vssd1 vccd1 vccd1 _09437_/Y sky130_fd_sc_hd__a21oi_2
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09368_ _09368_/A _09368_/B vssd1 vssd1 vccd1 vccd1 _09369_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_117_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout18_A _12009_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09299_ _09673_/A _09299_/B vssd1 vssd1 vccd1 vccd1 _09307_/A sky130_fd_sc_hd__xor2_1
X_08319_ _08316_/A _08316_/B _08318_/Y vssd1 vssd1 vccd1 vccd1 _08328_/A sky130_fd_sc_hd__o21ai_1
X_11330_ _11331_/A _11331_/B _11331_/C vssd1 vssd1 vccd1 vccd1 _11330_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA_60 _09661_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11261_ _07262_/A _12422_/A _11258_/Y _11260_/Y vssd1 vssd1 vccd1 vccd1 _11264_/A
+ sky130_fd_sc_hd__a211o_1
X_11192_ _11393_/A _11192_/B vssd1 vssd1 vccd1 vccd1 _11193_/B sky130_fd_sc_hd__xnor2_2
X_13000_ hold169/X _13000_/A2 _13257_/A2 _13310_/Q vssd1 vssd1 vccd1 vccd1 hold170/A
+ sky130_fd_sc_hd__a22o_1
X_10212_ _10212_/A _10212_/B vssd1 vssd1 vccd1 vccd1 _10215_/A sky130_fd_sc_hd__or2_1
X_10143_ _10143_/A _10143_/B vssd1 vssd1 vccd1 vccd1 _10143_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_30_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_17 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10074_ _10075_/A _10075_/B vssd1 vssd1 vccd1 vccd1 _10224_/A sky130_fd_sc_hd__and2_1
XFILLER_0_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10976_ _10976_/A _10976_/B _10976_/C vssd1 vssd1 vccd1 vccd1 _10984_/A sky130_fd_sc_hd__or3_1
XFILLER_0_97_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12715_ _12721_/A _12715_/B vssd1 vssd1 vccd1 vccd1 _12717_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_127_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12646_ _12646_/A _12646_/B vssd1 vssd1 vccd1 vccd1 _12647_/B sky130_fd_sc_hd__nand2_2
XANTENNA__12051__A1 _11892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12577_ _12582_/B _12577_/B vssd1 vssd1 vccd1 vccd1 new_PC[17] sky130_fd_sc_hd__xnor2_4
XANTENNA__06970__D _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10601__A2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11528_ _11528_/A _11712_/A vssd1 vssd1 vccd1 vccd1 _11528_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_53_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13000__B1 _13257_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11459_ _06719_/X _11995_/B _11457_/Y _06721_/B _11458_/Y vssd1 vssd1 vccd1 vccd1
+ _11459_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08540__A _09404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13129_ _13129_/A _13129_/B vssd1 vssd1 vccd1 vccd1 _13129_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12997__A _13001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08670_ _08719_/A _08719_/B _08653_/X vssd1 vssd1 vccd1 vccd1 _08721_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_17_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09371__A _09371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07621_ fanout61/X _10245_/B2 _10245_/A1 fanout53/X vssd1 vssd1 vccd1 vccd1 _07622_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11406__A _11406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07552_ fanout46/X _09325_/A _07172_/Y _07830_/B vssd1 vssd1 vccd1 vccd1 _07553_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07483_ _08656_/A _07483_/B vssd1 vssd1 vccd1 vccd1 _07682_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09222_ _11813_/S _09222_/B vssd1 vssd1 vccd1 vccd1 _09222_/Y sky130_fd_sc_hd__nand2_8
XFILLER_0_63_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09153_ _12438_/A _09222_/B vssd1 vssd1 vccd1 vccd1 _09153_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_8_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11141__A _11820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10053__B1 _07282_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08104_ _08334_/A _08104_/B vssd1 vssd1 vccd1 vccd1 _08108_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11250__C1 _06946_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09084_ _09085_/A _09085_/B vssd1 vssd1 vccd1 vccd1 _09084_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_102_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08035_ _10207_/A _08035_/B vssd1 vssd1 vccd1 vccd1 _08081_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09546__A _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11553__A0 _11829_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07066__A _09947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09986_ _09854_/A _09854_/B _09852_/Y vssd1 vssd1 vccd1 vccd1 _09993_/A sky130_fd_sc_hd__a21o_1
X_08937_ _08937_/A _08937_/B vssd1 vssd1 vccd1 vccd1 _08939_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_99_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08868_ _08868_/A _08868_/B vssd1 vssd1 vccd1 vccd1 _08869_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07524__A2 _09661_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07819_ _07819_/A _07819_/B vssd1 vssd1 vccd1 vccd1 _07874_/A sky130_fd_sc_hd__xnor2_1
X_08799_ _08805_/A _08799_/B _08799_/C vssd1 vssd1 vccd1 vccd1 _08800_/B sky130_fd_sc_hd__nand3_1
X_10830_ _10834_/A vssd1 vssd1 vccd1 vccd1 _10833_/A sky130_fd_sc_hd__inv_2
XFILLER_0_67_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10761_ _10636_/A _10635_/B _10635_/A vssd1 vssd1 vccd1 vccd1 _10766_/A sky130_fd_sc_hd__o21bai_2
XANTENNA__12281__B2 _12335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12281__A1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07288__B2 _08112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07288__A1 _07217_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10692_ hold279/A _12271_/A1 _10810_/B _10691_/Y _12376_/C1 vssd1 vssd1 vccd1 vccd1
+ _10692_/X sky130_fd_sc_hd__a311o_1
XANTENNA__10831__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12500_ _12670_/B _12501_/B vssd1 vssd1 vccd1 vccd1 _12511_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_66_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12431_ _12348_/B _12392_/Y _12394_/B vssd1 vssd1 vccd1 vccd1 _12431_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10595__A1 _10595_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12362_ _06673_/A _12360_/X _12361_/Y vssd1 vssd1 vccd1 vccd1 _12381_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__06799__B1 _06797_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11313_ _11313_/A _11313_/B vssd1 vssd1 vccd1 vccd1 _11326_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__10595__B2 _07198_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12293_ _12346_/A _12292_/C _12292_/A vssd1 vssd1 vccd1 vccd1 _12294_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_120_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11244_ _11137_/A _11137_/B _11135_/A vssd1 vssd1 vccd1 vccd1 _11245_/B sky130_fd_sc_hd__o21a_1
XANTENNA__09737__B1 _12064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09456__A _09779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10347__B2 _10473_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11175_ _11318_/B _11175_/B vssd1 vssd1 vccd1 vccd1 _11196_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10126_ _10124_/A _10124_/B _10127_/B vssd1 vssd1 vccd1 vccd1 _10126_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__08960__A1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08960__B2 _09661_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10057_ _12233_/A fanout86/X fanout82/X _12087_/A vssd1 vssd1 vccd1 vccd1 _10058_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09504__A3 _12158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap118_A _07195_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13049__B1 _09302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10959_ _12233_/B fanout28/X fanout26/X _12233_/A vssd1 vssd1 vccd1 vccd1 _10960_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06981__C _07097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12629_ _12633_/A _12620_/B _12624_/A _12624_/B vssd1 vssd1 vccd1 vccd1 _12630_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_110_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold105 hold105/A vssd1 vssd1 vccd1 vccd1 hold105/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 hold143/X vssd1 vssd1 vccd1 vccd1 hold116/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold138 hold138/A vssd1 vssd1 vccd1 vccd1 hold138/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12327__A2 _09228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold127 hold200/X vssd1 vssd1 vccd1 vccd1 hold127/X sky130_fd_sc_hd__buf_1
Xhold149 hold149/A vssd1 vssd1 vccd1 vccd1 hold149/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10338__A1 _10595_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10338__B2 _10338_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11535__B1 _12356_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09840_ _09683_/A _09683_/B _09681_/Y vssd1 vssd1 vccd1 vccd1 _09842_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_0_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06983_ _06983_/A _06983_/B _06983_/C vssd1 vssd1 vccd1 vccd1 _07070_/A sky130_fd_sc_hd__nand3_4
X_09771_ _09936_/A _09771_/B vssd1 vssd1 vccd1 vccd1 _09775_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08951__B2 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08951__A1 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08722_ _10010_/B _10010_/C vssd1 vssd1 vccd1 vccd1 _10151_/B sky130_fd_sc_hd__and2_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09900__B1 _11554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout172_A _12826_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08653_ _08654_/B _08654_/A vssd1 vssd1 vccd1 vccd1 _08653_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09259__A2 _09257_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08584_ _08605_/A vssd1 vssd1 vccd1 vccd1 _08584_/Y sky130_fd_sc_hd__inv_2
X_07604_ _07604_/A _07604_/B vssd1 vssd1 vccd1 vccd1 _07615_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_119_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07535_ _07535_/A _07535_/B vssd1 vssd1 vccd1 vccd1 _07537_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_91_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07466_ _07466_/A _07466_/B vssd1 vssd1 vccd1 vccd1 _07495_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_107_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09205_ _09203_/X _09204_/X _09403_/S vssd1 vssd1 vccd1 vccd1 _09205_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07397_ _09341_/A _07397_/B vssd1 vssd1 vccd1 vccd1 _07434_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10577__A1 _12446_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09431__A2 _08664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09136_ _09136_/A _09136_/B vssd1 vssd1 vccd1 vccd1 _09137_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_114_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10914__S _11029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09067_ _09278_/A _09067_/B vssd1 vssd1 vccd1 vccd1 _09069_/B sky130_fd_sc_hd__and2_1
XFILLER_0_102_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08018_ _08598_/B _10595_/A1 _10338_/B2 _08538_/A1 vssd1 vssd1 vccd1 vccd1 _08019_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09969_ _10092_/A _09969_/B vssd1 vssd1 vccd1 vccd1 _09973_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09215__S _11138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12980_ hold237/A _13000_/A2 _13257_/A2 hold221/X vssd1 vssd1 vccd1 vccd1 hold222/A
+ sky130_fd_sc_hd__a22o_1
X_11931_ _12093_/A _11931_/B vssd1 vssd1 vccd1 vccd1 _11932_/B sky130_fd_sc_hd__xnor2_1
X_11862_ _11776_/A _11776_/B _11767_/A vssd1 vssd1 vccd1 vccd1 _11874_/A sky130_fd_sc_hd__o21ai_1
X_10813_ _10813_/A _12422_/A vssd1 vssd1 vccd1 vccd1 _10813_/Y sky130_fd_sc_hd__nand2_1
X_11793_ _11793_/A _11793_/B _11793_/C vssd1 vssd1 vccd1 vccd1 _11794_/B sky130_fd_sc_hd__or3_1
XFILLER_0_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10744_ _10476_/A fanout12/X fanout7/X _08411_/B vssd1 vssd1 vccd1 vccd1 _10745_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12006__A1 _11929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10675_ reg1_val[10] curr_PC[10] vssd1 vssd1 vccd1 vccd1 _10679_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_40_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12414_ hold258/A _12414_/B vssd1 vssd1 vccd1 vccd1 _12414_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13394_ _13396_/CLK hold168/X vssd1 vssd1 vccd1 vccd1 hold298/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09885__S _11138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12345_ _12345_/A _12345_/B vssd1 vssd1 vccd1 vccd1 _12346_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12276_ _09221_/Y _09880_/Y _09886_/X _12379_/B2 _12275_/Y vssd1 vssd1 vccd1 vccd1
+ _12277_/C sky130_fd_sc_hd__a221o_1
XANTENNA__08090__A _08664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11227_ _11227_/A _11333_/A vssd1 vssd1 vccd1 vccd1 _11434_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12190__B1 _11637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11158_ _12365_/A _11127_/X _11128_/X _11157_/X _11126_/X vssd1 vssd1 vccd1 vccd1
+ _11158_/X sky130_fd_sc_hd__a311o_1
X_10109_ _10944_/B2 fanout32/X fanout30/X _07097_/X vssd1 vssd1 vccd1 vccd1 _10110_/B
+ sky130_fd_sc_hd__a22o_1
X_11089_ _11309_/A fanout10/X fanout5/X _11198_/A vssd1 vssd1 vccd1 vccd1 _11090_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10779__B _10900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09489__A2 fanout86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11296__A2 _07171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06992__B _12644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07320_ _09669_/B2 fanout59/X fanout57/X _09301_/A vssd1 vssd1 vccd1 vccd1 _07321_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09661__A2 _08199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07251_ reg1_val[11] _07248_/B _07585_/B1 vssd1 vssd1 vccd1 vccd1 _07252_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_6_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07182_ _11134_/A _11242_/A reg1_val[16] _07141_/C _07585_/B1 vssd1 vssd1 vccd1 vccd1
+ _07184_/B sky130_fd_sc_hd__o41a_4
XFILLER_0_60_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11756__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12515__A _12680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09823_ _09673_/A _09673_/B _09671_/Y vssd1 vssd1 vccd1 vccd1 _09827_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__10731__B2 _07013_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10731__A1 _11946_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09754_ _06800_/Y _12144_/A1 _12420_/A0 _09745_/B _09753_/X vssd1 vssd1 vccd1 vccd1
+ _09754_/X sky130_fd_sc_hd__o221a_1
X_06966_ _12644_/A _06967_/B vssd1 vssd1 vccd1 vccd1 _09671_/A sky130_fd_sc_hd__xor2_4
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06897_ _11239_/A _11131_/A _11022_/A _06897_/D vssd1 vssd1 vccd1 vccd1 _06900_/B
+ sky130_fd_sc_hd__and4bb_1
X_09685_ _09685_/A _09685_/B vssd1 vssd1 vccd1 vccd1 _09686_/B sky130_fd_sc_hd__xor2_2
X_08705_ _08706_/A _08706_/B vssd1 vssd1 vccd1 vccd1 _08802_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_96_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08636_ _08630_/A _08630_/B _08628_/Y vssd1 vssd1 vccd1 vccd1 _08637_/C sky130_fd_sc_hd__o21ba_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout11 _08876_/Y vssd1 vssd1 vccd1 vccd1 _08877_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout22 _12428_/B vssd1 vssd1 vccd1 vccd1 _11946_/C sky130_fd_sc_hd__clkbuf_16
X_08567_ _08567_/A _08567_/B vssd1 vssd1 vccd1 vccd1 _08568_/C sky130_fd_sc_hd__xor2_2
Xfanout55 fanout56/X vssd1 vssd1 vccd1 vccd1 _12233_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout44 _07157_/Y vssd1 vssd1 vccd1 vccd1 _07417_/B sky130_fd_sc_hd__buf_6
X_08498_ _08498_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _08500_/B sky130_fd_sc_hd__xnor2_1
Xfanout33 _07201_/X vssd1 vssd1 vccd1 vccd1 fanout33/X sky130_fd_sc_hd__buf_8
X_07518_ _07518_/A _07518_/B vssd1 vssd1 vccd1 vccd1 _07734_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout66 _06997_/Y vssd1 vssd1 vccd1 vccd1 _12087_/A sky130_fd_sc_hd__buf_4
XFILLER_0_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout99 _07096_/Y vssd1 vssd1 vccd1 vccd1 _11406_/A sky130_fd_sc_hd__buf_4
Xfanout77 _07270_/X vssd1 vssd1 vccd1 vccd1 _11093_/A sky130_fd_sc_hd__buf_6
X_07449_ _10871_/A fanout82/X _10974_/A fanout86/X vssd1 vssd1 vccd1 vccd1 _07450_/B
+ sky130_fd_sc_hd__o22a_1
Xfanout88 _11284_/A vssd1 vssd1 vccd1 vccd1 _09341_/A sky130_fd_sc_hd__buf_12
X_10460_ _10461_/A _10461_/B vssd1 vssd1 vccd1 vccd1 _10618_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09119_ _09119_/A _09119_/B vssd1 vssd1 vccd1 vccd1 _09122_/A sky130_fd_sc_hd__xor2_2
XANTENNA__07415__A1 _07830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10391_ _11868_/A fanout28/X fanout26/X fanout62/X vssd1 vssd1 vccd1 vccd1 _10392_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08612__B1 _06992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07415__B2 _08576_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12130_ _12063_/A _12060_/Y _12062_/B vssd1 vssd1 vccd1 vccd1 _12134_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_102_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12061_ reg1_val[24] curr_PC[24] vssd1 vssd1 vccd1 vccd1 _12062_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11012_ _10546_/X _11009_/A _11229_/A _11011_/X vssd1 vssd1 vccd1 vccd1 _11012_/Y
+ sky130_fd_sc_hd__a31oi_1
XANTENNA__07718__A2 _08289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10599__B _12087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12963_ hold60/X hold284/X vssd1 vssd1 vccd1 vccd1 _13229_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07254__A _10749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_28 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11914_ _12421_/A1 _11913_/X _06686_/B vssd1 vssd1 vccd1 vccd1 _11914_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09340__A1 _08112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09340__B2 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12894_ hold285/A hold106/X vssd1 vssd1 vccd1 vccd1 _13163_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_68_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ _07051_/X fanout41/X _07316_/Y fanout43/X vssd1 vssd1 vccd1 vccd1 _11846_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_68_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _11776_/A _11776_/B vssd1 vssd1 vccd1 vccd1 _11790_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_83_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10727_ _10728_/A _10728_/B vssd1 vssd1 vccd1 vccd1 _10727_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__12319__B _12319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08851__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10658_ _10658_/A _10658_/B vssd1 vssd1 vccd1 vccd1 _10658_/X sky130_fd_sc_hd__and2_1
XFILLER_0_51_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07406__A1 _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13377_ _13379_/CLK _13377_/D vssd1 vssd1 vccd1 vccd1 hold292/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10589_ _07417_/B _07256_/Y _07262_/X fanout41/X vssd1 vssd1 vccd1 vccd1 _10590_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12335__A _12335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10554__S _12054_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07406__B2 _08613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12328_ _06630_/X _11995_/B _12327_/Y _06632_/B _12422_/A vssd1 vssd1 vccd1 vccd1
+ _12328_/X sky130_fd_sc_hd__a221o_1
XANTENNA__11753__A3 _11720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07957__A2 _08199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12259_ _12192_/X _12193_/Y _12195_/B vssd1 vssd1 vccd1 vccd1 _12259_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_76_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10713__A1 _07097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10713__B2 _07256_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06820_ _09418_/A _09418_/B _06819_/X vssd1 vssd1 vccd1 vccd1 _06820_/X sky130_fd_sc_hd__a21o_1
X_06751_ reg1_val[11] _10813_/A vssd1 vssd1 vccd1 vccd1 _10808_/S sky130_fd_sc_hd__and2_1
X_06682_ _06723_/A _12675_/B vssd1 vssd1 vccd1 vccd1 _06682_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10477__B1 _10207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09470_ _09471_/A _09471_/B vssd1 vssd1 vccd1 vccd1 _09621_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__08134__A2 _10221_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08421_ _08421_/A _08421_/B vssd1 vssd1 vccd1 vccd1 _08423_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07893__A1 _07148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07893__B2 _07959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09095__B1 _09672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08352_ _08352_/A _08352_/B vssd1 vssd1 vccd1 vccd1 _08405_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08283_ _08283_/A _08283_/B vssd1 vssd1 vccd1 vccd1 _08323_/A sky130_fd_sc_hd__xnor2_1
X_07303_ _09667_/A _07303_/B vssd1 vssd1 vccd1 vccd1 _07306_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07234_ _07212_/A _07212_/B _07230_/B _11381_/A vssd1 vssd1 vccd1 vccd1 _07234_/Y
+ sky130_fd_sc_hd__a211oi_2
XANTENNA_fanout135_A _08454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07165_ _07165_/A _07166_/B vssd1 vssd1 vccd1 vccd1 _07165_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07096_ _07097_/A _07097_/B vssd1 vssd1 vccd1 vccd1 _07096_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_42_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout223 _07165_/A vssd1 vssd1 vccd1 vccd1 _11028_/S sky130_fd_sc_hd__buf_2
Xfanout212 _09419_/B vssd1 vssd1 vccd1 vccd1 _09383_/S sky130_fd_sc_hd__clkbuf_4
Xfanout201 _10243_/A vssd1 vssd1 vccd1 vccd1 _08580_/A sky130_fd_sc_hd__buf_12
Xfanout234 _09423_/X vssd1 vssd1 vccd1 vccd1 _12271_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout245 _12631_/S vssd1 vssd1 vccd1 vccd1 _12638_/S sky130_fd_sc_hd__clkbuf_8
Xfanout256 _13000_/A2 vssd1 vssd1 vccd1 vccd1 _12804_/A sky130_fd_sc_hd__clkbuf_4
Xfanout278 _06585_/Y vssd1 vssd1 vccd1 vccd1 _13001_/A sky130_fd_sc_hd__buf_4
Xfanout267 _06783_/A vssd1 vssd1 vccd1 vccd1 _06766_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__10180__A2 _12446_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09806_ _09806_/A _09807_/B vssd1 vssd1 vccd1 vccd1 _09931_/A sky130_fd_sc_hd__nor2_1
Xfanout289 reg1_val[1] vssd1 vssd1 vccd1 vccd1 _12644_/A sky130_fd_sc_hd__buf_12
XANTENNA__08373__A2 _08457_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07998_ _08006_/A _08006_/B vssd1 vssd1 vccd1 vccd1 _08009_/A sky130_fd_sc_hd__nand2b_1
X_06949_ _06949_/A instruction[4] vssd1 vssd1 vccd1 vccd1 _09237_/B sky130_fd_sc_hd__nand2_2
X_09737_ _09733_/X _09736_/X _12064_/S vssd1 vssd1 vccd1 vccd1 _09737_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout48_A _07131_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09668_ _09668_/A _09668_/B vssd1 vssd1 vccd1 vccd1 _09675_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07333__B1 _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ _06809_/Y _12420_/A0 _09589_/Y _09598_/X vssd1 vssd1 vccd1 vccd1 _09599_/X
+ sky130_fd_sc_hd__o211a_1
X_08619_ _08619_/A _08619_/B vssd1 vssd1 vccd1 vccd1 _08625_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_77_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09086__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11630_ _11630_/A _11630_/B _11630_/C vssd1 vssd1 vccd1 vccd1 _11631_/B sky130_fd_sc_hd__or3_1
XFILLER_0_126_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11561_ _09242_/B _11548_/X _11560_/X vssd1 vssd1 vccd1 vccd1 _11561_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09625__A2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07636__B2 _07134_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07636__A1 _07121_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10512_ fanout52/X fanout47/X fanout45/X _11476_/A vssd1 vssd1 vccd1 vccd1 _10513_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_80_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13300_ _13304_/CLK hold223/X vssd1 vssd1 vccd1 vccd1 hold221/A sky130_fd_sc_hd__dfxtp_1
X_11492_ _11492_/A _11492_/B vssd1 vssd1 vccd1 vccd1 _11493_/B sky130_fd_sc_hd__or2_1
XFILLER_0_33_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13231_ hold284/A _13230_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13231_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_107_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10443_ _10435_/Y _10436_/X _10442_/X vssd1 vssd1 vccd1 vccd1 _10443_/X sky130_fd_sc_hd__o21a_1
X_13162_ _13162_/A hold286/X vssd1 vssd1 vccd1 vccd1 _13373_/D sky130_fd_sc_hd__and2_1
X_10374_ _10501_/A _10501_/B vssd1 vssd1 vccd1 vccd1 _10376_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12113_ _12113_/A _12300_/A vssd1 vssd1 vccd1 vccd1 _12114_/B sky130_fd_sc_hd__nor2_1
XANTENNA__12145__B1 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13093_ _12224_/A _13101_/B2 hold117/X vssd1 vssd1 vccd1 vccd1 hold118/A sky130_fd_sc_hd__o21a_1
X_12044_ _11883_/A _11964_/A _11963_/A vssd1 vssd1 vccd1 vccd1 _12044_/Y sky130_fd_sc_hd__a21oi_1
X_12946_ _13193_/A _13194_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13198_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_99_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12877_ hold284/X hold60/X vssd1 vssd1 vccd1 vccd1 _13229_/A sky130_fd_sc_hd__nand2b_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ hold188/A _11990_/A1 _11907_/B _11648_/A vssd1 vssd1 vccd1 vccd1 _11828_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12049__B _12049_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11759_ _12096_/A _11759_/B vssd1 vssd1 vccd1 vccd1 _11760_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_83_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13176__A2 _13223_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12384__B1 _12335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08052__B2 _09404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08052__A1 _08649_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06998__A _06998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08970_ _09064_/B _08970_/B vssd1 vssd1 vccd1 vccd1 _08983_/A sky130_fd_sc_hd__nand2_1
X_07921_ _10243_/A _07921_/B vssd1 vssd1 vccd1 vccd1 _07924_/A sky130_fd_sc_hd__xnor2_1
X_07852_ _10246_/A _07852_/B vssd1 vssd1 vccd1 vccd1 _07887_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12439__A1 _12438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06803_ reg2_val[2] _06810_/B vssd1 vssd1 vccd1 vccd1 _06803_/X sky130_fd_sc_hd__and2_2
XANTENNA__13100__A2 _06577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09522_ _09522_/A _09522_/B vssd1 vssd1 vccd1 vccd1 _09525_/A sky130_fd_sc_hd__xnor2_1
X_07783_ _07753_/Y _07756_/X _07802_/B vssd1 vssd1 vccd1 vccd1 _07783_/X sky130_fd_sc_hd__a21o_1
X_06734_ reg2_val[14] _06810_/B vssd1 vssd1 vccd1 vccd1 _06734_/X sky130_fd_sc_hd__and2_1
XFILLER_0_78_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06665_ instruction[36] _06675_/B vssd1 vssd1 vccd1 vccd1 _12696_/B sky130_fd_sc_hd__and2_4
X_09453_ _09452_/B _09453_/B vssd1 vssd1 vccd1 vccd1 _09454_/B sky130_fd_sc_hd__and2b_1
XANTENNA__07622__A _10479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09384_ _09382_/X _09383_/X _09725_/S vssd1 vssd1 vccd1 vccd1 _09384_/X sky130_fd_sc_hd__mux2_1
X_08404_ _08403_/A _08403_/B _08403_/C vssd1 vssd1 vccd1 vccd1 _08433_/B sky130_fd_sc_hd__a21o_1
X_06596_ instruction[14] _06590_/X _06595_/X _06716_/B vssd1 vssd1 vccd1 vccd1 reg1_idx[3]
+ sky130_fd_sc_hd__o211a_4
XFILLER_0_108_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08335_ _07983_/A _07195_/X _07274_/Y _12642_/A vssd1 vssd1 vccd1 vccd1 _08336_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07618__A1 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07618__B2 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10622__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08266_ _08267_/B _08266_/B vssd1 vssd1 vccd1 vccd1 _08268_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_117_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07217_ _07215_/A _07214_/X _07215_/Y _06983_/A vssd1 vssd1 vccd1 vccd1 _07217_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_0_61_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08197_ _08193_/A _08193_/B _08264_/A vssd1 vssd1 vccd1 vccd1 _08211_/A sky130_fd_sc_hd__o21ba_1
X_07148_ _09728_/S _07149_/B vssd1 vssd1 vccd1 vccd1 _07148_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__09791__A1 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09240__B1 _09238_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09791__B2 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07079_ _07080_/A _07080_/B vssd1 vssd1 vccd1 vccd1 _07079_/X sky130_fd_sc_hd__and2_2
X_10090_ _09923_/A _09923_/B _09920_/A vssd1 vssd1 vccd1 vccd1 _10102_/A sky130_fd_sc_hd__a21o_1
XANTENNA__11038__B _12422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12800_ hold67/X vssd1 vssd1 vccd1 vccd1 _12800_/Y sky130_fd_sc_hd__inv_2
X_10992_ _10990_/A _10990_/B _10993_/B vssd1 vssd1 vccd1 vccd1 _11108_/A sky130_fd_sc_hd__a21o_1
XANTENNA__08628__A _09302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12731_ reg1_val[18] _12755_/B vssd1 vssd1 vccd1 vccd1 _12732_/B sky130_fd_sc_hd__or2_1
XANTENNA__10861__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _12662_/A _12662_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[4] sky130_fd_sc_hd__xnor2_4
XFILLER_0_32_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11613_ _11613_/A _11613_/B vssd1 vssd1 vccd1 vccd1 _11616_/C sky130_fd_sc_hd__or2_1
XFILLER_0_65_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12593_ reg1_val[20] curr_PC[20] _12638_/S vssd1 vssd1 vccd1 vccd1 _12595_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07609__B2 _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11544_ reg1_val[18] curr_PC[18] vssd1 vssd1 vccd1 vccd1 _11545_/B sky130_fd_sc_hd__or2_1
XFILLER_0_25_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11475_ _11476_/A _12335_/B _11591_/A vssd1 vssd1 vccd1 vccd1 _11477_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_80_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13214_ hold254/X _13223_/A2 _13213_/X _13223_/B2 vssd1 vssd1 vccd1 vccd1 hold255/A
+ sky130_fd_sc_hd__a22o_1
X_10426_ reg1_val[8] curr_PC[8] vssd1 vssd1 vccd1 vccd1 _10426_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08034__A1 _09770_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08034__B2 _09940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10357_ _11476_/A fanout47/X fanout45/X _11406_/A vssd1 vssd1 vccd1 vccd1 _10358_/B
+ sky130_fd_sc_hd__o22a_1
X_13145_ hold252/X _13144_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13145_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13076_ hold133/A _12805_/A _13101_/A2 hold113/X _13259_/A vssd1 vssd1 vccd1 vccd1
+ hold114/A sky130_fd_sc_hd__o221a_1
X_10288_ _06781_/A _10153_/Y _06779_/X vssd1 vssd1 vccd1 vccd1 _10288_/Y sky130_fd_sc_hd__a21oi_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12027_ _12027_/A _12027_/B _12027_/C vssd1 vssd1 vccd1 vccd1 _12028_/B sky130_fd_sc_hd__or3_1
XANTENNA__08337__A2 _10221_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09922__A _09922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09298__B1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12841__A1 _07256_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12929_ _13148_/A _13149_/A _13148_/B vssd1 vssd1 vccd1 vccd1 _13154_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__07848__B2 _08538_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07848__A1 _09943_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08120_ _08120_/A _08120_/B vssd1 vssd1 vccd1 vccd1 _08165_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_22_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10080__B2 _10225_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10080__A1 _10337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08051_ _08051_/A _08051_/B vssd1 vssd1 vccd1 vccd1 _08085_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07002_ _07248_/A _07083_/C vssd1 vssd1 vccd1 vccd1 _07008_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_24_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08576__A2 _08576_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07617__A _10749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08953_ _08954_/A _08954_/B vssd1 vssd1 vccd1 vccd1 _09066_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07904_ _08561_/A2 fanout75/X _09940_/B2 _08289_/B vssd1 vssd1 vccd1 vccd1 _07905_/B
+ sky130_fd_sc_hd__o22a_1
X_08884_ _07584_/A _07584_/B _07581_/A vssd1 vssd1 vccd1 vccd1 _08896_/A sky130_fd_sc_hd__a21oi_1
X_07835_ _09669_/B2 fanout98/X fanout84/X _09301_/A vssd1 vssd1 vccd1 vccd1 _07836_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13085__A1 _11929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07766_ _07824_/B vssd1 vssd1 vccd1 vccd1 _07766_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09289__B1 _10240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06717_ _06723_/A _12650_/B vssd1 vssd1 vccd1 vccd1 _06717_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09505_ _09505_/A _09505_/B vssd1 vssd1 vccd1 vccd1 _09507_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07839__A1 _09298_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07839__B2 _09298_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07071__B _07907_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09436_ _09436_/A vssd1 vssd1 vccd1 vccd1 _09436_/Y sky130_fd_sc_hd__inv_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07697_ _09947_/A _07697_/B vssd1 vssd1 vccd1 vccd1 _07701_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06648_ _06723_/A _12689_/B vssd1 vssd1 vccd1 vccd1 _06648_/Y sky130_fd_sc_hd__nor2_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06579_ instruction[6] vssd1 vssd1 vccd1 vccd1 _09233_/B sky130_fd_sc_hd__inv_2
X_09367_ _09368_/A _09368_/B vssd1 vssd1 vccd1 vccd1 _09367_/X sky130_fd_sc_hd__and2_1
XFILLER_0_105_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_50 reg1_val[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09298_ _09298_/A1 fanout13/X fanout8/X _09298_/B2 vssd1 vssd1 vccd1 vccd1 _09299_/B
+ sky130_fd_sc_hd__o22a_1
X_08318_ _08364_/A _08364_/B vssd1 vssd1 vccd1 vccd1 _08318_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_104_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_61 reg1_val[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08249_ _08313_/A _08313_/B _08245_/X vssd1 vssd1 vccd1 vccd1 _08260_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11260_ _12421_/A1 _11259_/X _06733_/B vssd1 vssd1 vccd1 vccd1 _11260_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11191_ _12087_/A fanout47/X fanout45/X _12009_/A vssd1 vssd1 vccd1 vccd1 _11192_/B
+ sky130_fd_sc_hd__o22a_1
X_10211_ _10211_/A _10211_/B vssd1 vssd1 vccd1 vccd1 _10212_/B sky130_fd_sc_hd__and2_1
X_10142_ _09546_/X _09705_/X _09706_/X _10331_/A _10542_/A vssd1 vssd1 vccd1 vccd1
+ _10143_/B sky130_fd_sc_hd__a2111oi_2
X_10073_ _07073_/X fanout8/X _10072_/Y _10243_/A vssd1 vssd1 vccd1 vccd1 _10075_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07262__A _07262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10975_ _10975_/A _10975_/B vssd1 vssd1 vccd1 vccd1 _10976_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12823__A1 _12823_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12714_ reg1_val[14] _12714_/B vssd1 vssd1 vccd1 vccd1 _12715_/B sky130_fd_sc_hd__or2_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12645_ reg1_val[1] _12645_/B vssd1 vssd1 vccd1 vccd1 _12646_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09047__A3 _08983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12576_ _12639_/A _12570_/B _12582_/A vssd1 vssd1 vccd1 vccd1 _12577_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_53_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11527_ _11528_/A _11712_/A vssd1 vssd1 vccd1 vccd1 _11527_/X sky130_fd_sc_hd__and2_1
XFILLER_0_53_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11458_ _07097_/A _09257_/S _12638_/S vssd1 vssd1 vccd1 vccd1 _11458_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09917__A _11393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11389_ _11389_/A _11389_/B vssd1 vssd1 vccd1 vccd1 _11401_/A sky130_fd_sc_hd__xnor2_1
X_10409_ _10409_/A _10409_/B vssd1 vssd1 vccd1 vccd1 _10411_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13128_ _13128_/A _13128_/B vssd1 vssd1 vccd1 vccd1 _13129_/B sky130_fd_sc_hd__nand2_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08540__B _08540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13059_ _07297_/B _12826_/B hold146/X vssd1 vssd1 vccd1 vccd1 _13339_/D sky130_fd_sc_hd__a21boi_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09652__A _09944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13067__A1 _07267_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09371__B _09371_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07620_ _07620_/A _07620_/B vssd1 vssd1 vccd1 vccd1 _07624_/A sky130_fd_sc_hd__xor2_2
XANTENNA__08191__B1 _10338_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11406__B _12017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11078__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07172__A _07172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07551_ _07959_/A _07554_/B vssd1 vssd1 vccd1 vccd1 _07706_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_124_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07482_ _06993_/A fanout59/X fanout57/X _08613_/A vssd1 vssd1 vccd1 vccd1 _07483_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09221_ _12359_/A _09221_/B vssd1 vssd1 vccd1 vccd1 _09221_/Y sky130_fd_sc_hd__nor2_8
XFILLER_0_63_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09152_ _12054_/S _09221_/B vssd1 vssd1 vccd1 vccd1 _09152_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_84_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08103_ _08561_/B1 _08289_/B fanout75/X _08576_/A2 vssd1 vssd1 vccd1 vccd1 _08104_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout215_A _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09083_ _10092_/A _09083_/B vssd1 vssd1 vccd1 vccd1 _09085_/B sky130_fd_sc_hd__xnor2_1
X_08034_ _09770_/B2 _08411_/B _10476_/A _09940_/B2 vssd1 vssd1 vccd1 vccd1 _08035_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09546__B _09548_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11553__A1 _11995_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07347__A _09834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09985_ _09847_/A _09846_/B _09844_/Y vssd1 vssd1 vccd1 vccd1 _09995_/A sky130_fd_sc_hd__a21o_1
X_08936_ _09922_/A _08936_/B vssd1 vssd1 vccd1 vccd1 _08937_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_98_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08867_ _08867_/A _08867_/B vssd1 vssd1 vccd1 vccd1 _08868_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_98_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07818_ _08708_/A _08708_/B _08706_/A _08706_/B vssd1 vssd1 vccd1 vccd1 _07818_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_08798_ _08799_/B _08799_/C _08805_/A vssd1 vssd1 vccd1 vccd1 _08800_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07082__A _09944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07749_ _07749_/A _07749_/B vssd1 vssd1 vccd1 vccd1 _07813_/B sky130_fd_sc_hd__xor2_1
X_10760_ _10620_/A _10620_/B _10637_/X vssd1 vssd1 vccd1 vccd1 _10770_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12281__A2 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout30_A _07218_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07288__A2 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10691_ _12271_/A1 _10810_/B hold279/A vssd1 vssd1 vccd1 vccd1 _10691_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09419_ _12054_/S _09419_/B vssd1 vssd1 vccd1 vccd1 _09419_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12428__A fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12430_ _12430_/A _12430_/B _12430_/C vssd1 vssd1 vccd1 vccd1 _12430_/X sky130_fd_sc_hd__or3_1
XFILLER_0_75_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10595__A2 _08877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12361_ _06673_/A _12360_/X _09225_/Y vssd1 vssd1 vccd1 vccd1 _12361_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11312_ _11313_/A _11313_/B vssd1 vssd1 vccd1 vccd1 _11312_/X sky130_fd_sc_hd__and2b_1
X_12292_ _12292_/A _12346_/A _12292_/C vssd1 vssd1 vccd1 vccd1 _12346_/B sky130_fd_sc_hd__nor3_1
XANTENNA__08641__A _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11243_ _11243_/A _11243_/B vssd1 vssd1 vccd1 vccd1 _11245_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_31_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10347__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11174_ _11174_/A _11174_/B vssd1 vssd1 vccd1 vccd1 _11175_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_100_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10125_ _09980_/A _09980_/B _09978_/Y vssd1 vssd1 vccd1 vccd1 _10127_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__08960__A2 fanout86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10056_ _10056_/A _10056_/B vssd1 vssd1 vccd1 vccd1 _10089_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09472__A _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13049__B2 _13101_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07920__B1 fanout72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10958_ _11929_/A _10958_/B vssd1 vssd1 vccd1 vccd1 _10962_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10807__B1 _12205_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12628_ _12628_/A _12628_/B vssd1 vssd1 vccd1 vccd1 _12630_/A sky130_fd_sc_hd__nor2_2
X_10889_ _10890_/A _10890_/B vssd1 vssd1 vccd1 vccd1 _10889_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__11242__A _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12559_ _12560_/A _12560_/B _12560_/C vssd1 vssd1 vccd1 vccd1 _12567_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_81_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold106 hold106/A vssd1 vssd1 vccd1 vccd1 hold106/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold117 hold117/A vssd1 vssd1 vccd1 vccd1 hold117/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12980__B1 _13257_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold139 hold139/A vssd1 vssd1 vccd1 vccd1 hold139/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 hold128/A vssd1 vssd1 vccd1 vccd1 hold128/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10338__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07203__A2 _07195_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06982_ _06983_/A _06983_/B _06983_/C vssd1 vssd1 vccd1 vccd1 _06987_/A sky130_fd_sc_hd__and3_4
X_09770_ _07217_/Y _07362_/B fanout16/X _09770_/B2 vssd1 vssd1 vccd1 vccd1 _09771_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08951__A2 _07068_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11299__B1 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08721_ _08721_/A _08721_/B vssd1 vssd1 vccd1 vccd1 _10010_/C sky130_fd_sc_hd__xnor2_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09900__A1 _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08652_ _08652_/A _08652_/B vssd1 vssd1 vccd1 vccd1 _08654_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07911__B1 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07603_ fanout68/X _09298_/A1 fanout56/X _09298_/B2 vssd1 vssd1 vccd1 vccd1 _07604_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout165_A _12447_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08583_ _08583_/A _08596_/A vssd1 vssd1 vccd1 vccd1 _08605_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_88_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07534_ _07534_/A _07534_/B vssd1 vssd1 vccd1 vccd1 _07535_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_49_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07465_ _07563_/B _07563_/A vssd1 vssd1 vccd1 vccd1 _07466_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_8_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07630__A _09779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09204_ reg1_val[12] reg1_val[19] _09211_/S vssd1 vssd1 vccd1 vccd1 _09204_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_60_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07396_ _07217_/Y _08112_/B fanout25/X _07221_/X vssd1 vssd1 vccd1 vccd1 _07397_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_115_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09135_ _09136_/A _09136_/B vssd1 vssd1 vccd1 vccd1 _09135_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_17_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09066_ _09066_/A _09066_/B _09066_/C vssd1 vssd1 vccd1 vccd1 _09067_/B sky130_fd_sc_hd__or3_1
XFILLER_0_4_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08017_ _08073_/A _08073_/B vssd1 vssd1 vccd1 vccd1 _08017_/X sky130_fd_sc_hd__and2_1
XFILLER_0_12_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09968_ fanout61/X fanout36/X fanout33/X fanout53/X vssd1 vssd1 vccd1 vccd1 _09969_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout78_A _08289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08919_ _07676_/A _07676_/B _08918_/X vssd1 vssd1 vccd1 vccd1 _08919_/X sky130_fd_sc_hd__a21o_1
X_11930_ _07175_/Y fanout12/X fanout7/X _07171_/Y vssd1 vssd1 vccd1 vccd1 _11931_/B
+ sky130_fd_sc_hd__o22a_1
X_09899_ _09899_/A _09899_/B vssd1 vssd1 vccd1 vccd1 _09899_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_87_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10231__A _11398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07902__B1 _10476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11861_ _11861_/A _11861_/B vssd1 vssd1 vccd1 vccd1 _11876_/A sky130_fd_sc_hd__nand2_1
X_11792_ _11793_/A _11793_/B _11793_/C vssd1 vssd1 vccd1 vccd1 _11881_/B sky130_fd_sc_hd__o21ai_1
X_10812_ hold288/A _12271_/A1 _10924_/B _12416_/C1 vssd1 vssd1 vccd1 vccd1 _10812_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10743_ _10597_/A _10597_/B _10599_/X vssd1 vssd1 vccd1 vccd1 _10756_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_67_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11062__A _11393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10674_ reg1_val[10] curr_PC[10] vssd1 vssd1 vccd1 vccd1 _10674_/X sky130_fd_sc_hd__and2_1
XFILLER_0_70_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12413_ _12412_/A _12411_/X _12412_/Y _12446_/C1 vssd1 vssd1 vccd1 vccd1 _12425_/C
+ sky130_fd_sc_hd__o211a_1
X_13393_ _13396_/CLK hold142/X vssd1 vssd1 vccd1 vccd1 hold305/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12344_ _12345_/A _12345_/B vssd1 vssd1 vccd1 vccd1 _12391_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__10568__A2 _11829_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08371__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12275_ _06643_/X _12273_/Y _12274_/X vssd1 vssd1 vccd1 vccd1 _12275_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11226_ _11007_/A _11118_/A _11118_/B vssd1 vssd1 vccd1 vccd1 _11226_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__07197__A1 _07233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11157_ _11157_/A _11157_/B _11156_/X vssd1 vssd1 vccd1 vccd1 _11157_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10108_ _11398_/A _10108_/B vssd1 vssd1 vccd1 vccd1 _10112_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07715__A _10092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11088_ _11088_/A _11088_/B vssd1 vssd1 vccd1 vccd1 _11098_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08146__B1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10039_ _10039_/A _10039_/B vssd1 vssd1 vccd1 vccd1 _10039_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__09894__B1 _07117_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07450__A _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_20 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07250_ _10749_/A vssd1 vssd1 vccd1 vccd1 _10748_/A sky130_fd_sc_hd__inv_6
XFILLER_0_45_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07181_ _11134_/A _11242_/A _07141_/C _07585_/B1 vssd1 vssd1 vccd1 vccd1 _07188_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_54_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11756__A1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11756__B2 _11868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09822_ _09822_/A _11497_/A vssd1 vssd1 vccd1 vccd1 _09828_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10731__A2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10192__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09753_ _11138_/A _09257_/S _09422_/B _06802_/B _09752_/X vssd1 vssd1 vccd1 vccd1
+ _09753_/X sky130_fd_sc_hd__o221a_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout282_A _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06965_ _12642_/A reg1_val[31] _12359_/A vssd1 vssd1 vccd1 vccd1 _06967_/B sky130_fd_sc_hd__and3_4
X_08704_ _08706_/A _08706_/B vssd1 vssd1 vccd1 vccd1 _08704_/Y sky130_fd_sc_hd__nor2_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06896_ _06753_/Y _10672_/A _06896_/C _10291_/A vssd1 vssd1 vccd1 vccd1 _06900_/A
+ sky130_fd_sc_hd__and4bb_1
X_09684_ _09685_/A _09685_/B vssd1 vssd1 vccd1 vccd1 _09684_/Y sky130_fd_sc_hd__nor2_1
X_08635_ _08640_/A _08640_/B vssd1 vssd1 vccd1 vccd1 _08637_/B sky130_fd_sc_hd__or2_1
XFILLER_0_96_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ _08587_/A _08587_/B vssd1 vssd1 vccd1 vccd1 _08568_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout12 fanout13/X vssd1 vssd1 vccd1 vccd1 fanout12/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__07360__A _12224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07517_ _07518_/A _07518_/B vssd1 vssd1 vccd1 vccd1 _07529_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08456__A _08575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout56 _07050_/Y vssd1 vssd1 vccd1 vccd1 fanout56/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout23 _07362_/B vssd1 vssd1 vccd1 vccd1 fanout23/X sky130_fd_sc_hd__buf_6
Xfanout45 fanout46/X vssd1 vssd1 vccd1 vccd1 fanout45/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_64_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout34 _07201_/X vssd1 vssd1 vccd1 vccd1 fanout34/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08497_ _08497_/A _08497_/B vssd1 vssd1 vccd1 vccd1 _08500_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout67 fanout68/X vssd1 vssd1 vccd1 vccd1 _12233_/A sky130_fd_sc_hd__buf_6
Xfanout89 _11284_/A vssd1 vssd1 vccd1 vccd1 _11582_/A sky130_fd_sc_hd__buf_12
Xfanout78 _08289_/B vssd1 vssd1 vccd1 vccd1 fanout78/X sky130_fd_sc_hd__buf_6
XANTENNA__07073__C_N _10243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07448_ _07451_/A _07451_/B vssd1 vssd1 vccd1 vccd1 _07463_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_9_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07379_ _10749_/A _07379_/B vssd1 vssd1 vccd1 vccd1 _07384_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09118_ _09119_/A _09119_/B vssd1 vssd1 vccd1 vccd1 _09118_/X sky130_fd_sc_hd__and2_1
XFILLER_0_103_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10390_ _10390_/A _10390_/B vssd1 vssd1 vccd1 vccd1 _10393_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07415__A2 _09822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09049_ _09936_/A _09049_/B vssd1 vssd1 vccd1 vccd1 _09053_/A sky130_fd_sc_hd__xnor2_2
X_12060_ reg1_val[24] curr_PC[24] vssd1 vssd1 vccd1 vccd1 _12060_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_102_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11011_ _10781_/Y _11229_/A _11010_/Y vssd1 vssd1 vccd1 vccd1 _11011_/X sky130_fd_sc_hd__a21o_1
XANTENNA__11263__A1_N _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10183__B1 _11752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08128__B1 fanout72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12962_ _12880_/B _13225_/B _12878_/X vssd1 vssd1 vccd1 vccd1 _13230_/A sky130_fd_sc_hd__a21o_1
XANTENNA__11132__C1 _09225_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12893_ hold270/X hold50/X vssd1 vssd1 vccd1 vccd1 _13168_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12587__S _12638_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11913_ _09228_/X _09234_/X _11913_/S vssd1 vssd1 vccd1 vccd1 _11913_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09340__A2 _11198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11844_ _11844_/A _11844_/B vssd1 vssd1 vccd1 vccd1 _11848_/A sky130_fd_sc_hd__xnor2_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07270__A _07270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _11775_/A _11775_/B vssd1 vssd1 vccd1 vccd1 _11776_/B sky130_fd_sc_hd__or2_1
XFILLER_0_83_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10726_ _10726_/A _10726_/B vssd1 vssd1 vccd1 vccd1 _10728_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08851__B2 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08851__A1 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10657_ _10415_/A _10415_/B _10539_/A vssd1 vssd1 vccd1 vccd1 _10658_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13376_ _13379_/CLK _13376_/D vssd1 vssd1 vccd1 vccd1 hold275/A sky130_fd_sc_hd__dfxtp_1
X_10588_ _10588_/A _10588_/B vssd1 vssd1 vccd1 vccd1 _10592_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12335__B _12335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07406__A2 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12327_ _06630_/X _09228_/X _12421_/A1 vssd1 vssd1 vccd1 vccd1 _12327_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10136__A _10136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_528 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12258_ _12364_/A _12258_/B _12258_/C vssd1 vssd1 vccd1 vccd1 _12258_/X sky130_fd_sc_hd__or3_1
X_11209_ _11093_/A _12087_/B _11094_/A _11095_/Y vssd1 vssd1 vccd1 vccd1 _11210_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_76_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10713__A2 _07417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12189_ _06883_/X _12188_/X _12404_/S vssd1 vssd1 vccd1 vccd1 _12189_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10174__B1 _11829_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07445__A _10749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06750_ _06815_/A _06723_/A _12702_/B _06749_/X vssd1 vssd1 vccd1 vccd1 _10813_/A
+ sky130_fd_sc_hd__a31o_4
X_06681_ instruction[32] _06716_/B vssd1 vssd1 vccd1 vccd1 _12675_/B sky130_fd_sc_hd__and2_4
XFILLER_0_92_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09660__A _09794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08420_ _08420_/A _08420_/B vssd1 vssd1 vccd1 vccd1 _08421_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_86_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07893__A2 _07959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09095__A1 _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08351_ _08351_/A _08351_/B vssd1 vssd1 vccd1 vccd1 _08405_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_19_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07302_ _10871_/A fanout74/X fanout72/X fanout78/X vssd1 vssd1 vccd1 vccd1 _07303_/B
+ sky130_fd_sc_hd__o22a_1
X_08282_ _08282_/A _08282_/B vssd1 vssd1 vccd1 vccd1 _08689_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_116_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07233_ _07233_/A _07233_/B vssd1 vssd1 vccd1 vccd1 _07233_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_73_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13121__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07164_ _07172_/A _07149_/A _07959_/A _07147_/B _12438_/A vssd1 vssd1 vccd1 vccd1
+ _07166_/B sky130_fd_sc_hd__o311a_2
XFILLER_0_42_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07095_ _07094_/A _06983_/A _06983_/B _07094_/B vssd1 vssd1 vccd1 vccd1 _07097_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout213 _07959_/A vssd1 vssd1 vccd1 vccd1 _09419_/B sky130_fd_sc_hd__clkbuf_4
Xfanout202 _10243_/A vssd1 vssd1 vccd1 vccd1 _09944_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout246 _06958_/A vssd1 vssd1 vccd1 vccd1 _12631_/S sky130_fd_sc_hd__buf_6
Xfanout235 _09423_/X vssd1 vssd1 vccd1 vccd1 _09425_/C sky130_fd_sc_hd__buf_4
Xfanout224 _07166_/A vssd1 vssd1 vccd1 vccd1 _11138_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout268 _06810_/B vssd1 vssd1 vccd1 vccd1 _06783_/A sky130_fd_sc_hd__clkbuf_8
Xfanout279 _13142_/A vssd1 vssd1 vccd1 vccd1 _13147_/A sky130_fd_sc_hd__buf_4
Xfanout257 hold191/X vssd1 vssd1 vccd1 vccd1 _13000_/A2 sky130_fd_sc_hd__clkbuf_8
X_09805_ _11179_/A _09805_/B vssd1 vssd1 vccd1 vccd1 _09807_/B sky130_fd_sc_hd__xnor2_1
X_07997_ _08059_/A _08059_/B _07976_/X vssd1 vssd1 vccd1 vccd1 _08006_/B sky130_fd_sc_hd__a21o_1
X_06948_ instruction[6] instruction[5] vssd1 vssd1 vccd1 vccd1 _09226_/B sky130_fd_sc_hd__or2_4
XFILLER_0_66_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09736_ _09734_/Y _09736_/B vssd1 vssd1 vccd1 vccd1 _09736_/X sky130_fd_sc_hd__and2b_1
XANTENNA__11665__B1 _11584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09667_ _09667_/A _09667_/B vssd1 vssd1 vccd1 vccd1 _09668_/B sky130_fd_sc_hd__xnor2_2
X_06879_ _12795_/A _07147_/B vssd1 vssd1 vccd1 vccd1 _06879_/X sky130_fd_sc_hd__or2_1
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08618_ _08618_/A _08618_/B _08618_/C vssd1 vssd1 vccd1 vccd1 _08630_/A sky130_fd_sc_hd__and3_2
XANTENNA__07333__A1 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07333__B2 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08530__B1 _08576_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12209__A2 _09257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07090__A _10243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09598_ _09743_/B _12144_/A1 _09422_/B _06809_/A _09593_/X vssd1 vssd1 vccd1 vccd1
+ _09598_/X sky130_fd_sc_hd__o221a_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08549_ _08521_/B _08521_/C _08521_/A vssd1 vssd1 vccd1 vccd1 _08549_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09086__A1 _09661_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09086__B2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12090__B1 _12335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11560_ _11558_/Y _11559_/X _11552_/X _11556_/X vssd1 vssd1 vccd1 vccd1 _11560_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07636__A2 _07554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout7_A fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10511_ _10511_/A _10511_/B vssd1 vssd1 vccd1 vccd1 _10514_/A sky130_fd_sc_hd__nor2_1
X_11491_ _11492_/A _11492_/B vssd1 vssd1 vccd1 vccd1 _11493_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_122_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13230_ _13230_/A _13230_/B vssd1 vssd1 vccd1 vccd1 _13230_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__11340__A _11526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10442_ _06770_/B _09422_/B _10437_/Y _06768_/Y _10441_/X vssd1 vssd1 vccd1 vccd1
+ _10442_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_33_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13161_ hold285/X _13209_/A2 _13160_/X _13171_/B2 vssd1 vssd1 vccd1 vccd1 hold286/A
+ sky130_fd_sc_hd__a22o_1
X_10373_ _11179_/A _10373_/B vssd1 vssd1 vccd1 vccd1 _10501_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_32_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12112_ _12110_/Y _12112_/B vssd1 vssd1 vccd1 vccd1 _12300_/B sky130_fd_sc_hd__nand2b_2
X_13092_ _13355_/Q _12805_/A _13250_/B hold116/X _13039_/A vssd1 vssd1 vccd1 vccd1
+ hold117/A sky130_fd_sc_hd__o221a_1
XFILLER_0_103_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12043_ _12043_/A _12043_/B vssd1 vssd1 vccd1 vccd1 _12043_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12145__A1 _06998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12145__B2 _10159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10156__B1 _09225_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07021__B1 _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09480__A _10749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12945_ hold96/X hold264/X vssd1 vssd1 vccd1 vccd1 _13193_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12876_ hold58/X hold282/X vssd1 vssd1 vccd1 vccd1 _12876_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_87_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ _11990_/A1 _11907_/B hold188/A vssd1 vssd1 vccd1 vccd1 _11827_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11234__B _11271_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11758_ _07051_/X fanout43/X fanout41/X _12169_/A vssd1 vssd1 vccd1 vccd1 _11759_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10709_ _10709_/A _10709_/B _10709_/C vssd1 vssd1 vccd1 vccd1 _10710_/B sky130_fd_sc_hd__or3_1
XFILLER_0_83_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08824__A _09922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11689_ _11689_/A _11689_/B vssd1 vssd1 vccd1 vccd1 _11695_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13359_ _13360_/CLK hold8/X vssd1 vssd1 vccd1 vccd1 hold296/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08052__A2 _08112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07920_ _08598_/B fanout76/X fanout72/X _08538_/A1 vssd1 vssd1 vccd1 vccd1 _07921_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07175__A _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10698__B2 _10788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07851_ _08515_/A2 _10595_/A1 fanout72/X _08540_/B vssd1 vssd1 vccd1 vccd1 _07852_/B
+ sky130_fd_sc_hd__o22a_1
X_06802_ _06800_/Y _06802_/B vssd1 vssd1 vccd1 vccd1 _09745_/B sky130_fd_sc_hd__nand2b_1
X_07782_ _07867_/A _07867_/B _07770_/X vssd1 vssd1 vccd1 vccd1 _07802_/B sky130_fd_sc_hd__a21oi_2
X_06733_ _11259_/S _06733_/B vssd1 vssd1 vccd1 vccd1 _11239_/A sky130_fd_sc_hd__nor2_2
X_09521_ _11770_/A _09521_/B vssd1 vssd1 vccd1 vccd1 _09522_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07903__A _10207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06664_ reg1_val[31] _07147_/B vssd1 vssd1 vccd1 vccd1 _06962_/B sky130_fd_sc_hd__xnor2_2
X_09452_ _09453_/B _09452_/B vssd1 vssd1 vccd1 vccd1 _09624_/A sky130_fd_sc_hd__and2b_1
X_06595_ instruction[21] _06944_/B vssd1 vssd1 vccd1 vccd1 _06595_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09383_ _09165_/X _09169_/X _09383_/S vssd1 vssd1 vccd1 vccd1 _09383_/X sky130_fd_sc_hd__mux2_1
X_08403_ _08403_/A _08403_/B _08403_/C vssd1 vssd1 vccd1 vccd1 _08403_/X sky130_fd_sc_hd__and3_1
XANTENNA_fanout245_A _12631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07618__A2 _09943_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08334_ _08334_/A _08392_/A _08392_/B vssd1 vssd1 vccd1 vccd1 _08345_/A sky130_fd_sc_hd__or3_1
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10622__A1 _10476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10622__B2 _08411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08265_ _08265_/A _08265_/B vssd1 vssd1 vccd1 vccd1 _08267_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07216_ _07215_/A _07214_/X _07215_/Y _06983_/A vssd1 vssd1 vccd1 vccd1 _10337_/A
+ sky130_fd_sc_hd__o22a_4
XFILLER_0_61_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08196_ _08263_/A _08263_/B vssd1 vssd1 vccd1 vccd1 _08264_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07147_ _12359_/A _07147_/B _07959_/A vssd1 vssd1 vccd1 vccd1 _07149_/B sky130_fd_sc_hd__and3_2
XANTENNA__08579__B1 _09325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10386__B1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07078_ _07078_/A _07088_/B _07078_/C vssd1 vssd1 vccd1 vccd1 _07080_/B sky130_fd_sc_hd__or3_4
XANTENNA__09791__A2 _10473_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10689__A1 _12421_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout60_A _07033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10991_ _10871_/A _12087_/B _10872_/A _10875_/A vssd1 vssd1 vccd1 vccd1 _10993_/B
+ sky130_fd_sc_hd__o31a_1
X_09719_ _09383_/X _09386_/X _09727_/S vssd1 vssd1 vccd1 vccd1 _09719_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08503__B1 _08561_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_6_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13392_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ reg1_val[18] _12755_/B vssd1 vssd1 vccd1 vccd1 _12732_/A sky130_fd_sc_hd__nand2_2
XANTENNA__10861__B2 _10974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10861__A1 _11093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12661_ _12659_/Y _12661_/B vssd1 vssd1 vccd1 vccd1 _12662_/B sky130_fd_sc_hd__and2b_1
X_11612_ _11612_/A _11612_/B _11612_/C vssd1 vssd1 vccd1 vccd1 _11613_/B sky130_fd_sc_hd__and3_1
XFILLER_0_108_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12592_ _12597_/C _12592_/B vssd1 vssd1 vccd1 vccd1 new_PC[19] sky130_fd_sc_hd__xnor2_4
XANTENNA__07609__A2 _07316_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11543_ reg1_val[18] curr_PC[18] vssd1 vssd1 vccd1 vccd1 _11545_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11474_ _07234_/Y _12158_/B _11473_/Y _11582_/A vssd1 vssd1 vccd1 vccd1 _11591_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_52_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13213_ hold266/A _13212_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13213_/X sky130_fd_sc_hd__mux2_1
X_10425_ _10313_/A _10310_/Y _10312_/B vssd1 vssd1 vccd1 vccd1 _10429_/A sky130_fd_sc_hd__o21a_1
XANTENNA__08034__A2 _08411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13144_ _13144_/A _13144_/B vssd1 vssd1 vccd1 vccd1 _13144_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10356_ _10356_/A _10356_/B vssd1 vssd1 vccd1 vccd1 _10367_/A sky130_fd_sc_hd__xor2_1
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06611__B _06675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13075_ _07230_/B _12826_/B hold134/X vssd1 vssd1 vccd1 vccd1 _13347_/D sky130_fd_sc_hd__a21boi_1
XFILLER_0_57_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10287_ _11893_/A _10287_/B _10287_/C vssd1 vssd1 vccd1 vccd1 _10287_/X sky130_fd_sc_hd__or3_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12026_ _12027_/A _12027_/B _12027_/C vssd1 vssd1 vccd1 vccd1 _12108_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__08819__A _09779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09298__A1 _09298_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09298__B2 _09298_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12928_ hold22/X hold294/A vssd1 vssd1 vccd1 vccd1 _13148_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07848__A2 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12841__A2 _12863_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12859_ _06998_/X _12871_/A2 hold65/X _13249_/A vssd1 vssd1 vccd1 vccd1 _13290_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_3_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08050_ _08051_/A _08051_/B vssd1 vssd1 vccd1 vccd1 _08050_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_113_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07001_ _12642_/A _12644_/A reg1_val[2] reg1_val[3] vssd1 vssd1 vccd1 vccd1 _07083_/C
+ sky130_fd_sc_hd__or4_2
XFILLER_0_12_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12804__A _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08952_ _09944_/A _08952_/B vssd1 vssd1 vccd1 vccd1 _08954_/B sky130_fd_sc_hd__xnor2_1
X_07903_ _10207_/A _07903_/B vssd1 vssd1 vccd1 vccd1 _07968_/A sky130_fd_sc_hd__xnor2_2
X_08883_ _08883_/A _08883_/B vssd1 vssd1 vccd1 vccd1 _08898_/A sky130_fd_sc_hd__xor2_1
X_07834_ _08656_/A _07834_/B _07834_/C vssd1 vssd1 vccd1 vccd1 _07837_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12817__C1 _13147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07765_ _08564_/A _07765_/B vssd1 vssd1 vccd1 vccd1 _07824_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09289__A1 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09289__B2 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06716_ instruction[27] _06716_/B vssd1 vssd1 vccd1 vccd1 _12650_/B sky130_fd_sc_hd__and2_4
XFILLER_0_79_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09504_ _09673_/A _07030_/B _12158_/B _09503_/Y vssd1 vssd1 vccd1 vccd1 _09505_/B
+ sky130_fd_sc_hd__a31o_2
XANTENNA__07839__A2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07696_ _09669_/B2 fanout51/X _09661_/B2 _09301_/A vssd1 vssd1 vccd1 vccd1 _07697_/B
+ sky130_fd_sc_hd__o22a_1
X_06647_ instruction[35] _06675_/B vssd1 vssd1 vccd1 vccd1 _12689_/B sky130_fd_sc_hd__and2_4
XFILLER_0_79_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09435_ _07172_/A _09434_/X _09248_/B vssd1 vssd1 vccd1 vccd1 _09436_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_63_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06578_ instruction[3] vssd1 vssd1 vccd1 vccd1 _06949_/A sky130_fd_sc_hd__inv_2
X_09366_ _09366_/A _09366_/B vssd1 vssd1 vccd1 vccd1 _09368_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_117_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_40 reg2_val[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08317_ _08317_/A _08317_/B vssd1 vssd1 vccd1 vccd1 _08364_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_299 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09297_ _09467_/B _09297_/B vssd1 vssd1 vccd1 vccd1 _09324_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_62_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_51 reg1_val[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08248_ _08575_/A _08248_/B vssd1 vssd1 vccd1 vccd1 _08313_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07472__B1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10359__B1 _07274_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10210_ _10211_/A _10211_/B vssd1 vssd1 vccd1 vccd1 _10212_/A sky130_fd_sc_hd__nor2_1
X_08179_ _08179_/A _08179_/B vssd1 vssd1 vccd1 vccd1 _08182_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_113_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11190_ _11190_/A _11190_/B vssd1 vssd1 vccd1 vccd1 _11193_/A sky130_fd_sc_hd__nor2_1
XANTENNA__09764__A2 _09760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10141_ _09999_/A _09999_/B _10140_/X vssd1 vssd1 vccd1 vccd1 _10143_/A sky130_fd_sc_hd__a21oi_2
X_10072_ _10072_/A fanout8/X vssd1 vssd1 vccd1 vccd1 _10072_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_100_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10974_ _10974_/A _12017_/A vssd1 vssd1 vccd1 vccd1 _10975_/B sky130_fd_sc_hd__nor2_1
XANTENNA__06750__A2 _06723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12823__A2 _13101_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12713_ reg1_val[14] _12714_/B vssd1 vssd1 vccd1 vccd1 _12721_/A sky130_fd_sc_hd__nand2_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12644_ _12644_/A _12645_/B vssd1 vssd1 vccd1 vccd1 _12646_/A sky130_fd_sc_hd__or2_1
XANTENNA__08374__A _08575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12575_ _12639_/A _12575_/B vssd1 vssd1 vccd1 vccd1 _12582_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_38_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11526_ _11526_/A _11618_/A vssd1 vssd1 vccd1 vccd1 _11712_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_4_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06805__A3 _12655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13000__A2 _13000_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11457_ _06719_/X _12420_/A0 _12421_/A1 vssd1 vssd1 vccd1 vccd1 _11457_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11388_ _11389_/A _11389_/B vssd1 vssd1 vccd1 vccd1 _11509_/B sky130_fd_sc_hd__nand2b_1
X_10408_ _10408_/A _10408_/B vssd1 vssd1 vccd1 vccd1 _10409_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_21_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10339_ _12157_/A _10339_/B vssd1 vssd1 vccd1 vccd1 _10341_/B sky130_fd_sc_hd__xnor2_1
X_13127_ _13147_/A hold249/X vssd1 vssd1 vccd1 vccd1 _13366_/D sky130_fd_sc_hd__and2_1
XFILLER_0_0_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ hold145/X _13094_/A2 _13101_/A2 hold98/X _13039_/A vssd1 vssd1 vccd1 vccd1
+ hold146/A sky130_fd_sc_hd__o221a_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12009_ _12009_/A _12009_/B vssd1 vssd1 vccd1 vccd1 _12010_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_84_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08191__A1 _08641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13067__A2 _12826_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08191__B2 _08627_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11078__B2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11078__A1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07550_ _07556_/B _07556_/C _07556_/A vssd1 vssd1 vccd1 vccd1 _07558_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_124_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09220_ _12064_/S _09216_/X _09219_/X _12446_/C1 vssd1 vssd1 vccd1 vccd1 _09220_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07481_ _07604_/A _07481_/B vssd1 vssd1 vccd1 vccd1 _07682_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_124_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09151_ _10049_/A _10321_/A _10321_/B _09150_/X vssd1 vssd1 vccd1 vccd1 _09151_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10589__B1 _07262_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11250__A1 _11820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07454__B1 _10245_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08102_ _08454_/A _08102_/B vssd1 vssd1 vccd1 vccd1 _08108_/A sky130_fd_sc_hd__xnor2_1
X_09082_ _08199_/B fanout84/X _11198_/A fanout33/X vssd1 vssd1 vccd1 vccd1 _09083_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08033_ _08334_/A _08033_/B vssd1 vssd1 vccd1 vccd1 _08036_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout110_A _07237_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09984_ _09984_/A _09984_/B vssd1 vssd1 vccd1 vccd1 _09997_/A sky130_fd_sc_hd__xor2_4
X_08935_ _07554_/B _12823_/A1 _07282_/Y _07175_/A vssd1 vssd1 vccd1 vccd1 _08936_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08866_ _08866_/A _08866_/B vssd1 vssd1 vccd1 vccd1 _08867_/B sky130_fd_sc_hd__xnor2_2
X_07817_ _08706_/A _08706_/B vssd1 vssd1 vccd1 vccd1 _07817_/Y sky130_fd_sc_hd__nand2_1
X_08797_ _08793_/A _08793_/B _08793_/C _08794_/A _08711_/A vssd1 vssd1 vccd1 vccd1
+ _08799_/C sky130_fd_sc_hd__a311o_2
X_07748_ _07748_/A _07748_/B vssd1 vssd1 vccd1 vccd1 _07813_/A sky130_fd_sc_hd__xor2_1
XANTENNA__10816__B2 _10159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07679_ _07679_/A _07679_/B vssd1 vssd1 vccd1 vccd1 _07745_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_109_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12018__B1 _08859_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10690_ hold294/A _10690_/B vssd1 vssd1 vccd1 vccd1 _10810_/B sky130_fd_sc_hd__or2_1
XANTENNA_fanout23_A _07362_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09418_ _09418_/A _09418_/B vssd1 vssd1 vccd1 vccd1 _09418_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12428__B _12428_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09349_ _09350_/A _09350_/B vssd1 vssd1 vccd1 vccd1 _09349_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_105_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12360_ _12359_/A _12358_/X _12359_/Y vssd1 vssd1 vccd1 vccd1 _12360_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10229__A _11844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11311_ _11311_/A _11311_/B vssd1 vssd1 vccd1 vccd1 _11313_/B sky130_fd_sc_hd__and2_1
XFILLER_0_90_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12291_ _12291_/A _12341_/A vssd1 vssd1 vccd1 vccd1 _12292_/C sky130_fd_sc_hd__and2_1
XANTENNA__08641__B _08641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11242_ _11242_/A curr_PC[15] vssd1 vssd1 vccd1 vccd1 _11243_/B sky130_fd_sc_hd__nor2_1
X_11173_ _11174_/A _11174_/B vssd1 vssd1 vccd1 vccd1 _11318_/B sky130_fd_sc_hd__or2_1
XFILLER_0_101_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10124_ _10124_/A _10124_/B vssd1 vssd1 vccd1 vccd1 _10127_/A sky130_fd_sc_hd__or2_2
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10055_ _10053_/X _10055_/B vssd1 vssd1 vccd1 vccd1 _10056_/B sky130_fd_sc_hd__and2b_1
XANTENNA__09472__B _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08369__A _08664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07273__A _11038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07920__B2 _08538_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07920__A1 _08598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10957_ fanout58/X fanout47/X fanout45/X _11868_/A vssd1 vssd1 vccd1 vccd1 _10958_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12627_ _12633_/A _12627_/B vssd1 vssd1 vccd1 vccd1 _12628_/B sky130_fd_sc_hd__nor2_1
XANTENNA__06617__A _06927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10888_ _10888_/A _10888_/B vssd1 vssd1 vccd1 vccd1 _10890_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_73_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12558_ _12567_/A _12558_/B vssd1 vssd1 vccd1 vccd1 _12560_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_80_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11509_ _11509_/A _11509_/B _11509_/C vssd1 vssd1 vccd1 vccd1 _11510_/B sky130_fd_sc_hd__and3_1
Xhold107 hold107/A vssd1 vssd1 vccd1 vccd1 hold107/X sky130_fd_sc_hd__dlygate4sd3_1
X_12489_ _12490_/A _12490_/B _12490_/C vssd1 vssd1 vccd1 vccd1 _12497_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_81_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold129 hold129/A vssd1 vssd1 vccd1 vccd1 hold129/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 hold118/A vssd1 vssd1 vccd1 vccd1 hold118/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ _07078_/A _07087_/A _07097_/A _07094_/A vssd1 vssd1 vccd1 vccd1 _06983_/C
+ sky130_fd_sc_hd__and4_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11299__B2 _11779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11299__A1 _07013_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10602__A _11393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08720_ _08720_/A _08720_/B vssd1 vssd1 vccd1 vccd1 _10010_/B sky130_fd_sc_hd__nor2_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09900__A2 _12446_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08651_ _08665_/A _08665_/B vssd1 vssd1 vccd1 vccd1 _08654_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07911__A1 _09669_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07911__B2 _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07602_ _07602_/A _07602_/B vssd1 vssd1 vccd1 vccd1 _07644_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_44_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08582_ _08583_/A _08582_/B _08582_/C vssd1 vssd1 vccd1 vccd1 _08596_/A sky130_fd_sc_hd__nand3_2
XANTENNA__12529__A _12689_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07533_ _07533_/A _07533_/B _07533_/C vssd1 vssd1 vccd1 vccd1 _07537_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_119_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07464_ _07466_/A _07464_/B vssd1 vssd1 vccd1 vccd1 _07563_/B sky130_fd_sc_hd__or2_1
XFILLER_0_9_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09203_ reg1_val[13] reg1_val[18] _09211_/S vssd1 vssd1 vccd1 vccd1 _09203_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10049__A _10049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07395_ _07400_/B _07395_/B vssd1 vssd1 vccd1 vccd1 _07434_/A sky130_fd_sc_hd__nor2_1
X_09134_ _09012_/A _09012_/B _09013_/X vssd1 vssd1 vccd1 vccd1 _09136_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_17_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12420__A0 _12420_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09065_ _09066_/A _09066_/B _09066_/C vssd1 vssd1 vccd1 vccd1 _09278_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08016_ _08016_/A _08016_/B vssd1 vssd1 vccd1 vccd1 _08073_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_102_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09967_ _09777_/Y _09780_/B _09776_/A vssd1 vssd1 vccd1 vccd1 _09980_/A sky130_fd_sc_hd__a21o_1
X_08918_ _07676_/A _07676_/B _08708_/A _08708_/B vssd1 vssd1 vccd1 vccd1 _08918_/X
+ sky130_fd_sc_hd__o22a_1
X_09898_ _09896_/Y _09898_/B vssd1 vssd1 vccd1 vccd1 _09899_/B sky130_fd_sc_hd__nand2b_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08849_ _08850_/A _08850_/B vssd1 vssd1 vccd1 vccd1 _08849_/X sky130_fd_sc_hd__and2b_1
XANTENNA__07902__A1 _10221_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07902__B2 _09770_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11860_ _11860_/A _11860_/B vssd1 vssd1 vccd1 vccd1 _11861_/B sky130_fd_sc_hd__nand2_1
X_11791_ _11881_/A _11791_/B vssd1 vssd1 vccd1 vccd1 _11793_/C sky130_fd_sc_hd__and2_1
X_10811_ _12271_/A1 _10924_/B hold288/A vssd1 vssd1 vccd1 vccd1 _10811_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10742_ _10742_/A _10742_/B vssd1 vssd1 vccd1 vccd1 _10758_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12158__B _12158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12006__A3 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10673_ _10672_/A _10672_/B _11637_/A vssd1 vssd1 vccd1 vccd1 _10673_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_47_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13392_ _13392_/CLK _13392_/D vssd1 vssd1 vccd1 vccd1 hold175/A sky130_fd_sc_hd__dfxtp_1
X_12412_ _12412_/A _12412_/B vssd1 vssd1 vccd1 vccd1 _12412_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12343_ _07316_/Y _11946_/C _12287_/A _12285_/A vssd1 vssd1 vccd1 vccd1 _12345_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08091__B1 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12274_ _07049_/A _09257_/S _09422_/B _06645_/B _12631_/S vssd1 vssd1 vccd1 vccd1
+ _12274_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_120_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11225_ _11223_/Y _11225_/B vssd1 vssd1 vccd1 vccd1 _11433_/A sky130_fd_sc_hd__nand2b_4
XFILLER_0_50_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11156_ _09222_/Y _11141_/B _11155_/Y _10159_/A _11153_/X vssd1 vssd1 vccd1 vccd1
+ _11156_/X sky130_fd_sc_hd__o221a_1
X_11087_ _11087_/A _11087_/B vssd1 vssd1 vccd1 vccd1 _11088_/B sky130_fd_sc_hd__xnor2_1
X_10107_ _07171_/A _07269_/Y _07274_/Y fanout38/X vssd1 vssd1 vccd1 vccd1 _10108_/B
+ sky130_fd_sc_hd__a22o_1
X_10038_ _10036_/Y _10038_/B vssd1 vssd1 vccd1 vccd1 _10039_/B sky130_fd_sc_hd__and2b_1
XANTENNA__08146__A1 _08576_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08146__B2 _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11150__A0 _12420_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09894__B2 _12422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11989_ hold219/A _11989_/B vssd1 vssd1 vccd1 vccd1 _12065_/B sky130_fd_sc_hd__or2_1
XFILLER_0_58_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07180_ _07242_/A vssd1 vssd1 vccd1 vccd1 _07180_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08562__A _08575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11756__A2 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10964__B1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10716__B1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10192__A1 _11406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09821_ _09821_/A _09821_/B vssd1 vssd1 vccd1 vccd1 _09830_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__10192__B2 _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ hold256/A _09750_/X _09751_/Y vssd1 vssd1 vccd1 vccd1 _09752_/X sky130_fd_sc_hd__a21o_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06964_ reg1_val[31] _12359_/A vssd1 vssd1 vccd1 vccd1 _06964_/X sky130_fd_sc_hd__and2_1
X_08703_ _08711_/A _08711_/B _08805_/A _08701_/X vssd1 vssd1 vccd1 vccd1 _08802_/A
+ sky130_fd_sc_hd__o31ai_4
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout275_A _13162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06895_ _11636_/A _11541_/A _11449_/A vssd1 vssd1 vccd1 vccd1 _06901_/B sky130_fd_sc_hd__and3_1
X_09683_ _09683_/A _09683_/B vssd1 vssd1 vccd1 vccd1 _09685_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08634_ _08656_/A _08634_/B vssd1 vssd1 vccd1 vccd1 _08640_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08565_ _08594_/A _08570_/B _08558_/X vssd1 vssd1 vccd1 vccd1 _08587_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_119_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout13 _08860_/Y vssd1 vssd1 vccd1 vccd1 fanout13/X sky130_fd_sc_hd__buf_4
XFILLER_0_76_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07516_ _07705_/A _07705_/B _07512_/X vssd1 vssd1 vccd1 vccd1 _07518_/B sky130_fd_sc_hd__o21ai_1
Xfanout24 _07361_/Y vssd1 vssd1 vccd1 vccd1 _07362_/B sky130_fd_sc_hd__clkbuf_8
Xfanout46 _07137_/X vssd1 vssd1 vccd1 vccd1 fanout46/X sky130_fd_sc_hd__buf_6
X_08496_ _08496_/A _08496_/B vssd1 vssd1 vccd1 vccd1 _08521_/A sky130_fd_sc_hd__xor2_1
Xfanout35 _07192_/Y vssd1 vssd1 vccd1 vccd1 _08199_/B sky130_fd_sc_hd__buf_8
XFILLER_0_9_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout68 _06991_/Y vssd1 vssd1 vccd1 vccd1 fanout68/X sky130_fd_sc_hd__buf_8
XFILLER_0_92_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout79 _07268_/Y vssd1 vssd1 vccd1 vccd1 _08289_/B sky130_fd_sc_hd__buf_8
Xfanout57 _07035_/X vssd1 vssd1 vccd1 vccd1 fanout57/X sky130_fd_sc_hd__buf_8
X_07447_ _09667_/A _07447_/B vssd1 vssd1 vccd1 vccd1 _07451_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07378_ _11309_/A _10473_/B2 _10240_/A fanout80/X vssd1 vssd1 vccd1 vccd1 _07379_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_122_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09117_ _09834_/A _09117_/B vssd1 vssd1 vccd1 vccd1 _09119_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_115_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09048_ _09822_/A _07362_/B fanout16/X _09677_/A vssd1 vssd1 vccd1 vccd1 _09049_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_60_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout90_A _09922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11010_ _10776_/X _10896_/X _10898_/B vssd1 vssd1 vccd1 vccd1 _11010_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__10242__A _10749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08128__B2 _08649_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08128__A1 _08657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12961_ _13220_/A _13221_/A _13220_/B vssd1 vssd1 vccd1 vccd1 _13225_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__09876__A1 _12404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11912_ hold266/A _12271_/A1 _11992_/B _12376_/C1 vssd1 vssd1 vccd1 vccd1 _11912_/X
+ sky130_fd_sc_hd__a31o_1
X_12892_ hold272/X hold20/X vssd1 vssd1 vccd1 vccd1 _13173_/A sky130_fd_sc_hd__nand2b_1
X_11843_ _12233_/A fanout23/X fanout15/X _12087_/A vssd1 vssd1 vccd1 vccd1 _11844_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07551__A _07959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12169__A _12169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _11773_/B _11774_/B vssd1 vssd1 vccd1 vccd1 _11775_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_83_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10725_ _10725_/A _12428_/B vssd1 vssd1 vccd1 vccd1 _10726_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08851__A2 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10656_ _10656_/A _10656_/B vssd1 vssd1 vccd1 vccd1 _10900_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_36_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08382__A _10207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13375_ _13379_/CLK _13375_/D vssd1 vssd1 vccd1 vccd1 hold272/A sky130_fd_sc_hd__dfxtp_1
X_10587_ _10587_/A vssd1 vssd1 vccd1 vccd1 _10588_/B sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_4_8_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12326_ hold287/A _12449_/B1 _12374_/B _12325_/Y _12376_/C1 vssd1 vssd1 vccd1 vccd1
+ _12326_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_50_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10136__B _10136_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12257_ _12364_/A _12258_/B _12258_/C vssd1 vssd1 vccd1 vccd1 _12257_/Y sky130_fd_sc_hd__o21ai_1
X_11208_ _11088_/A _11088_/B _11086_/X vssd1 vssd1 vccd1 vccd1 _11212_/A sky130_fd_sc_hd__a21o_1
X_12188_ _06672_/A _12124_/X _12143_/S vssd1 vssd1 vccd1 vccd1 _12188_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07726__A _09836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11139_ _11246_/S _10161_/X _11138_/X _11029_/S vssd1 vssd1 vccd1 vccd1 _11139_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10152__A _10788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09941__A _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06680_ _11995_/A _06680_/B vssd1 vssd1 vccd1 vccd1 _06700_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12320__C1 _06946_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10298__S _11138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08350_ _08350_/A _08350_/B vssd1 vssd1 vccd1 vccd1 _08351_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_74_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09095__A2 _12158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07301_ _10749_/A _07301_/B vssd1 vssd1 vccd1 vccd1 _07306_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08281_ _08779_/B _08769_/A vssd1 vssd1 vccd1 vccd1 _08281_/X sky130_fd_sc_hd__or2_1
X_07232_ _07233_/A _07233_/B vssd1 vssd1 vccd1 vccd1 _07232_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_61_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07163_ _07149_/A _07959_/A _12438_/A _07147_/B vssd1 vssd1 vccd1 vccd1 _07173_/B
+ sky130_fd_sc_hd__o211a_4
XFILLER_0_41_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07094_ _07094_/A _07094_/B vssd1 vssd1 vccd1 vccd1 _07094_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12542__A _12702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout214 _06817_/X vssd1 vssd1 vccd1 vccd1 _07959_/A sky130_fd_sc_hd__clkbuf_8
Xfanout203 _07063_/Y vssd1 vssd1 vccd1 vccd1 _10243_/A sky130_fd_sc_hd__buf_6
Xfanout247 _06911_/Y vssd1 vssd1 vccd1 vccd1 _06958_/A sky130_fd_sc_hd__buf_6
Xfanout236 _09226_/X vssd1 vssd1 vccd1 vccd1 _11637_/A sky130_fd_sc_hd__clkbuf_8
X_09804_ fanout63/X fanout78/X fanout74/X fanout62/X vssd1 vssd1 vccd1 vccd1 _09805_/B
+ sky130_fd_sc_hd__o22a_1
Xfanout269 _06607_/X vssd1 vssd1 vccd1 vccd1 _06810_/B sky130_fd_sc_hd__buf_4
Xfanout258 _13248_/A2 vssd1 vssd1 vccd1 vccd1 _13171_/B2 sky130_fd_sc_hd__buf_4
XANTENNA__10062__A _11179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07996_ _07996_/A _07996_/B vssd1 vssd1 vccd1 vccd1 _08059_/B sky130_fd_sc_hd__xnor2_2
X_06947_ instruction[6] instruction[5] _09234_/C vssd1 vssd1 vccd1 vccd1 _09242_/B
+ sky130_fd_sc_hd__or3_4
X_09735_ reg1_val[3] curr_PC[3] vssd1 vssd1 vccd1 vccd1 _09736_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11665__A1 _07218_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09666_ fanout61/X _07268_/Y fanout75/X fanout53/X vssd1 vssd1 vccd1 vccd1 _09667_/B
+ sky130_fd_sc_hd__o22a_1
X_06878_ _12406_/A _06877_/Y _06865_/X vssd1 vssd1 vccd1 vccd1 _06878_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08617_ _09673_/A _08617_/B vssd1 vssd1 vccd1 vccd1 _08618_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__07333__A2 _09943_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08530__B2 _08627_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08530__A1 _08641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ _12064_/S _09581_/Y _09596_/Y _09242_/B vssd1 vssd1 vccd1 vccd1 _09597_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08548_ _08521_/B _08521_/C _08521_/A vssd1 vssd1 vccd1 vccd1 _08683_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__09086__A2 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12090__B2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12090__A1 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08294__B1 _08501_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08479_ _08511_/A vssd1 vssd1 vccd1 vccd1 _08479_/Y sky130_fd_sc_hd__inv_2
X_11490_ _11490_/A _11490_/B vssd1 vssd1 vccd1 vccd1 _11492_/B sky130_fd_sc_hd__xor2_1
X_10510_ _10510_/A _10510_/B vssd1 vssd1 vccd1 vccd1 _10511_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_64_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11340__B _11340_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12378__C1 _12422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10441_ _07215_/A _06960_/X _10439_/Y _10440_/X vssd1 vssd1 vccd1 vccd1 _10441_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13160_ hold288/A _13159_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13160_/X sky130_fd_sc_hd__mux2_1
X_10372_ _12233_/A _08289_/B fanout74/X fanout65/X vssd1 vssd1 vccd1 vccd1 _10373_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_60_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12111_ _12111_/A _12111_/B _12111_/C vssd1 vssd1 vccd1 vccd1 _12112_/B sky130_fd_sc_hd__nand3_1
XANTENNA__10671__S _12054_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13091_ _07155_/C _13101_/B2 hold14/X vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__o21a_1
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12042_ _12042_/A _12113_/A vssd1 vssd1 vccd1 vccd1 _12043_/B sky130_fd_sc_hd__nor2_2
XANTENNA__12145__A2 _09257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold290 hold290/A vssd1 vssd1 vccd1 vccd1 hold290/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07021__A1 _09669_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07021__B2 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12944_ _13188_/B _13189_/A _12888_/X vssd1 vssd1 vccd1 vccd1 _13194_/A sky130_fd_sc_hd__a21o_1
XANTENNA__11656__A1 _09238_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07281__A _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12875_ hold287/A hold28/X vssd1 vssd1 vccd1 vccd1 _13238_/A sky130_fd_sc_hd__nand2b_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _13317_/Q _11826_/B vssd1 vssd1 vccd1 vccd1 _11907_/B sky130_fd_sc_hd__or2_1
X_11757_ _12335_/B _11757_/B vssd1 vssd1 vccd1 vccd1 _11761_/B sky130_fd_sc_hd__xnor2_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12081__A1 _12631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13222__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10708_ _10709_/A _10709_/B _10709_/C vssd1 vssd1 vccd1 vccd1 _10882_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11688_ _11692_/B _11587_/B _11594_/B _11595_/B _11595_/A vssd1 vssd1 vccd1 vccd1
+ _11701_/A sky130_fd_sc_hd__a32oi_4
XFILLER_0_83_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12369__C1 _09242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10639_ _10519_/A _10519_/C _10519_/B vssd1 vssd1 vccd1 vccd1 _10649_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_11_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12384__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13358_ _13358_/CLK _13358_/D vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09936__A _09936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12309_ _12399_/A _12307_/X _12308_/Y vssd1 vssd1 vccd1 vccd1 _12309_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07260__A1 _07270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13289_ _13379_/CLK _13289_/D vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07850_ _07850_/A _07850_/B vssd1 vssd1 vccd1 vccd1 _07853_/B sky130_fd_sc_hd__xor2_1
X_06801_ reg1_val[3] _07165_/A vssd1 vssd1 vccd1 vccd1 _06802_/B sky130_fd_sc_hd__nand2_1
X_07781_ _07781_/A _07781_/B vssd1 vssd1 vccd1 vccd1 _07867_/B sky130_fd_sc_hd__xnor2_2
X_06732_ _11242_/A _07262_/A vssd1 vssd1 vccd1 vccd1 _06733_/B sky130_fd_sc_hd__nor2_1
X_09520_ fanout32/X _07269_/Y _07274_/Y fanout29/X vssd1 vssd1 vccd1 vccd1 _09521_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06663_ _12795_/A _07147_/B vssd1 vssd1 vccd1 vccd1 _06963_/B sky130_fd_sc_hd__xnor2_2
X_09451_ _09922_/A _09451_/B vssd1 vssd1 vccd1 vccd1 _09452_/B sky130_fd_sc_hd__xor2_1
X_06594_ instruction[13] _06590_/X _06593_/X _06716_/B vssd1 vssd1 vccd1 vccd1 reg1_idx[2]
+ sky130_fd_sc_hd__o211a_4
X_09382_ _09162_/X _09164_/X _09383_/S vssd1 vssd1 vccd1 vccd1 _09382_/X sky130_fd_sc_hd__mux2_1
X_08402_ _08402_/A _08402_/B vssd1 vssd1 vccd1 vccd1 _08403_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__12072__A1 _11554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08333_ _08564_/A _08333_/B vssd1 vssd1 vccd1 vccd1 _08392_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11441__A _11840_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout238_A _08502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08264_ _08264_/A _08264_/B vssd1 vssd1 vccd1 vccd1 _08266_/B sky130_fd_sc_hd__nor2_1
XANTENNA_fanout140_A _07172_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10622__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07215_ _07215_/A _07215_/B vssd1 vssd1 vccd1 vccd1 _07215_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_6_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08195_ _08580_/A _08195_/B vssd1 vssd1 vccd1 vccd1 _08263_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10386__A1 _11764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07146_ reg1_val[27] _07146_/B vssd1 vssd1 vccd1 vccd1 _07146_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_42_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08579__B2 _09943_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08579__A1 _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11583__B1 _08974_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10386__B2 _11592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07077_ _07088_/B _07078_/C _07078_/A vssd1 vssd1 vccd1 vccd1 _07080_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_100_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08200__A0 _10092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09718_ _09380_/X _09382_/X _09725_/S vssd1 vssd1 vccd1 vccd1 _09718_/X sky130_fd_sc_hd__mux2_1
X_07979_ _08540_/B _10338_/B2 _08457_/A2 _08515_/A2 vssd1 vssd1 vccd1 vccd1 _07980_/B
+ sky130_fd_sc_hd__o22a_1
X_10990_ _10990_/A _10990_/B vssd1 vssd1 vccd1 vccd1 _10993_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_97_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout53_A _07072_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08503__B2 _08627_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08503__A1 _08641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09649_ _07608_/A _07608_/B _09943_/B2 vssd1 vssd1 vccd1 vccd1 _09652_/B sky130_fd_sc_hd__a21o_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10861__A2 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ reg1_val[4] _12660_/B vssd1 vssd1 vccd1 vccd1 _12661_/B sky130_fd_sc_hd__nand2_1
X_11611_ _11612_/A _11612_/B _11612_/C vssd1 vssd1 vccd1 vccd1 _11613_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__06667__A2_N _06766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12591_ _12598_/A _12591_/B vssd1 vssd1 vccd1 vccd1 _12592_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_108_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08806__A2 _08799_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11542_ _11541_/A _11541_/B _09225_/Y vssd1 vssd1 vccd1 vccd1 _11542_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_80_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13012__B1 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11473_ _11473_/A _12158_/B vssd1 vssd1 vccd1 vccd1 _11473_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13212_ _13212_/A _13212_/B vssd1 vssd1 vccd1 vccd1 _13212_/Y sky130_fd_sc_hd__xnor2_1
X_10424_ _10423_/A _10423_/B _10423_/Y _11637_/A vssd1 vssd1 vccd1 vccd1 _10424_/X
+ sky130_fd_sc_hd__a211o_1
X_13143_ _13143_/A _13143_/B vssd1 vssd1 vccd1 vccd1 _13144_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_60_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10355_ _10355_/A _10355_/B vssd1 vssd1 vccd1 vccd1 _10356_/B sky130_fd_sc_hd__xnor2_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07276__A _09667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13074_ hold100/X _12805_/A _13250_/B hold133/X _13142_/A vssd1 vssd1 vccd1 vccd1
+ hold134/A sky130_fd_sc_hd__o221a_1
X_10286_ _11893_/A _10287_/B _10287_/C vssd1 vssd1 vccd1 vccd1 _10286_/Y sky130_fd_sc_hd__o21ai_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12025_ _12101_/B _12025_/B vssd1 vssd1 vccd1 vccd1 _12027_/C sky130_fd_sc_hd__nor2_1
XANTENNA__13217__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11526__A _11526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09298__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12927_ _13143_/A _13144_/A _13143_/B vssd1 vssd1 vccd1 vccd1 _13149_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__10301__A1 _11990_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12858_ hold64/X _12862_/B vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__or2_1
XFILLER_0_29_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11809_ _11809_/A _11809_/B vssd1 vssd1 vccd1 vccd1 _11810_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_8_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12789_ reg1_val[30] _12790_/B vssd1 vssd1 vccd1 vccd1 _12789_/X sky130_fd_sc_hd__and2_1
XFILLER_0_44_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07000_ _09672_/A _07000_/B vssd1 vssd1 vccd1 vccd1 _07041_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_12_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11565__B1 _11752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12092__A _12093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08951_ fanout65/X _07068_/Y _09650_/A fanout59/X vssd1 vssd1 vccd1 vccd1 _08952_/B
+ sky130_fd_sc_hd__o22a_1
X_07902_ _10221_/B2 _08411_/B _10476_/A _09770_/B2 vssd1 vssd1 vccd1 vccd1 _07903_/B
+ sky130_fd_sc_hd__o22a_1
X_08882_ _08882_/A _08882_/B vssd1 vssd1 vccd1 vccd1 _08883_/B sky130_fd_sc_hd__xnor2_1
X_07833_ _07834_/B _07834_/C _08656_/A vssd1 vssd1 vccd1 vccd1 _07837_/A sky130_fd_sc_hd__o21a_1
XANTENNA_fanout188_A _12803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07764_ _08540_/B fanout76/X fanout72/X _08515_/A2 vssd1 vssd1 vccd1 vccd1 _07765_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09289__A2 _10473_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06715_ _11553_/S _06715_/B vssd1 vssd1 vccd1 vccd1 _11541_/A sky130_fd_sc_hd__or2_2
X_09503_ _07038_/X _12158_/B _09673_/A vssd1 vssd1 vccd1 vccd1 _09503_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07695_ _09672_/A _07695_/B vssd1 vssd1 vccd1 vccd1 _07701_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06646_ _12406_/A _06874_/A vssd1 vssd1 vccd1 vccd1 _06673_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_78_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09434_ _09197_/X _09250_/B _09725_/S vssd1 vssd1 vccd1 vccd1 _09434_/X sky130_fd_sc_hd__mux2_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06577_ _06577_/A vssd1 vssd1 vccd1 vccd1 _06577_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09365_ _09366_/B _09366_/A vssd1 vssd1 vccd1 vccd1 _09365_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_117_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_30 reg2_val[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_41 _07097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08316_ _08316_/A _08316_/B vssd1 vssd1 vccd1 vccd1 _08364_/A sky130_fd_sc_hd__xnor2_2
X_09296_ _09295_/B _09296_/B vssd1 vssd1 vccd1 vccd1 _09297_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_52 reg1_val[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08247_ _08649_/A2 _10595_/A1 fanout72/X _08657_/B vssd1 vssd1 vccd1 vccd1 _08248_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07472__B2 _07134_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07472__A1 _07121_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09749__B1 _12205_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10359__B2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10359__A1 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12714__B _12714_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08178_ _08174_/A _08174_/B _08171_/X vssd1 vssd1 vccd1 vccd1 _08182_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07129_ _07129_/A _07129_/B _07129_/C _07129_/D vssd1 vssd1 vccd1 vccd1 _07136_/B
+ sky130_fd_sc_hd__or4_2
XANTENNA__07096__A _07097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10140_ _09862_/A _09862_/B _09999_/A _09999_/B vssd1 vssd1 vccd1 vccd1 _10140_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10071_ _10246_/A _10071_/B vssd1 vssd1 vccd1 vccd1 _10075_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09921__B1 _07274_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10973_ _10973_/A _10973_/B vssd1 vssd1 vccd1 vccd1 _10975_/A sky130_fd_sc_hd__nor2_1
XANTENNA__06750__A3 _12702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12712_ _12717_/B _12712_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[13] sky130_fd_sc_hd__and2_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07160__B1 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12643_ _12647_/A _12643_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[0] sky130_fd_sc_hd__and2_4
XFILLER_0_26_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12574_ reg1_val[17] curr_PC[17] _12638_/S vssd1 vssd1 vccd1 vccd1 _12575_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_38_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11525_ _11523_/Y _11525_/B vssd1 vssd1 vccd1 vccd1 _11711_/A sky130_fd_sc_hd__nand2b_4
XFILLER_0_92_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11456_ _12444_/B _11454_/Y _11455_/Y _09242_/B vssd1 vssd1 vccd1 vccd1 _11456_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08390__A _08564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11387_ _11387_/A _11387_/B vssd1 vssd1 vccd1 vccd1 _11389_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_104_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11020__S _11813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10407_ _10408_/A _10408_/B vssd1 vssd1 vccd1 vccd1 _10407_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_68_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10338_ _10595_/A1 fanout23/X fanout15/X _10338_/B2 vssd1 vssd1 vccd1 vccd1 _10339_/B
+ sky130_fd_sc_hd__o22a_1
X_13126_ hold248/X _13254_/A2 _13125_/X _06577_/A vssd1 vssd1 vccd1 vccd1 hold249/A
+ sky130_fd_sc_hd__a22o_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _10246_/A _12826_/B hold151/X vssd1 vssd1 vccd1 vccd1 _13338_/D sky130_fd_sc_hd__a21boi_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12008_ _07170_/A _12007_/Y _12006_/X vssd1 vssd1 vccd1 vccd1 _12084_/B sky130_fd_sc_hd__a21o_2
X_10269_ _10270_/A _10270_/B vssd1 vssd1 vccd1 vccd1 _10413_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08191__A2 _10595_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11078__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07480_ fanout63/X _09298_/B2 _09298_/A1 fanout61/X vssd1 vssd1 vccd1 vccd1 _07481_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_124_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12087__A _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10589__A1 _07417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09150_ _09234_/C _09239_/B vssd1 vssd1 vccd1 vccd1 _09150_/X sky130_fd_sc_hd__or2_4
XFILLER_0_71_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10589__B2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07454__A1 _10245_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07454__B2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08101_ _10221_/B2 _08484_/B _09479_/B1 _09770_/B2 vssd1 vssd1 vccd1 vccd1 _08102_/B
+ sky130_fd_sc_hd__o22a_1
X_09081_ _10623_/A _09081_/B vssd1 vssd1 vccd1 vccd1 _09085_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08032_ _08561_/A2 _08289_/B fanout75/X _08561_/B1 vssd1 vssd1 vccd1 vccd1 _08033_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06813__A _12644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09983_ _09981_/Y _09983_/B vssd1 vssd1 vccd1 vccd1 _09984_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_3_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08934_ _08934_/A _08934_/B vssd1 vssd1 vccd1 vccd1 _08937_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12550__A _12708_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08865_ _08866_/A _08866_/B vssd1 vssd1 vccd1 vccd1 _08865_/X sky130_fd_sc_hd__or2_1
XFILLER_0_79_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07816_ _07816_/A _07816_/B vssd1 vssd1 vccd1 vccd1 _08706_/B sky130_fd_sc_hd__xor2_4
X_08796_ _07950_/B _08012_/Y _07948_/X vssd1 vssd1 vccd1 vccd1 _08799_/B sky130_fd_sc_hd__a21o_1
X_07747_ _08708_/A _08708_/B vssd1 vssd1 vccd1 vccd1 _07747_/Y sky130_fd_sc_hd__nand2_1
X_07678_ _07678_/A _07678_/B vssd1 vssd1 vccd1 vccd1 _07745_/A sky130_fd_sc_hd__xor2_4
XANTENNA__08475__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12018__B2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12018__A1 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06629_ _06627_/Y _06724_/B1 _06766_/B reg2_val[28] vssd1 vssd1 vccd1 vccd1 _08973_/B
+ sky130_fd_sc_hd__a2bb2o_4
X_09417_ hold301/A hold293/A _11538_/A _12205_/B1 _09416_/Y vssd1 vssd1 vccd1 vccd1
+ _09429_/B sky130_fd_sc_hd__a311o_1
X_09348_ _09109_/A _09109_/B _09107_/Y vssd1 vssd1 vccd1 vccd1 _09350_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_124_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08642__A0 _09302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11310_ _11309_/A _12017_/A _11309_/C vssd1 vssd1 vccd1 vccd1 _11311_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06799__A3 _12660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09279_ _09279_/A _09279_/B vssd1 vssd1 vccd1 vccd1 _09280_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_105_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06723__A _06723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12290_ _12291_/A _12341_/A vssd1 vssd1 vccd1 vccd1 _12346_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12444__B _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11241_ _11242_/A curr_PC[15] vssd1 vssd1 vccd1 vccd1 _11243_/A sky130_fd_sc_hd__and2_1
XFILLER_0_31_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11172_ _12336_/A _11172_/B vssd1 vssd1 vccd1 vccd1 _11174_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10123_ _09925_/A _09925_/B _09928_/A vssd1 vssd1 vccd1 vccd1 _10128_/A sky130_fd_sc_hd__a21o_2
X_10054_ _07282_/Y _11946_/C _09956_/Y _09958_/Y vssd1 vssd1 vccd1 vccd1 _10055_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__07554__A _07959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07920__A2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10956_ _10956_/A _10956_/B vssd1 vssd1 vccd1 vccd1 _10967_/B sky130_fd_sc_hd__or2_1
XFILLER_0_85_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10807__A2 _11990_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10887_ _10766_/A _10766_/B _10764_/Y vssd1 vssd1 vccd1 vccd1 _10888_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_85_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12626_ _12639_/A _12627_/B vssd1 vssd1 vccd1 vccd1 _12628_/A sky130_fd_sc_hd__and2_1
XANTENNA__11768__B1 _12335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12557_ _12714_/B _12557_/B vssd1 vssd1 vccd1 vccd1 _12558_/B sky130_fd_sc_hd__or2_1
XFILLER_0_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08633__B1 _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11508_ _11509_/A _11509_/B _11509_/C vssd1 vssd1 vccd1 vccd1 _11510_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__10991__A1 _10871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12488_ _12497_/A _12488_/B vssd1 vssd1 vccd1 vccd1 _12490_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10440__B1 _12416_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold108 hold108/A vssd1 vssd1 vccd1 vccd1 hold108/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12980__A2 _13000_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11439_ _10548_/B _11009_/Y _11435_/Y _11438_/Y vssd1 vssd1 vccd1 vccd1 _11440_/B
+ sky130_fd_sc_hd__o31ai_4
Xhold119 hold119/A vssd1 vssd1 vccd1 vccd1 hold119/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09944__A _09944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11535__A3 _11567_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13109_ _13147_/A hold236/X vssd1 vssd1 vccd1 vccd1 _13362_/D sky130_fd_sc_hd__and2_1
XFILLER_0_0_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06980_ _07097_/A _07094_/A vssd1 vssd1 vccd1 vccd1 _06980_/X sky130_fd_sc_hd__and2_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11299__A2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09900__A3 _09899_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08650_ _08658_/A _08650_/B vssd1 vssd1 vccd1 vccd1 _08665_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07911__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07601_ _07601_/A _07601_/B _07601_/C vssd1 vssd1 vccd1 vccd1 _07602_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08581_ _08608_/A _08608_/B _08578_/C vssd1 vssd1 vccd1 vccd1 _08582_/C sky130_fd_sc_hd__a21o_1
XANTENNA__11456__C1 _09242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08295__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07532_ _07490_/A _07490_/B _07489_/X vssd1 vssd1 vccd1 vccd1 _07533_/C sky130_fd_sc_hd__o21bai_1
XFILLER_0_119_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11433__B _11526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07463_ _07463_/A _07463_/B _07531_/A vssd1 vssd1 vccd1 vccd1 _07464_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_119_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09202_ _09200_/X _09201_/X _09403_/S vssd1 vssd1 vccd1 vccd1 _09202_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07394_ _07394_/A _07394_/B vssd1 vssd1 vccd1 vccd1 _07395_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_8_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09133_ _09001_/A _09001_/B _08999_/Y vssd1 vssd1 vccd1 vccd1 _09136_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12420__A1 _09422_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13140__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout220_A _07172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09064_ _08964_/X _09064_/B vssd1 vssd1 vccd1 vccd1 _09069_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_102_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08015_ _08015_/A _08015_/B vssd1 vssd1 vccd1 vccd1 _08073_/A sky130_fd_sc_hd__and2_1
XFILLER_0_102_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09966_ _10124_/B _09966_/B vssd1 vssd1 vccd1 vccd1 _09982_/A sky130_fd_sc_hd__or2_1
X_09897_ reg1_val[4] curr_PC[4] vssd1 vssd1 vccd1 vccd1 _09898_/B sky130_fd_sc_hd__nand2_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08917_ _08917_/A _08917_/B vssd1 vssd1 vccd1 vccd1 _09549_/A sky130_fd_sc_hd__xnor2_4
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08848_ _10092_/A _08848_/B vssd1 vssd1 vccd1 vccd1 _08850_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07902__A2 _08411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08779_ _08779_/A _08779_/B vssd1 vssd1 vccd1 vccd1 _08779_/X sky130_fd_sc_hd__or2_1
X_11790_ _11790_/A _11790_/B vssd1 vssd1 vccd1 vccd1 _11791_/B sky130_fd_sc_hd__or2_1
X_10810_ hold279/A _10810_/B vssd1 vssd1 vccd1 vccd1 _10924_/B sky130_fd_sc_hd__or2_1
X_10741_ _10741_/A _10741_/B vssd1 vssd1 vccd1 vccd1 _10742_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08863__B1 _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12411_ reg1_val[30] _12444_/C vssd1 vssd1 vccd1 vccd1 _12411_/X sky130_fd_sc_hd__xor2_1
X_10672_ _10672_/A _10672_/B vssd1 vssd1 vccd1 vccd1 _10672_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_35_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13391_ _13392_/CLK _13391_/D vssd1 vssd1 vccd1 vccd1 hold297/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12342_ _12391_/A _12342_/B vssd1 vssd1 vccd1 vccd1 _12345_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_50_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08091__B2 _08649_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08091__A1 _08657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12273_ _06645_/B _11829_/B _11554_/A vssd1 vssd1 vccd1 vccd1 _12273_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11224_ _11224_/A _11224_/B _11224_/C vssd1 vssd1 vccd1 vccd1 _11225_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_50_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11922__B1 _06958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11155_ _11455_/B vssd1 vssd1 vccd1 vccd1 _11155_/Y sky130_fd_sc_hd__inv_2
X_11086_ _11087_/B _11087_/A vssd1 vssd1 vccd1 vccd1 _11086_/X sky130_fd_sc_hd__and2b_1
X_10106_ _09838_/A _09838_/B _09960_/B _09961_/B _09961_/A vssd1 vssd1 vccd1 vccd1
+ _10120_/A sky130_fd_sc_hd__a32oi_4
X_10037_ reg1_val[5] curr_PC[5] vssd1 vssd1 vccd1 vccd1 _10038_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08146__A2 _08289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11150__A1 _09422_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11988_ _10444_/Y _11987_/Y _12444_/B vssd1 vssd1 vccd1 vccd1 _11988_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_86_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10939_ _12336_/A _10939_/B vssd1 vssd1 vccd1 vccd1 _10943_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09004__A _09341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12609_ _12607_/X _12609_/B vssd1 vssd1 vccd1 vccd1 _12621_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_109_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12365__A _12365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10964__A1 _06998_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10964__B2 _07032_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12084__B _12084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10716__A1 _11592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10716__B2 _10944_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11913__A0 _09228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12812__B _12820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09820_ _09820_/A _09820_/B vssd1 vssd1 vccd1 vccd1 _09821_/B sky130_fd_sc_hd__nor2_1
XANTENNA__06810__B _06810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07194__A _07195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10192__A2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06963_ _12438_/A _06963_/B vssd1 vssd1 vccd1 vccd1 _06963_/Y sky130_fd_sc_hd__nand2_1
X_09751_ hold256/A _09750_/X _09238_/Y vssd1 vssd1 vccd1 vccd1 _09751_/Y sky130_fd_sc_hd__o21ai_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08702_ _07877_/X _08702_/B vssd1 vssd1 vccd1 vccd1 _08805_/A sky130_fd_sc_hd__nand2b_2
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06894_ _09218_/A _09419_/B vssd1 vssd1 vccd1 vccd1 _06894_/Y sky130_fd_sc_hd__nor2_1
X_09682_ _09682_/A _09682_/B vssd1 vssd1 vccd1 vccd1 _09683_/B sky130_fd_sc_hd__xnor2_2
X_08633_ _06992_/A _08613_/B _08613_/C _09677_/A _06993_/Y vssd1 vssd1 vccd1 vccd1
+ _08634_/B sky130_fd_sc_hd__o32ai_4
XANTENNA_fanout268_A _06810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13135__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08564_ _08564_/A _08564_/B vssd1 vssd1 vccd1 vccd1 _08570_/B sky130_fd_sc_hd__xnor2_2
X_07515_ _07515_/A _07515_/B vssd1 vssd1 vccd1 vccd1 _07705_/B sky130_fd_sc_hd__xnor2_1
Xfanout14 _12335_/A vssd1 vssd1 vccd1 vccd1 fanout14/X sky130_fd_sc_hd__clkbuf_8
Xfanout47 _07830_/B vssd1 vssd1 vccd1 vccd1 fanout47/X sky130_fd_sc_hd__clkbuf_8
Xfanout36 _07192_/Y vssd1 vssd1 vccd1 vccd1 fanout36/X sky130_fd_sc_hd__buf_4
X_08495_ _08495_/A _08495_/B vssd1 vssd1 vccd1 vccd1 _08745_/A sky130_fd_sc_hd__xor2_1
XANTENNA__08845__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout25 _07235_/Y vssd1 vssd1 vccd1 vccd1 fanout25/X sky130_fd_sc_hd__buf_6
Xfanout58 _07035_/X vssd1 vssd1 vccd1 vccd1 fanout58/X sky130_fd_sc_hd__buf_4
XFILLER_0_91_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout69 _09936_/A vssd1 vssd1 vccd1 vccd1 _12336_/A sky130_fd_sc_hd__buf_8
X_07446_ _07198_/Y fanout78/X fanout74/X _10599_/A vssd1 vssd1 vccd1 vccd1 _07447_/B
+ sky130_fd_sc_hd__o22a_1
X_07377_ _07377_/A _07377_/B vssd1 vssd1 vccd1 vccd1 _07430_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09116_ _07830_/B _10599_/A _10500_/A fanout46/X vssd1 vssd1 vccd1 vccd1 _09117_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_5_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09047_ _09064_/B _08970_/B _08983_/B _08984_/B _08984_/A vssd1 vssd1 vccd1 vccd1
+ _09063_/A sky130_fd_sc_hd__a32o_2
XFILLER_0_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06720__B _07097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09949_ _09949_/A _09949_/B vssd1 vssd1 vccd1 vccd1 _09961_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08128__A2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12960_ hold64/X hold278/X vssd1 vssd1 vccd1 vccd1 _13220_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11911_ _12271_/A1 _11992_/B hold266/A vssd1 vssd1 vccd1 vccd1 _11911_/Y sky130_fd_sc_hd__a21oi_1
X_12891_ hold275/X hold36/X vssd1 vssd1 vccd1 vccd1 _13178_/A sky130_fd_sc_hd__nand2b_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _12050_/A _12050_/B vssd1 vssd1 vccd1 vccd1 _11892_/B sky130_fd_sc_hd__and2_1
XANTENNA__07551__B _07554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12169__B _12335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _11774_/B _11773_/B vssd1 vssd1 vccd1 vccd1 _11775_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_83_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ _11844_/A _10724_/B vssd1 vssd1 vccd1 vccd1 _10726_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10655_ _10655_/A _10655_/B _10655_/C vssd1 vssd1 vccd1 vccd1 _10656_/B sky130_fd_sc_hd__nand3_2
X_13374_ _13390_/CLK _13374_/D vssd1 vssd1 vccd1 vccd1 hold270/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12325_ _12449_/B1 _12374_/B hold287/A vssd1 vssd1 vccd1 vccd1 _12325_/Y sky130_fd_sc_hd__a21oi_1
X_10586_ _11398_/A _10586_/B vssd1 vssd1 vccd1 vccd1 _10587_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_50_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_543 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12256_ _06874_/A _12254_/X _12255_/Y vssd1 vssd1 vccd1 vccd1 _12256_/X sky130_fd_sc_hd__o21a_1
X_11207_ _11207_/A _11207_/B vssd1 vssd1 vccd1 vccd1 _11214_/A sky130_fd_sc_hd__nand2_2
X_12187_ _12306_/A _12185_/X _12186_/Y vssd1 vssd1 vccd1 vccd1 _12215_/A sky130_fd_sc_hd__o21a_1
XANTENNA__07218__S _11584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10174__A2 _11554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11138_ _11138_/A _11138_/B vssd1 vssd1 vccd1 vccd1 _11138_/X sky130_fd_sc_hd__or2_1
XANTENNA__07575__B1 fanout72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11069_ _11770_/A _11069_/B vssd1 vssd1 vccd1 vccd1 _11070_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11123__A1 max_cap3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08838__A _09944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12871__A1 _08974_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07300_ fanout98/X _10473_/B2 _10240_/A fanout84/X vssd1 vssd1 vccd1 vccd1 _07301_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_128_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08573__A _08664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08280_ _08280_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08769_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07231_ _07231_/A _11473_/A vssd1 vssd1 vccd1 vccd1 _07231_/X sky130_fd_sc_hd__or2_2
XFILLER_0_74_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10608__A _11770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07189__A _09667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07162_ _07162_/A _07162_/B vssd1 vssd1 vccd1 vccd1 _07371_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_42_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07093_ _06983_/A _06983_/B _07094_/B vssd1 vssd1 vccd1 vccd1 _07093_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_42_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout204 _08658_/A vssd1 vssd1 vccd1 vccd1 _08575_/A sky130_fd_sc_hd__buf_12
XFILLER_0_10_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout226 _10165_/S vssd1 vssd1 vccd1 vccd1 _11247_/A sky130_fd_sc_hd__clkbuf_8
X_09803_ _09807_/A vssd1 vssd1 vccd1 vccd1 _09806_/A sky130_fd_sc_hd__inv_2
Xfanout215 _12808_/A vssd1 vssd1 vccd1 vccd1 _09404_/S sky130_fd_sc_hd__buf_6
Xfanout237 _06993_/Y vssd1 vssd1 vccd1 vccd1 _08613_/A sky130_fd_sc_hd__buf_6
XFILLER_0_10_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout259 _13248_/A2 vssd1 vssd1 vccd1 vccd1 _13223_/B2 sky130_fd_sc_hd__buf_4
Xfanout248 _12218_/A vssd1 vssd1 vccd1 vccd1 _11752_/S sky130_fd_sc_hd__buf_12
X_07995_ _09836_/A _07993_/B _08066_/A vssd1 vssd1 vccd1 vccd1 _08059_/A sky130_fd_sc_hd__o21ai_2
X_06946_ _09234_/C _09234_/B _09233_/B vssd1 vssd1 vccd1 vccd1 _06946_/X sky130_fd_sc_hd__and3b_4
X_09734_ reg1_val[3] curr_PC[3] vssd1 vssd1 vccd1 vccd1 _09734_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13103__A2 fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07318__B1 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11665__A2 _08974_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06877_ _06877_/A _06877_/B vssd1 vssd1 vccd1 vccd1 _06877_/Y sky130_fd_sc_hd__nand2_1
X_09665_ _09665_/A _09665_/B vssd1 vssd1 vccd1 vccd1 _09668_/A sky130_fd_sc_hd__nand2_1
X_08616_ _07030_/Y _07166_/Y _07173_/Y _07038_/X vssd1 vssd1 vccd1 vccd1 _08617_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08530__A2 _08561_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ _12064_/S _09596_/B vssd1 vssd1 vccd1 vccd1 _09596_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08547_ _08550_/B _08550_/C _08550_/A vssd1 vssd1 vccd1 vccd1 _08739_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__08818__B1 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12090__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09491__B1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08294__A1 _08641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08294__B2 _08627_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08478_ _08580_/A _08478_/B vssd1 vssd1 vccd1 vccd1 _08511_/A sky130_fd_sc_hd__xor2_2
X_07429_ _07429_/A _07429_/B vssd1 vssd1 vccd1 vccd1 _07678_/A sky130_fd_sc_hd__and2_2
X_10440_ hold252/A _09425_/C _10438_/X _12416_/C1 vssd1 vssd1 vccd1 vccd1 _10440_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10928__A1 _12144_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10371_ _10950_/A _10371_/B vssd1 vssd1 vccd1 vccd1 _10501_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_33_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12110_ _12111_/A _12111_/B _12111_/C vssd1 vssd1 vccd1 vccd1 _12110_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__06731__A _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13090_ hold13/X _12805_/A _13250_/B _13355_/Q _13039_/A vssd1 vssd1 vccd1 vccd1
+ hold14/A sky130_fd_sc_hd__o221a_1
X_12041_ _12041_/A _12041_/B vssd1 vssd1 vccd1 vccd1 _12300_/A sky130_fd_sc_hd__or2_2
Xhold280 hold280/A vssd1 vssd1 vccd1 vccd1 hold280/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 hold291/A vssd1 vssd1 vccd1 vccd1 hold291/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07038__S _09673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07021__A2 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08658__A _08658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12853__A1 _07013_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12943_ _13183_/A _13184_/A _13183_/B vssd1 vssd1 vccd1 vccd1 _13189_/A sky130_fd_sc_hd__a21bo_1
X_12874_ _12874_/A _12874_/B vssd1 vssd1 vccd1 vccd1 _13243_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11825_ _11825_/A _11825_/B vssd1 vssd1 vccd1 vccd1 _11825_/X sky130_fd_sc_hd__or2_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11756_ fanout58/X fanout10/X fanout5/X _11868_/A vssd1 vssd1 vccd1 vccd1 _11757_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707_ _10707_/A _10707_/B vssd1 vssd1 vccd1 vccd1 _10709_/C sky130_fd_sc_hd__xor2_1
X_11687_ _11687_/A _11687_/B vssd1 vssd1 vccd1 vccd1 _11703_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_102_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10638_ _10638_/A _10638_/B vssd1 vssd1 vccd1 vccd1 _10651_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10569_ hold252/A hold281/A _10569_/C vssd1 vssd1 vccd1 vccd1 _10690_/B sky130_fd_sc_hd__or3_1
X_13357_ _13358_/CLK _13357_/D vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__dfxtp_1
X_13288_ _13385_/CLK _13288_/D vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__dfxtp_1
X_12308_ _12399_/A _12307_/X _09150_/X vssd1 vssd1 vccd1 vccd1 _12308_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12239_ _12239_/A _12239_/B _12239_/C vssd1 vssd1 vccd1 vccd1 _12240_/B sky130_fd_sc_hd__nor3_1
XANTENNA__13097__A1 _09936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06800_ reg1_val[3] _07165_/A vssd1 vssd1 vccd1 vccd1 _06800_/Y sky130_fd_sc_hd__nor2_1
X_07780_ _07776_/Y _07845_/B _07775_/Y vssd1 vssd1 vccd1 vccd1 _07867_/A sky130_fd_sc_hd__a21o_1
X_06731_ _11242_/A _07262_/A vssd1 vssd1 vccd1 vccd1 _11259_/S sky130_fd_sc_hd__and2_1
XANTENNA__10855__B1 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09450_ _07554_/B _07232_/X _07238_/Y _07175_/A vssd1 vssd1 vccd1 vccd1 _09451_/B
+ sky130_fd_sc_hd__a22o_1
X_06662_ instruction[41] _06927_/A _06617_/B _06660_/X vssd1 vssd1 vccd1 vccd1 _07147_/B
+ sky130_fd_sc_hd__a31o_4
X_08401_ _08431_/B _08431_/A vssd1 vssd1 vccd1 vccd1 _08403_/B sky130_fd_sc_hd__nand2b_1
X_06593_ instruction[20] _06944_/B vssd1 vssd1 vccd1 vccd1 _06593_/X sky130_fd_sc_hd__or2_1
X_09381_ _09379_/X _09380_/X _09725_/S vssd1 vssd1 vccd1 vccd1 _09381_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10607__B1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09473__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08332_ _08540_/B _08561_/A2 _08561_/B1 _08515_/A2 vssd1 vssd1 vccd1 vccd1 _08333_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08263_ _08263_/A _08263_/B vssd1 vssd1 vccd1 vccd1 _08264_/B sky130_fd_sc_hd__and2_1
X_07214_ _07133_/A _06974_/B _07215_/B vssd1 vssd1 vccd1 vccd1 _07214_/X sky130_fd_sc_hd__o21a_1
XANTENNA_fanout133_A _10245_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08194_ _08598_/B _08457_/A2 _08501_/B1 _08538_/A1 vssd1 vssd1 vccd1 vccd1 _08195_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07145_ reg1_val[26] _07585_/B1 _07154_/B vssd1 vssd1 vccd1 vccd1 _07146_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08579__A2 _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11583__B2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11583__A1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10386__A2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07076_ _07087_/A _07094_/B vssd1 vssd1 vccd1 vccd1 _07078_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_15_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07787__B1 _07283_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09862__A _09862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07978_ _08580_/A _07978_/B vssd1 vssd1 vccd1 vccd1 _08023_/A sky130_fd_sc_hd__xnor2_1
X_06929_ instruction[12] _06933_/B vssd1 vssd1 vccd1 vccd1 dest_idx[1] sky130_fd_sc_hd__and2_4
X_09717_ _12364_/A _09717_/B _09717_/C vssd1 vssd1 vccd1 vccd1 _09717_/X sky130_fd_sc_hd__or3_1
XANTENNA__08478__A _08580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12835__A1 _07274_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08503__A2 _08561_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10846__B1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09648_ _10748_/A _09648_/B vssd1 vssd1 vccd1 vccd1 _09653_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ reg1_val[2] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _09580_/B sky130_fd_sc_hd__nand2_1
X_11610_ _11610_/A _11610_/B vssd1 vssd1 vccd1 vccd1 _11612_/C sky130_fd_sc_hd__xnor2_1
X_12590_ _12598_/C _12590_/B vssd1 vssd1 vccd1 vccd1 _12597_/C sky130_fd_sc_hd__nand2_2
XANTENNA__11632__A _11813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11541_ _11541_/A _11541_/B vssd1 vssd1 vccd1 vccd1 _11541_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13260__B2 _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06817__A2 _06766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11472_ _12050_/A _11567_/B _11567_/C vssd1 vssd1 vccd1 vccd1 _11472_/X sky130_fd_sc_hd__and3_1
XFILLER_0_18_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13211_ _13211_/A _13211_/B vssd1 vssd1 vccd1 vccd1 _13212_/B sky130_fd_sc_hd__nand2_1
X_10423_ _10423_/A _10423_/B vssd1 vssd1 vccd1 vccd1 _10423_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10682__S _11029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10354_ _10247_/A _10249_/B _10355_/B vssd1 vssd1 vccd1 vccd1 _10354_/Y sky130_fd_sc_hd__a21oi_1
X_13142_ _13142_/A hold253/X vssd1 vssd1 vccd1 vccd1 _13369_/D sky130_fd_sc_hd__and2_1
XANTENNA__07778__B1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11079__A _11182_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08990__A2 _11946_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13073_ _11182_/A _13089_/A2 hold101/X vssd1 vssd1 vccd1 vccd1 hold102/A sky130_fd_sc_hd__o21a_1
X_10285_ _10187_/X _10581_/A _10284_/Y vssd1 vssd1 vccd1 vccd1 _10285_/Y sky130_fd_sc_hd__a21oi_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12024_ _12024_/A _12024_/B vssd1 vssd1 vccd1 vccd1 _12025_/B sky130_fd_sc_hd__and2_1
XANTENNA__08388__A _08580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12926_ hold32/X hold252/X vssd1 vssd1 vccd1 vccd1 _13143_/B sky130_fd_sc_hd__nand2b_1
X_12857_ _07032_/Y _12863_/A2 hold78/X _13249_/A vssd1 vssd1 vccd1 vccd1 _13289_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11808_ _11807_/A _11807_/B _09150_/X vssd1 vssd1 vccd1 vccd1 _11808_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_95_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12788_ _12788_/A _12788_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[29] sky130_fd_sc_hd__xnor2_4
XANTENNA__09455__B1 _12823_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11739_ hold262/A _11739_/B vssd1 vssd1 vccd1 vccd1 _11822_/B sky130_fd_sc_hd__or2_1
XFILLER_0_71_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09947__A _09947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13409_ instruction[10] vssd1 vssd1 vccd1 vccd1 pred_idx[2] sky130_fd_sc_hd__buf_12
XANTENNA__09758__A1 _12446_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08950_ _10749_/A _08950_/B vssd1 vssd1 vccd1 vccd1 _08954_/A sky130_fd_sc_hd__xnor2_1
X_07901_ _07932_/A _07932_/B vssd1 vssd1 vccd1 vccd1 _07901_/Y sky130_fd_sc_hd__nor2_1
X_08881_ _08882_/A _08882_/B vssd1 vssd1 vccd1 vccd1 _08881_/X sky130_fd_sc_hd__or2_1
XANTENNA__12312__S _12404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12820__B _12820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07832_ _07983_/A _07907_/B _07907_/C vssd1 vssd1 vccd1 vccd1 _07834_/C sky130_fd_sc_hd__and3_1
XFILLER_0_47_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08194__B1 _08501_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12817__A1 _07134_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09502_ _09671_/A _09502_/B vssd1 vssd1 vccd1 vccd1 _09505_/A sky130_fd_sc_hd__xnor2_2
X_07763_ _07763_/A _07763_/B vssd1 vssd1 vccd1 vccd1 _07824_/A sky130_fd_sc_hd__xor2_2
XANTENNA__10828__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06714_ reg1_val[18] _07088_/A vssd1 vssd1 vccd1 vccd1 _06715_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_79_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07694_ _06993_/Y fanout63/X fanout57/X _06993_/A vssd1 vssd1 vccd1 vccd1 _07695_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_94_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout250_A _06782_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06645_ _06643_/X _06645_/B vssd1 vssd1 vccd1 vccd1 _06874_/A sky130_fd_sc_hd__nand2b_2
X_09433_ _12365_/A _09433_/B vssd1 vssd1 vccd1 vccd1 _09433_/Y sky130_fd_sc_hd__nand2_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09364_ _09364_/A _09364_/B vssd1 vssd1 vccd1 vccd1 _09366_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06576_ hold165/A vssd1 vssd1 vccd1 vccd1 _06576_/Y sky130_fd_sc_hd__inv_2
X_08315_ _08315_/A _08315_/B vssd1 vssd1 vccd1 vccd1 _08316_/B sky130_fd_sc_hd__or2_1
XANTENNA_31 reg2_val[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_20 reg1_val[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09295_ _09296_/B _09295_/B vssd1 vssd1 vccd1 vccd1 _09467_/B sky130_fd_sc_hd__and2b_1
XANTENNA_42 _07221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_53 reg1_val[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ _08246_/A _08246_/B vssd1 vssd1 vccd1 vccd1 _08313_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07472__A2 _07959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08177_ _08177_/A _08177_/B vssd1 vssd1 vccd1 vccd1 _08779_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__11556__B2 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11556__A1 _10159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10359__A2 _07269_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07128_ _07129_/C _07129_/D vssd1 vssd1 vccd1 vccd1 _07128_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_42_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07059_ _07059_/A _07059_/B vssd1 vssd1 vccd1 vccd1 _07102_/B sky130_fd_sc_hd__xor2_1
X_10070_ _10245_/A1 fanout14/X fanout13/X _10245_/B2 vssd1 vssd1 vccd1 vccd1 _10071_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09921__B2 _07554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09921__A1 _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10972_ _10972_/A _10972_/B vssd1 vssd1 vccd1 vccd1 _10973_/B sky130_fd_sc_hd__and2_1
XANTENNA__06684__A_N _07014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08936__A _09922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12711_ _12711_/A _12711_/B _12711_/C vssd1 vssd1 vccd1 vccd1 _12712_/B sky130_fd_sc_hd__nand3_1
XANTENNA__07840__A _09673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12642_ _12642_/A _12642_/B vssd1 vssd1 vccd1 vccd1 _12643_/B sky130_fd_sc_hd__or2_1
XANTENNA__07160__B2 _07959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07160__A1 _07148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12573_ _12582_/A _12573_/B vssd1 vssd1 vccd1 vccd1 new_PC[16] sky130_fd_sc_hd__and2_4
XFILLER_0_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11081__B fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11524_ _11524_/A _11524_/B _11524_/C vssd1 vssd1 vccd1 vccd1 _11525_/B sky130_fd_sc_hd__nand3_2
XANTENNA__12992__B1 _13257_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11455_ _12064_/S _11455_/B vssd1 vssd1 vccd1 vccd1 _11455_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10706__A _10707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10406_ _10268_/A _10268_/B _10266_/Y vssd1 vssd1 vccd1 vccd1 _10408_/B sky130_fd_sc_hd__a21boi_1
X_11386_ _11387_/A _11387_/B vssd1 vssd1 vccd1 vccd1 _11509_/A sky130_fd_sc_hd__or2_1
XFILLER_0_104_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10337_ _10337_/A _12428_/B vssd1 vssd1 vccd1 vccd1 _10341_/A sky130_fd_sc_hd__nand2_1
X_13125_ hold290/A _13124_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13125_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10268_ _10268_/A _10268_/B vssd1 vssd1 vccd1 vccd1 _10270_/B sky130_fd_sc_hd__xnor2_2
X_13056_ hold150/X _13094_/A2 _13101_/A2 hold145/X _13259_/A vssd1 vssd1 vccd1 vccd1
+ hold151/A sky130_fd_sc_hd__o221a_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12007_ _12093_/A fanout7/X vssd1 vssd1 vccd1 vccd1 _12007_/Y sky130_fd_sc_hd__nor2_1
X_10199_ _11592_/A _07213_/Y fanout30/X _10944_/B2 vssd1 vssd1 vccd1 vccd1 _10200_/B
+ sky130_fd_sc_hd__a22o_2
XANTENNA__11483__B1 _08859_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12909_ hold235/X hold70/X vssd1 vssd1 vccd1 vccd1 _13110_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__08846__A _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12087__B _12087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10589__A2 _07256_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09677__A _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08100_ _08097_/Y _08155_/B _08096_/Y vssd1 vssd1 vccd1 vccd1 _08116_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07454__A2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09080_ fanout53/X fanout86/X fanout82/X fanout51/X vssd1 vssd1 vccd1 vccd1 _09081_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08031_ _08454_/A _08031_/B vssd1 vssd1 vccd1 vccd1 _08036_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06813__B _07149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09982_ _09982_/A _09982_/B vssd1 vssd1 vccd1 vccd1 _09983_/B sky130_fd_sc_hd__nand2_1
X_08933_ _08933_/A _08933_/B vssd1 vssd1 vccd1 vccd1 _08934_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11447__A _11813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07914__B1 _07097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08864_ _09947_/A _08864_/B vssd1 vssd1 vccd1 vccd1 _08866_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_74_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08795_ _08795_/A _08795_/B vssd1 vssd1 vccd1 vccd1 _12129_/C sky130_fd_sc_hd__nor2_1
X_07815_ _07813_/A _07813_/B _07814_/Y vssd1 vssd1 vccd1 vccd1 _08706_/A sky130_fd_sc_hd__a21bo_2
X_07746_ _07816_/A _07816_/B _07680_/X vssd1 vssd1 vccd1 vccd1 _08708_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__11182__A _11182_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ hold293/A _11538_/A hold301/A vssd1 vssd1 vccd1 vccd1 _09416_/Y sky130_fd_sc_hd__a21oi_1
X_07677_ _07677_/A _07677_/B vssd1 vssd1 vccd1 vccd1 _08708_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_109_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12018__A2 _07608_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06628_ reg2_val[28] _06766_/B _06724_/B1 _06627_/Y vssd1 vssd1 vccd1 vccd1 _06867_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_09347_ _09347_/A _09347_/B vssd1 vssd1 vccd1 vccd1 _09350_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12974__B1 fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09278_ _09278_/A _09278_/B _09278_/C vssd1 vssd1 vccd1 vccd1 _09279_/B sky130_fd_sc_hd__and3_1
XFILLER_0_117_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08229_ _08278_/A _08278_/B vssd1 vssd1 vccd1 vccd1 _08229_/X sky130_fd_sc_hd__or2_1
XANTENNA__06723__B _12645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11240_ _11239_/A _11239_/B _11239_/Y _09225_/Y vssd1 vssd1 vccd1 vccd1 _11265_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11171_ fanout52/X fanout23/X fanout16/X _11476_/A vssd1 vssd1 vccd1 vccd1 _11172_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10122_ _09984_/A _09983_/B _09981_/Y vssd1 vssd1 vccd1 vccd1 _10132_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_100_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10053_ _09956_/Y _09958_/Y _07282_/Y _11946_/C vssd1 vssd1 vccd1 vccd1 _10053_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07554__B _07554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11465__B1 _09238_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11092__A _12336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10955_ _10956_/A _10956_/B vssd1 vssd1 vccd1 vccd1 _10967_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_58_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08330__B1 _09940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10886_ _10886_/A _10886_/B vssd1 vssd1 vccd1 vccd1 _10888_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12625_ reg1_val[25] curr_PC[25] _12638_/S vssd1 vssd1 vccd1 vccd1 _12627_/B sky130_fd_sc_hd__mux2_1
X_12556_ _12714_/B _12557_/B vssd1 vssd1 vccd1 vccd1 _12567_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11820__A _11820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08633__A1 _06992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09497__A _09667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11507_ _11399_/A _11399_/B _11396_/A vssd1 vssd1 vccd1 vccd1 _11509_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08633__B2 _06993_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06633__B _06675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12487_ _12660_/B _12487_/B vssd1 vssd1 vccd1 vccd1 _12488_/B sky130_fd_sc_hd__or2_1
XFILLER_0_80_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10991__A2 _12087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11438_ _11011_/X _11801_/A _11802_/A vssd1 vssd1 vccd1 vccd1 _11438_/Y sky130_fd_sc_hd__a21oi_1
Xhold109 hold109/A vssd1 vssd1 vccd1 vccd1 hold109/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11369_ _09225_/Y _11348_/Y _11349_/X _11368_/X vssd1 vssd1 vccd1 vccd1 _11369_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13108_ hold235/X _13254_/A2 _13107_/X _06577_/A vssd1 vssd1 vccd1 vccd1 hold236/A
+ sky130_fd_sc_hd__a22o_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13039_ _13039_/A hold120/X vssd1 vssd1 vccd1 vccd1 _13329_/D sky130_fd_sc_hd__and2_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08580_ _08580_/A _08580_/B vssd1 vssd1 vccd1 vccd1 _08582_/B sky130_fd_sc_hd__xor2_1
X_07600_ _07601_/A _07601_/B _07601_/C vssd1 vssd1 vccd1 vccd1 _07602_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_89_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09649__B1 _09943_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07531_ _07531_/A _07531_/B vssd1 vssd1 vccd1 vccd1 _07533_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_88_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06808__B _07172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07462_ _07540_/A _07540_/B _07458_/X vssd1 vssd1 vccd1 vccd1 _07563_/A sky130_fd_sc_hd__o21ai_2
X_09201_ _11134_/A reg1_val[17] _09211_/S vssd1 vssd1 vccd1 vccd1 _09201_/X sky130_fd_sc_hd__mux2_1
X_07393_ _07394_/A _07394_/B vssd1 vssd1 vccd1 vccd1 _07400_/B sky130_fd_sc_hd__and2_1
XFILLER_0_9_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09132_ _08939_/A _08939_/B _08942_/A vssd1 vssd1 vccd1 vccd1 _09137_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_8_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout213_A _07959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09063_ _09063_/A _09063_/B vssd1 vssd1 vccd1 vccd1 _09130_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_102_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08014_ _08014_/A _08014_/B vssd1 vssd1 vccd1 vccd1 _08015_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_102_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09965_ _09965_/A _09965_/B vssd1 vssd1 vccd1 vccd1 _09966_/B sky130_fd_sc_hd__and2_1
XFILLER_0_0_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11177__A _11582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10081__A _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09896_ reg1_val[4] curr_PC[4] vssd1 vssd1 vccd1 vccd1 _09896_/Y sky130_fd_sc_hd__nor2_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08916_ _08917_/A _08917_/B vssd1 vssd1 vccd1 vccd1 _08916_/X sky130_fd_sc_hd__and2_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08847_ _08199_/B _11093_/A _10974_/A fanout33/X vssd1 vssd1 vccd1 vccd1 _08848_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_99_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07390__A _10092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08778_ _08176_/Y _08229_/X _08175_/Y vssd1 vssd1 vccd1 vccd1 _08791_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_95_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07729_ _07806_/A _07806_/B _07722_/X vssd1 vssd1 vccd1 vccd1 _07750_/A sky130_fd_sc_hd__a21oi_1
X_10740_ _10740_/A _10740_/B vssd1 vssd1 vccd1 vccd1 _10741_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_95_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11998__A1 _10159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11998__B2 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08863__A1 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10671_ _06836_/Y _10670_/Y _12054_/S vssd1 vssd1 vccd1 vccd1 _10672_/B sky130_fd_sc_hd__mux2_1
XANTENNA__08863__B2 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12410_ _09040_/C _12408_/X _12409_/Y vssd1 vssd1 vccd1 vccd1 _12425_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_35_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13390_ _13390_/CLK _13390_/D vssd1 vssd1 vccd1 vccd1 hold258/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09812__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12341_ _12341_/A _12341_/B vssd1 vssd1 vccd1 vccd1 _12342_/B sky130_fd_sc_hd__or2_1
XFILLER_0_63_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08091__A2 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12272_ hold282/A _12449_/B1 _12324_/B _12271_/Y _12376_/C1 vssd1 vssd1 vccd1 vccd1
+ _12272_/X sky130_fd_sc_hd__a311o_1
X_11223_ _11224_/A _11224_/B _11224_/C vssd1 vssd1 vccd1 vccd1 _11223_/Y sky130_fd_sc_hd__a21oi_1
X_11154_ _11247_/A _09407_/X _09251_/A vssd1 vssd1 vccd1 vccd1 _11455_/B sky130_fd_sc_hd__o21a_1
X_11085_ _11201_/A _11085_/B vssd1 vssd1 vccd1 vccd1 _11087_/B sky130_fd_sc_hd__nor2_1
X_10105_ _10105_/A _10105_/B vssd1 vssd1 vccd1 vccd1 _10121_/A sky130_fd_sc_hd__and2_2
X_10036_ reg1_val[5] curr_PC[5] vssd1 vssd1 vccd1 vccd1 _10036_/Y sky130_fd_sc_hd__nor2_1
X_11987_ _11987_/A _11987_/B vssd1 vssd1 vccd1 vccd1 _11987_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10938_ _11406_/A _07362_/B fanout16/X _11309_/A vssd1 vssd1 vccd1 vccd1 _10939_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_105_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10869_ _10990_/B _10869_/B vssd1 vssd1 vccd1 vccd1 _10877_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_39_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12608_ _12633_/A _12608_/B vssd1 vssd1 vccd1 vccd1 _12609_/B sky130_fd_sc_hd__or2_1
XFILLER_0_30_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12539_ _12539_/A _12539_/B _12539_/C vssd1 vssd1 vccd1 vccd1 _12540_/B sky130_fd_sc_hd__nand3_1
XANTENNA__10964__A2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09955__A _11179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10716__A2 _07171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06962_ _12404_/S _06962_/B vssd1 vssd1 vccd1 vccd1 _06962_/Y sky130_fd_sc_hd__nor2_1
X_09750_ hold295/A hold235/A hold245/A _09425_/C vssd1 vssd1 vccd1 vccd1 _09750_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09681_ _09682_/A _09682_/B vssd1 vssd1 vccd1 vccd1 _09681_/Y sky130_fd_sc_hd__nand2b_1
X_08701_ _07950_/B _08702_/B _07877_/X vssd1 vssd1 vccd1 vccd1 _08701_/X sky130_fd_sc_hd__a21o_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06893_ _06992_/A _12808_/A vssd1 vssd1 vccd1 vccd1 _08663_/A sky130_fd_sc_hd__nor2_2
X_08632_ _09673_/A _08632_/B vssd1 vssd1 vccd1 vccd1 _08640_/A sky130_fd_sc_hd__xor2_2
XANTENNA__06819__A _12644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout163_A _12322_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08563_ _08593_/A _08593_/B vssd1 vssd1 vccd1 vccd1 _08594_/A sky130_fd_sc_hd__nor2_2
X_08494_ _08495_/A _08495_/B vssd1 vssd1 vccd1 vccd1 _08749_/A sky130_fd_sc_hd__or2_1
X_07514_ _10207_/A _07514_/B vssd1 vssd1 vccd1 vccd1 _07705_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08845__A1 _09661_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout26 _07235_/Y vssd1 vssd1 vccd1 vccd1 fanout26/X sky130_fd_sc_hd__clkbuf_8
Xfanout15 fanout16/X vssd1 vssd1 vccd1 vccd1 fanout15/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_71_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout37 _07174_/X vssd1 vssd1 vccd1 vccd1 _07175_/A sky130_fd_sc_hd__buf_6
XFILLER_0_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08845__B2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07445_ _10749_/A _07445_/B vssd1 vssd1 vccd1 vccd1 _07451_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12556__A _12714_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout59 _07033_/X vssd1 vssd1 vccd1 vccd1 fanout59/X sky130_fd_sc_hd__buf_8
Xfanout48 _07131_/Y vssd1 vssd1 vccd1 vccd1 _07830_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07376_ _07376_/A _07376_/B vssd1 vssd1 vccd1 vccd1 _07377_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09115_ _09341_/A _09115_/B vssd1 vssd1 vccd1 vccd1 _09119_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09046_ _09027_/A _09027_/B _09028_/Y vssd1 vssd1 vccd1 vccd1 _09144_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_4_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10168__B1 _12205_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09948_ _09949_/A _09949_/B vssd1 vssd1 vccd1 vccd1 _09948_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout76_A _11093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09879_ _11028_/S _09726_/X _11247_/C vssd1 vssd1 vccd1 vccd1 _09879_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__08533__B1 _09940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11910_ hold268/A _11910_/B vssd1 vssd1 vccd1 vccd1 _11992_/B sky130_fd_sc_hd__or2_1
X_12890_ hold292/A hold87/X vssd1 vssd1 vccd1 vccd1 _13183_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07832__B _07907_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _11841_/A _11841_/B _11841_/C _11807_/B vssd1 vssd1 vccd1 vccd1 _12050_/B
+ sky130_fd_sc_hd__nor4b_2
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _11929_/A _11772_/B vssd1 vssd1 vccd1 vccd1 _11773_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10723_ _07269_/Y _07596_/A _07596_/B _07360_/X _07262_/X vssd1 vssd1 vccd1 vccd1
+ _10724_/B sky130_fd_sc_hd__a32o_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12466__A _12645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10654_ _10655_/A _10655_/B _10655_/C vssd1 vssd1 vccd1 vccd1 _10656_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_36_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10585_ _10944_/B2 _07171_/A _07175_/A _07097_/X vssd1 vssd1 vccd1 vccd1 _10586_/B
+ sky130_fd_sc_hd__a22o_1
X_13373_ _13373_/CLK _13373_/D vssd1 vssd1 vccd1 vccd1 hold285/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12324_ hold282/A _12324_/B vssd1 vssd1 vccd1 vccd1 _12374_/B sky130_fd_sc_hd__or2_1
XFILLER_0_106_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12148__A1 _09242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10714__A _12096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12255_ _06874_/A _12254_/X _11637_/A vssd1 vssd1 vccd1 vccd1 _12255_/Y sky130_fd_sc_hd__a21oi_1
X_11206_ _11107_/A _11107_/B _11105_/Y vssd1 vssd1 vccd1 vccd1 _11215_/A sky130_fd_sc_hd__a21bo_1
X_12186_ _12306_/A _12185_/X _09150_/X vssd1 vssd1 vccd1 vccd1 _12186_/Y sky130_fd_sc_hd__a21oi_1
X_11137_ _11137_/A _11137_/B vssd1 vssd1 vccd1 vccd1 _11137_/X sky130_fd_sc_hd__xor2_1
XANTENNA__07575__A1 _10871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07575__B2 _08199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11068_ _12169_/A fanout32/X fanout30/X _06998_/X vssd1 vssd1 vccd1 vccd1 _11069_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12320__A1 _12412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11659__B1 _12471_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10019_ _10297_/S _09402_/X _10018_/X vssd1 vssd1 vccd1 vccd1 _10020_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07230_ _11381_/A _07230_/B vssd1 vssd1 vccd1 vccd1 _11473_/A sky130_fd_sc_hd__and2_1
XFILLER_0_41_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12387__A1 _08859_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07161_ _09779_/A _07161_/B vssd1 vssd1 vccd1 vccd1 _07162_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_26_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10937__A2 _11050_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07263__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07092_ _10350_/A _07092_/B vssd1 vssd1 vccd1 vccd1 _07092_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_42_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06821__B _10297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout205 _07604_/A vssd1 vssd1 vccd1 vccd1 _09673_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout227 _07117_/C vssd1 vssd1 vccd1 vccd1 _10165_/S sky130_fd_sc_hd__clkbuf_4
X_09802_ _11582_/A _09802_/B vssd1 vssd1 vccd1 vccd1 _09807_/A sky130_fd_sc_hd__xnor2_1
Xfanout216 _09103_/A vssd1 vssd1 vccd1 vccd1 _12808_/A sky130_fd_sc_hd__buf_8
Xfanout238 _08502_/A vssd1 vssd1 vccd1 vccd1 _08664_/A sky130_fd_sc_hd__buf_12
Xfanout249 _12444_/B vssd1 vssd1 vccd1 vccd1 _12064_/S sky130_fd_sc_hd__clkbuf_8
X_07994_ _08065_/A _08065_/B _08065_/C vssd1 vssd1 vccd1 vccd1 _08066_/A sky130_fd_sc_hd__a21o_1
X_06945_ instruction[23] _06590_/X _06944_/X _06716_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[5]
+ sky130_fd_sc_hd__o211a_4
XANTENNA__12847__C1 _13019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09733_ _09581_/A _09578_/Y _09580_/B vssd1 vssd1 vccd1 vccd1 _09733_/X sky130_fd_sc_hd__o21a_1
XANTENNA__08515__B1 _08649_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07318__A1 _06993_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07318__B2 _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06876_ _06867_/Y _06875_/X _06673_/A vssd1 vssd1 vccd1 vccd1 _06877_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11455__A _12064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09664_ _09664_/A _09664_/B vssd1 vssd1 vccd1 vccd1 _09665_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_96_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09595_ _11813_/S _09562_/Y _09594_/X _09222_/B vssd1 vssd1 vccd1 vccd1 _09602_/B
+ sky130_fd_sc_hd__o211a_1
X_08615_ _09672_/A _08615_/B _08615_/C vssd1 vssd1 vccd1 vccd1 _08618_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08546_ _08567_/B _08567_/A vssd1 vssd1 vccd1 vccd1 _08550_/C sky130_fd_sc_hd__and2b_1
XANTENNA__08818__A1 _07134_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08818__B2 _07166_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12286__A _12286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09491__A1 _09661_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09491__B2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08294__A2 _08457_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08477_ _08598_/B _08561_/B1 _08576_/A2 _08538_/A1 vssd1 vssd1 vccd1 vccd1 _08478_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_119_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07428_ _07428_/A _07428_/B _07428_/C vssd1 vssd1 vccd1 vccd1 _07429_/B sky130_fd_sc_hd__or3_1
XFILLER_0_9_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07359_ reg1_val[28] _07359_/B vssd1 vssd1 vccd1 vccd1 _07361_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_115_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10370_ _07255_/Y _10476_/B _10476_/C _10476_/A _12233_/B vssd1 vssd1 vccd1 vccd1
+ _10371_/B sky130_fd_sc_hd__o32a_1
XFILLER_0_33_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06731__B _07262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09029_ _09029_/A _09029_/B vssd1 vssd1 vccd1 vccd1 _09031_/B sky130_fd_sc_hd__xnor2_4
Xhold270 hold270/A vssd1 vssd1 vccd1 vccd1 hold270/X sky130_fd_sc_hd__buf_1
X_12040_ _12040_/A _12040_/B _12040_/C vssd1 vssd1 vccd1 vccd1 _12041_/B sky130_fd_sc_hd__and3_1
Xhold292 hold292/A vssd1 vssd1 vccd1 vccd1 hold292/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 hold281/A vssd1 vssd1 vccd1 vccd1 hold281/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_12_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12942_ hold87/X hold292/A vssd1 vssd1 vccd1 vccd1 _13183_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12853__A2 _12863_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12873_ hold258/A hold26/X vssd1 vssd1 vccd1 vccd1 _12874_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_99_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11824_ hold268/A _11650_/B _11910_/B _12376_/C1 vssd1 vssd1 vccd1 vccd1 _11825_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11755_ _12336_/A _11755_/B vssd1 vssd1 vccd1 vccd1 _11763_/A sky130_fd_sc_hd__xnor2_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10706_ _10707_/A _10707_/B vssd1 vssd1 vccd1 vccd1 _10882_/A sky130_fd_sc_hd__or2_1
XFILLER_0_126_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11686_ _11778_/B _11686_/B vssd1 vssd1 vccd1 vccd1 _11687_/B sky130_fd_sc_hd__or2_1
XANTENNA__12369__A1 _12412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10637_ _10638_/A _10638_/B vssd1 vssd1 vccd1 vccd1 _10637_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_11_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10568_ _06765_/B _11829_/B _11554_/A vssd1 vssd1 vccd1 vccd1 _10568_/Y sky130_fd_sc_hd__a21oi_1
X_13356_ _13358_/CLK hold118/X vssd1 vssd1 vccd1 vccd1 hold143/A sky130_fd_sc_hd__dfxtp_1
X_13287_ _13385_/CLK _13287_/D vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12135__S _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12307_ _12050_/X _12306_/X _11892_/A vssd1 vssd1 vccd1 vccd1 _12307_/X sky130_fd_sc_hd__a21o_1
X_10499_ _10634_/B _10499_/B vssd1 vssd1 vccd1 vccd1 _10516_/A sky130_fd_sc_hd__and2_1
XFILLER_0_121_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12238_ _12239_/A _12239_/B _12239_/C vssd1 vssd1 vccd1 vccd1 _12296_/B sky130_fd_sc_hd__o21a_1
XANTENNA__06641__B _12702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12169_ _12169_/A _12335_/B vssd1 vssd1 vccd1 vccd1 _12170_/B sky130_fd_sc_hd__nor2_1
XANTENNA__13097__A2 _12820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11275__A _11929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06730_ _06815_/A _12796_/A _06817_/B1 _06729_/X vssd1 vssd1 vccd1 vccd1 _07262_/A
+ sky130_fd_sc_hd__a31o_4
XANTENNA__10855__A1 _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06661_ _06582_/Y _06677_/B1 _06660_/X vssd1 vssd1 vccd1 vccd1 _06661_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__10855__B2 _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08400_ _08400_/A _08400_/B vssd1 vssd1 vccd1 vccd1 _08431_/B sky130_fd_sc_hd__xnor2_2
X_06592_ instruction[16] _06590_/X _06591_/X _06716_/B vssd1 vssd1 vccd1 vccd1 reg1_idx[5]
+ sky130_fd_sc_hd__o211a_4
X_09380_ _09158_/X _09161_/X _09383_/S vssd1 vssd1 vccd1 vccd1 _09380_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10607__B2 _11779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10607__A1 _07013_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12818__B _12820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09473__A1 _09822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08331_ _08580_/A _08331_/B vssd1 vssd1 vccd1 vccd1 _08392_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09473__B2 _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08262_ _08272_/A _08272_/B vssd1 vssd1 vccd1 vccd1 _08262_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07484__B1 _07172_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07213_ _07213_/A _07213_/B vssd1 vssd1 vccd1 vccd1 _07213_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_6_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08193_ _08193_/A _08193_/B vssd1 vssd1 vccd1 vccd1 _08263_/A sky130_fd_sc_hd__xnor2_1
X_07144_ _11134_/A _11242_/A _07141_/C _07143_/X _07585_/B1 vssd1 vssd1 vccd1 vccd1
+ _07154_/B sky130_fd_sc_hd__o41a_1
XANTENNA__07787__A1 _09934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11583__A2 _08859_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07075_ _06983_/A _06983_/B _06980_/X _07094_/B vssd1 vssd1 vccd1 vccd1 _07088_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07787__B2 _08199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10543__B1 _10542_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ _08538_/A1 _10595_/A1 fanout72/X _08598_/B vssd1 vssd1 vccd1 vccd1 _07978_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11185__A _12093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06928_ instruction[11] _06933_/B vssd1 vssd1 vccd1 vccd1 dest_idx[0] sky130_fd_sc_hd__and2_4
X_09716_ _12364_/A _09717_/B _09717_/C vssd1 vssd1 vccd1 vccd1 _09716_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__12835__A2 _12863_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10846__A1 _11764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10846__B2 _11592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06859_ _11814_/A _06858_/Y _06857_/Y vssd1 vssd1 vccd1 vccd1 _06860_/B sky130_fd_sc_hd__o21a_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09647_ fanout65/X _10473_/B2 _10240_/A fanout59/X vssd1 vssd1 vccd1 vccd1 _09648_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ reg1_val[2] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _09578_/Y sky130_fd_sc_hd__nor2_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08529_ _08664_/A _08529_/B vssd1 vssd1 vccd1 vccd1 _08535_/A sky130_fd_sc_hd__xnor2_2
X_11540_ _06852_/X _11539_/Y _11813_/S vssd1 vssd1 vccd1 vccd1 _11541_/B sky130_fd_sc_hd__mux2_1
XANTENNA__06726__B _06727_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13260__A2 _12803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout5_A fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13012__A2 _13171_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11471_ _11471_/A _11471_/B vssd1 vssd1 vccd1 vccd1 dest_val[17] sky130_fd_sc_hd__nor2_8
XFILLER_0_33_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13210_ _13210_/A hold267/X vssd1 vssd1 vccd1 vccd1 _13383_/D sky130_fd_sc_hd__and2_1
X_10422_ _06832_/X _10421_/X _12054_/S vssd1 vssd1 vccd1 vccd1 _10423_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_61_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10353_ _10353_/A _10353_/B vssd1 vssd1 vccd1 vccd1 _10355_/B sky130_fd_sc_hd__xor2_2
X_13141_ hold252/X _13254_/A2 _13140_/X _12804_/A vssd1 vssd1 vccd1 vccd1 hold253/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07778__B2 _09298_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07778__A1 _09298_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13072_ _13345_/Q _12805_/A _13250_/B hold100/X _13039_/A vssd1 vssd1 vccd1 vccd1
+ hold101/A sky130_fd_sc_hd__o221a_1
XFILLER_0_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12023_ _12024_/A _12024_/B vssd1 vssd1 vccd1 vccd1 _12101_/B sky130_fd_sc_hd__nor2_1
X_10284_ _10187_/X _10581_/A _12356_/B1 vssd1 vssd1 vccd1 vccd1 _10284_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11807__B _11807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12925_ _13138_/A _13139_/A _13138_/B vssd1 vssd1 vccd1 vccd1 _13144_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__07163__C1 _07147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12856_ hold77/X _12870_/B vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__or2_1
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _11807_/A _11807_/B vssd1 vssd1 vccd1 vccd1 _11807_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09455__A1 _07417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13251__A2 _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12787_ _12787_/A _12787_/B vssd1 vssd1 vccd1 vccd1 _12788_/B sky130_fd_sc_hd__or2_2
XANTENNA__09455__B2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11738_ _11738_/A _11738_/B vssd1 vssd1 vccd1 vccd1 _11747_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_22_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11669_ _11783_/A _11669_/B vssd1 vssd1 vccd1 vccd1 _11674_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13408_ instruction[9] vssd1 vssd1 vccd1 vccd1 pred_idx[1] sky130_fd_sc_hd__buf_12
XFILLER_0_114_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13339_ _13358_/CLK _13339_/D vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08966__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07900_ _08000_/A _08000_/B _07897_/A vssd1 vssd1 vccd1 vccd1 _07932_/B sky130_fd_sc_hd__a21oi_2
X_08880_ _09010_/A _08880_/B vssd1 vssd1 vccd1 vccd1 _08882_/B sky130_fd_sc_hd__xor2_2
X_07831_ _07020_/A _07020_/B _06993_/A vssd1 vssd1 vccd1 vccd1 _07834_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__08194__B2 _08538_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08194__A1 _08598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12278__B1 _12277_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12817__A2 _12805_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09501_ _09672_/A _09502_/B vssd1 vssd1 vccd1 vccd1 _09501_/Y sky130_fd_sc_hd__nor2_1
X_07762_ _07763_/A _07763_/B vssd1 vssd1 vccd1 vccd1 _07762_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10828__A1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10828__B2 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06713_ reg1_val[18] _07088_/A vssd1 vssd1 vccd1 vccd1 _11553_/S sky130_fd_sc_hd__and2_1
XFILLER_0_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07693_ _07703_/B _07703_/A vssd1 vssd1 vccd1 vccd1 _07693_/X sky130_fd_sc_hd__and2b_1
XANTENNA__11733__A _11820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06644_ _07049_/A reg1_val[27] vssd1 vssd1 vccd1 vccd1 _06645_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09432_ _09432_/A _09432_/B vssd1 vssd1 vccd1 vccd1 _09433_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06575_ hold38/X vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__inv_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09363_ _09137_/A _09137_/B _09135_/Y vssd1 vssd1 vccd1 vccd1 _09364_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_19_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout243_A _12520_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08314_ _08314_/A _08314_/B vssd1 vssd1 vccd1 vccd1 _08315_/B sky130_fd_sc_hd__and2_1
XANTENNA__12450__B1 _09238_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_32 reg2_val[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 reg1_val[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_10 reg1_val[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09294_ _10479_/A _09294_/B vssd1 vssd1 vccd1 vccd1 _09296_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12564__A _12719_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_43 _10476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_54 reg1_val[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08245_ _08246_/A _08246_/B vssd1 vssd1 vccd1 vccd1 _08245_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09749__A2 _12322_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08176_ _08177_/A _08177_/B vssd1 vssd1 vccd1 vccd1 _08176_/Y sky130_fd_sc_hd__nand2_1
X_07127_ _07585_/B1 _07112_/B _07210_/B reg1_val[22] vssd1 vssd1 vccd1 vccd1 _07129_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_88_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07058_ _07059_/A _07059_/B vssd1 vssd1 vccd1 vccd1 _07363_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_11_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09921__A2 _10234_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06735__A2 _06723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10971_ _10972_/A _10972_/B vssd1 vssd1 vccd1 vccd1 _10973_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_97_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11643__A _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12710_ _12711_/A _12711_/B _12711_/C vssd1 vssd1 vccd1 vccd1 _12717_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07696__B1 _09661_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06737__A _11134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12641_ _12642_/A _12642_/B vssd1 vssd1 vccd1 vccd1 _12647_/A sky130_fd_sc_hd__nand2_2
XANTENNA__07160__A2 _07417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09437__A1 _11138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12572_ _12572_/A _12572_/B _12572_/C vssd1 vssd1 vccd1 vccd1 _12573_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_93_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08952__A _09944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11523_ _11524_/A _11524_/B _11524_/C vssd1 vssd1 vccd1 vccd1 _11523_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11454_ _11454_/A _11454_/B vssd1 vssd1 vccd1 vccd1 _11454_/Y sky130_fd_sc_hd__xnor2_1
X_10405_ _10405_/A _10405_/B vssd1 vssd1 vccd1 vccd1 _10408_/A sky130_fd_sc_hd__xnor2_1
X_11385_ _11385_/A _11385_/B vssd1 vssd1 vccd1 vccd1 _11387_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_104_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10336_ _12087_/B _10336_/B vssd1 vssd1 vccd1 vccd1 _10343_/A sky130_fd_sc_hd__xnor2_1
X_13124_ _13124_/A _13124_/B vssd1 vssd1 vccd1 vccd1 _13124_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10507__B1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10722__A _12087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10267_ _10267_/A _10267_/B vssd1 vssd1 vccd1 vccd1 _10268_/B sky130_fd_sc_hd__xnor2_2
X_13055_ _07091_/B _12820_/B hold159/X vssd1 vssd1 vccd1 vccd1 _13337_/D sky130_fd_sc_hd__a21boi_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12006_ _11929_/A _07168_/C fanout8/X _12093_/A vssd1 vssd1 vccd1 vccd1 _12006_/X
+ sky130_fd_sc_hd__o31a_1
X_10198_ _10198_/A _10198_/B vssd1 vssd1 vccd1 vccd1 _10201_/A sky130_fd_sc_hd__nor2_2
XANTENNA__11029__S _11029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11483__B2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11483__A1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13244__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12908_ hold295/A hold92/X vssd1 vssd1 vccd1 vccd1 _13115_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11272__B _12050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12839_ _07262_/X _12863_/A2 hold21/X _13249_/A vssd1 vssd1 vccd1 vccd1 _13280_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09677__B _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08030_ _08501_/B1 _08484_/B _09479_/B1 _10221_/B2 vssd1 vssd1 vccd1 vccd1 _08031_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10616__B _10707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_5_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13385_/CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA__10746__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09981_ _09982_/A _09982_/B vssd1 vssd1 vccd1 vccd1 _09981_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_12_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07611__B1 _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08932_ _08933_/A _08933_/B vssd1 vssd1 vccd1 vccd1 _08934_/A sky130_fd_sc_hd__and2_1
XANTENNA__11171__B1 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08102__A _08454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08863_ fanout68/X _09669_/B2 _09301_/A fanout65/X vssd1 vssd1 vccd1 vccd1 _08864_/B
+ sky130_fd_sc_hd__o22a_1
X_08794_ _08794_/A _08794_/B vssd1 vssd1 vccd1 vccd1 _08795_/B sky130_fd_sc_hd__xor2_4
XANTENNA__09116__B1 _10500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07814_ _07876_/B _07876_/A vssd1 vssd1 vccd1 vccd1 _07814_/Y sky130_fd_sc_hd__nand2b_1
X_07745_ _07745_/A _07745_/B vssd1 vssd1 vccd1 vccd1 _07816_/B sky130_fd_sc_hd__xor2_4
XANTENNA__11474__B2 _11582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09415_ _09222_/Y _09414_/X _09409_/Y vssd1 vssd1 vccd1 vccd1 _09415_/Y sky130_fd_sc_hd__a21oi_1
X_07676_ _07676_/A _07676_/B vssd1 vssd1 vccd1 vccd1 _09037_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_94_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06627_ _06723_/A _12708_/B vssd1 vssd1 vccd1 vccd1 _06627_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10079__A _12157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12423__B1 _12412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09346_ _11770_/A _09346_/B vssd1 vssd1 vccd1 vccd1 _09347_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12974__B2 _13000_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09277_ _09278_/A _09278_/B _09278_/C vssd1 vssd1 vccd1 vccd1 _09279_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08228_ _08278_/A _08278_/B vssd1 vssd1 vccd1 vccd1 _08228_/X sky130_fd_sc_hd__and2_1
XFILLER_0_99_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08159_ _08159_/A _08159_/B vssd1 vssd1 vccd1 vccd1 _08230_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11170_ _11318_/A _11170_/B vssd1 vssd1 vccd1 vccd1 _11174_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_101_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10121_ _10121_/A _10121_/B vssd1 vssd1 vccd1 vccd1 _10134_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_30_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10052_ _09302_/A _09947_/B _09948_/Y vssd1 vssd1 vccd1 vccd1 _10056_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_98_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06711__A2_N _06783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10954_ _10954_/A _10954_/B vssd1 vssd1 vccd1 vccd1 _10956_/B sky130_fd_sc_hd__xor2_2
XANTENNA__08330__A1 _08598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08330__B2 _08538_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10885_ _10885_/A _10885_/B vssd1 vssd1 vccd1 vccd1 _10886_/B sky130_fd_sc_hd__xnor2_1
X_12624_ _12624_/A _12624_/B vssd1 vssd1 vccd1 vccd1 new_PC[24] sky130_fd_sc_hd__xor2_4
XFILLER_0_72_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11768__A2 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12555_ _11134_/A curr_PC[14] _12638_/S vssd1 vssd1 vccd1 vccd1 _12557_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_53_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06914__B _12218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11506_ _11406_/A _12017_/A _11407_/A _11408_/Y vssd1 vssd1 vccd1 vccd1 _11511_/A
+ sky130_fd_sc_hd__o31a_1
XANTENNA__10717__A _12093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12486_ _12660_/B _12487_/B vssd1 vssd1 vccd1 vccd1 _12497_/A sky130_fd_sc_hd__nand2_1
X_11437_ _11226_/X _11623_/B _11436_/X vssd1 vssd1 vccd1 vccd1 _11802_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11368_ _06946_/X _11355_/X _11362_/X _11367_/Y vssd1 vssd1 vccd1 vccd1 _11368_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_1_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13107_ hold245/A _13106_/X fanout2/X vssd1 vssd1 vccd1 vccd1 _13107_/X sky130_fd_sc_hd__mux2_1
X_10319_ curr_PC[7] _10448_/C _10821_/A vssd1 vssd1 vccd1 vccd1 _10319_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11299_ _07013_/X fanout43/X fanout42/X _11779_/A vssd1 vssd1 vccd1 vccd1 _11300_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13038_ hold119/X _13254_/A2 _12820_/B _12642_/A vssd1 vssd1 vccd1 vccd1 hold120/A
+ sky130_fd_sc_hd__a22o_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08857__A _09673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09649__A1 _07608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07761__A _08454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11456__A1 _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07530_ _07530_/A _07530_/B vssd1 vssd1 vccd1 vccd1 _07531_/B sky130_fd_sc_hd__and2_1
XFILLER_0_76_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07461_ _07461_/A _07461_/B vssd1 vssd1 vccd1 vccd1 _07540_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12405__B1 _11637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09200_ _11242_/A reg1_val[16] _09211_/S vssd1 vssd1 vccd1 vccd1 _09200_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07392_ _09836_/A _07392_/B vssd1 vssd1 vccd1 vccd1 _07394_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12826__B _12826_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09131_ _09018_/A _09018_/B _09017_/A vssd1 vssd1 vccd1 vccd1 _09141_/A sky130_fd_sc_hd__a21bo_2
XANTENNA__13003__A _13019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09062_ _09063_/B _09063_/A vssd1 vssd1 vccd1 vccd1 _09357_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_32_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07001__A _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout206_A _08658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08013_ _08013_/A _08013_/B vssd1 vssd1 vccd1 vccd1 _08794_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__09585__B1 _07959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08927__A3 _08868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11392__B1 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09964_ _09965_/A _09965_/B vssd1 vssd1 vccd1 vccd1 _10124_/B sky130_fd_sc_hd__nor2_1
X_09895_ _09733_/X _09734_/Y _09736_/B vssd1 vssd1 vccd1 vccd1 _09899_/A sky130_fd_sc_hd__o21a_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08915_ _08917_/A _08917_/B vssd1 vssd1 vccd1 vccd1 _08915_/X sky130_fd_sc_hd__or2_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _10623_/A _08846_/B vssd1 vssd1 vccd1 vccd1 _08850_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08777_ _11809_/B _11810_/A vssd1 vssd1 vccd1 vccd1 _11893_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_95_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07728_ _07728_/A _07728_/B vssd1 vssd1 vccd1 vccd1 _07806_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_94_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07659_ _07659_/A _07659_/B vssd1 vssd1 vccd1 vccd1 _07660_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08863__A2 _09669_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout21_A _12009_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10670_ _06763_/Y _10553_/X _06765_/B vssd1 vssd1 vccd1 vccd1 _10670_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09329_ _09330_/A _09330_/B _09330_/C vssd1 vssd1 vccd1 vccd1 _09329_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_35_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06734__B _06810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09812__A1 _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09812__B2 _09943_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12340_ _12341_/A _12341_/B vssd1 vssd1 vccd1 vccd1 _12391_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_121_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12271_ _12271_/A1 _12324_/B hold282/A vssd1 vssd1 vccd1 vccd1 _12271_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11222_ _11222_/A _11222_/B vssd1 vssd1 vccd1 vccd1 _11224_/C sky130_fd_sc_hd__xor2_2
X_11153_ _11148_/Y _11149_/X _11152_/Y _11146_/X vssd1 vssd1 vccd1 vccd1 _11153_/X
+ sky130_fd_sc_hd__o211a_1
X_11084_ _11084_/A _11084_/B vssd1 vssd1 vccd1 vccd1 _11085_/B sky130_fd_sc_hd__and2_1
XFILLER_0_65_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10104_ _10104_/A _10104_/B vssd1 vssd1 vccd1 vccd1 _10105_/B sky130_fd_sc_hd__or2_1
XANTENNA__12332__C1 _12631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10035_ _09899_/A _09896_/Y _09898_/B vssd1 vssd1 vccd1 vccd1 _10039_/A sky130_fd_sc_hd__o21a_1
X_11986_ _11905_/A _11905_/B _11903_/A vssd1 vssd1 vccd1 vccd1 _11987_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_86_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10937_ _10824_/B _11050_/C _11538_/A vssd1 vssd1 vccd1 vccd1 _10937_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_14_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12607_ _12633_/A _12608_/B vssd1 vssd1 vccd1 vccd1 _12607_/X sky130_fd_sc_hd__and2_1
XFILLER_0_109_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10868_ _10868_/A _10868_/B vssd1 vssd1 vccd1 vccd1 _10869_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09301__A _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10799_ _10674_/X _10679_/X _10796_/Y _10797_/X vssd1 vssd1 vccd1 vccd1 _10800_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_30_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12538_ _12539_/A _12539_/B _12539_/C vssd1 vssd1 vccd1 vccd1 _12546_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_14_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12469_ _12469_/A _12469_/B vssd1 vssd1 vccd1 vccd1 _12470_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06961_ _11813_/S _09232_/A _09228_/B vssd1 vssd1 vccd1 vccd1 _06961_/X sky130_fd_sc_hd__or3_4
XANTENNA__09971__A _11770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09680_ _11946_/C _09680_/B vssd1 vssd1 vccd1 vccd1 _09682_/B sky130_fd_sc_hd__xnor2_2
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08700_ _07877_/A _07947_/A _07877_/C vssd1 vssd1 vccd1 vccd1 _08702_/B sky130_fd_sc_hd__a21o_1
X_06892_ instruction[3] instruction[4] vssd1 vssd1 vccd1 vccd1 _09232_/A sky130_fd_sc_hd__or2_4
X_08631_ _07038_/X _07148_/Y _07173_/Y _07030_/Y vssd1 vssd1 vccd1 vccd1 _08632_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06819__B _09728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08562_ _08575_/A _08562_/B vssd1 vssd1 vccd1 vccd1 _08593_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07513_ _10595_/A1 _08411_/B _10476_/A _10338_/B2 vssd1 vssd1 vccd1 vccd1 _07514_/B
+ sky130_fd_sc_hd__o22a_1
X_08493_ _08467_/B _08467_/C _08467_/A vssd1 vssd1 vccd1 vccd1 _08686_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_92_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout16 _07596_/Y vssd1 vssd1 vccd1 vccd1 fanout16/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_76_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout38 _07174_/X vssd1 vssd1 vccd1 vccd1 fanout38/X sky130_fd_sc_hd__buf_4
XFILLER_0_64_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout27 fanout28/X vssd1 vssd1 vccd1 vccd1 _08112_/B sky130_fd_sc_hd__buf_6
XANTENNA__08845__A2 fanout86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07444_ fanout80/X _10473_/B2 _10240_/A fanout76/X vssd1 vssd1 vccd1 vccd1 _07445_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout49 _11770_/A vssd1 vssd1 vccd1 vccd1 _09836_/A sky130_fd_sc_hd__buf_12
XFILLER_0_57_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07375_ _07443_/A _07375_/B vssd1 vssd1 vccd1 vccd1 _07376_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09114_ _08112_/B _11093_/A _10974_/A fanout25/X vssd1 vssd1 vccd1 vccd1 _09115_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_32_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09045_ _09032_/A _09032_/B _09030_/X vssd1 vssd1 vccd1 vccd1 _09146_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_103_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11365__B1 _11648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10092__A _10092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09947_ _09947_/A _09947_/B vssd1 vssd1 vccd1 vccd1 _09949_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12314__C1 _09225_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06792__B1 _06791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout69_A _09936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09878_ _06898_/C _09876_/X _09877_/Y vssd1 vssd1 vccd1 vccd1 _09878_/X sky130_fd_sc_hd__o21a_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08533__A1 _08649_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08533__B2 _08657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06729__B _06810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07832__C _07907_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08829_ _08829_/A _08829_/B vssd1 vssd1 vccd1 vccd1 _08900_/A sky130_fd_sc_hd__nor2_2
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _11840_/A _11840_/B _11840_/C _11567_/D vssd1 vssd1 vccd1 vccd1 _11841_/C
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_68_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ fanout45/X fanout12/X fanout7/X fanout47/X vssd1 vssd1 vccd1 vccd1 _11772_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _12087_/B _10722_/B vssd1 vssd1 vccd1 vccd1 _10728_/A sky130_fd_sc_hd__xnor2_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09121__A _11770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10653_ _10653_/A _10653_/B vssd1 vssd1 vccd1 vccd1 _10655_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_118_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10584_ _12157_/A _10584_/B vssd1 vssd1 vccd1 vccd1 _10588_/A sky130_fd_sc_hd__xnor2_1
X_13372_ _13392_/CLK _13372_/D vssd1 vssd1 vccd1 vccd1 hold288/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12323_ hold227/A _12447_/B1 _12370_/B _11648_/A vssd1 vssd1 vccd1 vccd1 _12323_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__07272__A1 _07195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07576__A _10092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12254_ instruction[7] _06884_/X _12253_/X vssd1 vssd1 vccd1 vccd1 _12254_/X sky130_fd_sc_hd__a21o_1
X_11205_ _11100_/A _11099_/B _11097_/Y vssd1 vssd1 vccd1 vccd1 _11217_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_102_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12185_ _12050_/A _12050_/B _12050_/C _12306_/B _11892_/A vssd1 vssd1 vccd1 vccd1
+ _12185_/X sky130_fd_sc_hd__a41o_1
XANTENNA__07024__A1 _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11136_ _11027_/A _11027_/B _11025_/A vssd1 vssd1 vccd1 vccd1 _11137_/B sky130_fd_sc_hd__o21a_1
XANTENNA__07575__A2 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11067_ _11067_/A _11067_/B vssd1 vssd1 vccd1 vccd1 _11070_/A sky130_fd_sc_hd__and2_1
XANTENNA__10730__A _11182_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10018_ _10294_/S _10018_/B vssd1 vssd1 vccd1 vccd1 _10018_/X sky130_fd_sc_hd__or2_1
XFILLER_0_25_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09730__S _11138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11969_ _11796_/X _11883_/A _11882_/A vssd1 vssd1 vccd1 vccd1 _11969_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_86_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11831__A1 _06984_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09031__A _09031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12387__A2 _11946_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07160_ _07148_/Y _07417_/B fanout42/X _07959_/A vssd1 vssd1 vccd1 vccd1 _07161_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07091_ _10243_/A _07091_/B vssd1 vssd1 vccd1 vccd1 _07092_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_54_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07263__A1 fanout86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07263__B2 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout228 _06792_/X vssd1 vssd1 vccd1 vccd1 _07117_/C sky130_fd_sc_hd__clkbuf_4
Xfanout217 _09725_/S vssd1 vssd1 vccd1 vccd1 _09727_/S sky130_fd_sc_hd__clkbuf_8
X_09801_ _11476_/A fanout28/X fanout26/X _11406_/A vssd1 vssd1 vccd1 vccd1 _09802_/B
+ sky130_fd_sc_hd__o22a_1
Xfanout206 _08658_/A vssd1 vssd1 vccd1 vccd1 _07604_/A sky130_fd_sc_hd__buf_6
XFILLER_0_10_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09732_ _12444_/B _09732_/B vssd1 vssd1 vccd1 vccd1 _09732_/X sky130_fd_sc_hd__or2_1
Xfanout239 _08502_/A vssd1 vssd1 vccd1 vccd1 _09672_/A sky130_fd_sc_hd__buf_8
XFILLER_0_5_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07993_ _09836_/A _07993_/B vssd1 vssd1 vccd1 vccd1 _08065_/C sky130_fd_sc_hd__xnor2_1
X_06944_ instruction[30] _06944_/B vssd1 vssd1 vccd1 vccd1 _06944_/X sky130_fd_sc_hd__or2_1
XANTENNA__08515__A1 _09404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07318__A2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06875_ _06868_/Y _06874_/Y _12313_/A vssd1 vssd1 vccd1 vccd1 _06875_/X sky130_fd_sc_hd__a21o_1
X_09663_ _09664_/A _09664_/B vssd1 vssd1 vccd1 vccd1 _09665_/A sky130_fd_sc_hd__or2_1
XANTENNA__08515__B2 _10245_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09594_ _12438_/A _09596_/B vssd1 vssd1 vccd1 vccd1 _09594_/X sky130_fd_sc_hd__or2_1
X_08614_ _08615_/B _08615_/C _09672_/A vssd1 vssd1 vccd1 vccd1 _08618_/A sky130_fd_sc_hd__a21o_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08545_ _08545_/A _08545_/B vssd1 vssd1 vccd1 vccd1 _08567_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_65_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08818__A2 _07417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12286__B _12335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09491__A2 _08199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08476_ _08480_/A _08480_/B vssd1 vssd1 vccd1 vccd1 _08476_/X sky130_fd_sc_hd__or2_1
XANTENNA__13024__B1 _13223_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07427_ _07428_/A _07428_/B _07428_/C vssd1 vssd1 vccd1 vccd1 _07429_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_9_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12378__A2 _11995_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07358_ _08870_/C _12779_/B _07585_/B1 vssd1 vssd1 vccd1 vccd1 _07359_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_33_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12506__S _12520_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07289_ _09341_/A _07289_/B vssd1 vssd1 vccd1 vccd1 _07373_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09028_ _09029_/B _09029_/A vssd1 vssd1 vccd1 vccd1 _09028_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_20_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold271 hold271/A vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold260 hold260/A vssd1 vssd1 vccd1 vccd1 hold260/X sky130_fd_sc_hd__buf_1
XANTENNA__07006__A1 _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold282 hold282/A vssd1 vssd1 vccd1 vccd1 hold282/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold293 hold293/A vssd1 vssd1 vccd1 vccd1 hold293/X sky130_fd_sc_hd__dlygate4sd3_1
X_12941_ _13178_/A _13179_/A _13178_/B vssd1 vssd1 vccd1 vccd1 _13184_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_99_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12872_ hold26/X hold258/A vssd1 vssd1 vccd1 vccd1 _12874_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_99_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11823_ _11650_/B _11910_/B hold268/A vssd1 vssd1 vccd1 vccd1 _11825_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__12066__A1 _12322_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11381__A _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _12087_/A fanout23/X fanout15/X _12009_/A vssd1 vssd1 vccd1 vccd1 _11755_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11685_ _11684_/B _11685_/B vssd1 vssd1 vccd1 vccd1 _11686_/B sky130_fd_sc_hd__and2b_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _10609_/A _10609_/B _10605_/X vssd1 vssd1 vccd1 vccd1 _10707_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10636_ _10636_/A _10636_/B vssd1 vssd1 vccd1 vccd1 _10638_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10725__A _10725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06922__B _12803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10567_ hold208/A _11990_/A1 _10685_/B _12205_/B1 vssd1 vssd1 vccd1 vccd1 _10567_/X
+ sky130_fd_sc_hd__a31o_1
X_13355_ _13358_/CLK hold15/X vssd1 vssd1 vccd1 vccd1 _13355_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08442__B1 _09940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13286_ _13379_/CLK _13286_/D vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__dfxtp_1
X_12306_ _12306_/A _12306_/B _12306_/C vssd1 vssd1 vccd1 vccd1 _12306_/X sky130_fd_sc_hd__and3_1
X_10498_ _10498_/A _10498_/B vssd1 vssd1 vccd1 vccd1 _10499_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12237_ _12237_/A _12237_/B vssd1 vssd1 vccd1 vccd1 _12239_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12168_ _07316_/Y _08875_/X _08990_/Y _07051_/X vssd1 vssd1 vccd1 vccd1 _12233_/D
+ sky130_fd_sc_hd__a22o_1
X_12099_ _12164_/B _12099_/B vssd1 vssd1 vccd1 vccd1 _12101_/C sky130_fd_sc_hd__and2_1
X_11119_ _10898_/A _11007_/A _11007_/B vssd1 vssd1 vccd1 vccd1 _11119_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_36_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10855__A2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06660_ reg2_val[31] _06783_/A vssd1 vssd1 vccd1 vccd1 _06660_/X sky130_fd_sc_hd__and2_1
XFILLER_0_36_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06591_ instruction[23] _06944_/B vssd1 vssd1 vccd1 vccd1 _06591_/X sky130_fd_sc_hd__or2_1
XFILLER_0_47_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12057__A1 _10049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10607__A2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09473__A2 _08877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08330_ _08598_/B _09770_/B2 _09940_/B2 _08538_/A1 vssd1 vssd1 vccd1 vccd1 _08331_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13006__B1 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08261_ _08286_/A _08286_/B _08250_/Y vssd1 vssd1 vccd1 vccd1 _08272_/B sky130_fd_sc_hd__a21boi_1
XANTENNA__07484__B2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07484__A1 _07830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07212_ _07212_/A _07212_/B _07212_/C vssd1 vssd1 vccd1 vccd1 _07213_/B sky130_fd_sc_hd__and3_1
XFILLER_0_6_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11568__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12834__B _12862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08192_ _09670_/A _08192_/B vssd1 vssd1 vccd1 vccd1 _08193_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07143_ _07143_/A _07357_/C vssd1 vssd1 vccd1 vccd1 _07143_/X sky130_fd_sc_hd__or2_1
XANTENNA_fanout119_A _07194_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07074_ _09944_/A _10072_/A _07073_/X vssd1 vssd1 vccd1 vccd1 _07074_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_42_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07787__A2 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07976_ _07966_/A _08062_/A _07996_/B vssd1 vssd1 vccd1 vccd1 _07976_/X sky130_fd_sc_hd__o21ba_1
X_06927_ _06927_/A _06927_/B _12218_/A vssd1 vssd1 vccd1 vccd1 _06933_/B sky130_fd_sc_hd__or3_4
X_09715_ _09715_/A _09715_/B vssd1 vssd1 vccd1 vccd1 _09715_/Y sky130_fd_sc_hd__nand2_1
X_09646_ _09646_/A _09646_/B vssd1 vssd1 vccd1 vccd1 _09686_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10846__A2 _07171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06858_ reg1_val[20] _07016_/A vssd1 vssd1 vccd1 vccd1 _06858_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_96_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06789_ _06790_/A _06790_/B vssd1 vssd1 vccd1 vccd1 _10014_/A sky130_fd_sc_hd__nor2_1
X_09577_ _09413_/A _09413_/B _09412_/B vssd1 vssd1 vccd1 vccd1 _09581_/A sky130_fd_sc_hd__o21a_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10059__B1 _10240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08528_ _06992_/A _10221_/B2 _09770_/B2 _08613_/A vssd1 vssd1 vccd1 vccd1 _08529_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_108_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08459_ _08485_/A _08485_/B vssd1 vssd1 vccd1 vccd1 _08497_/A sky130_fd_sc_hd__or2_1
XANTENNA__11559__B1 _11648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11470_ _10788_/A _11444_/Y _11445_/X _11469_/X _11443_/X vssd1 vssd1 vccd1 vccd1
+ _11471_/B sky130_fd_sc_hd__o311a_2
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06742__B _11038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10421_ _06773_/Y _10288_/Y _06775_/B vssd1 vssd1 vccd1 vccd1 _10421_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08975__A1 _12359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10352_ _10353_/A _10353_/B vssd1 vssd1 vccd1 vccd1 _10504_/A sky130_fd_sc_hd__nor2_1
X_13140_ hold281/A _13139_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13140_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12771__A2 _07357_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07778__A2 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13071_ _07200_/C _12826_/B hold80/X vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_21_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12022_ _12101_/A _12022_/B vssd1 vssd1 vccd1 vccd1 _12024_/B sky130_fd_sc_hd__or2_1
XFILLER_0_103_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10283_ _10661_/B _10283_/B vssd1 vssd1 vccd1 vccd1 _10581_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_88_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12924_ hold30/X hold281/X vssd1 vssd1 vccd1 vccd1 _13138_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_88_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07163__B1 _12438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12855_ _11946_/B _12863_/A2 hold25/X _13249_/A vssd1 vssd1 vccd1 vccd1 _13288_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11806_ _11965_/A _11806_/B vssd1 vssd1 vccd1 vccd1 _11807_/B sky130_fd_sc_hd__xnor2_4
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _12786_/A _12786_/B vssd1 vssd1 vccd1 vccd1 _12788_/A sky130_fd_sc_hd__nand2_2
X_11737_ _13317_/Q _11646_/B _11826_/B _11648_/A vssd1 vssd1 vccd1 vccd1 _11738_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09455__A2 _10337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11668_ _11667_/B _11668_/B vssd1 vssd1 vccd1 vccd1 _11669_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_43_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12654__B _12655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13407_ instruction[8] vssd1 vssd1 vccd1 vccd1 pred_idx[0] sky130_fd_sc_hd__buf_12
X_11599_ _11600_/A _11600_/B _11598_/Y vssd1 vssd1 vccd1 vccd1 _11698_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_113_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10619_ _10619_/A _10619_/B vssd1 vssd1 vccd1 vccd1 _10620_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09758__A3 _09738_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08415__B1 _08457_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13338_ _13358_/CLK _13338_/D vssd1 vssd1 vccd1 vccd1 hold145/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08966__A1 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08966__B2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13269_ _13365_/CLK _13269_/D vssd1 vssd1 vccd1 vccd1 hold111/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08194__A2 _08457_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07830_ _12808_/A _07830_/B vssd1 vssd1 vccd1 vccd1 _07936_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12278__A1 _12365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07761_ _08454_/A _07761_/B vssd1 vssd1 vccd1 vccd1 _07763_/B sky130_fd_sc_hd__xnor2_2
X_06712_ _06710_/Y _06724_/B1 _06783_/A reg2_val[18] vssd1 vssd1 vccd1 vccd1 _07088_/A
+ sky130_fd_sc_hd__a2bb2o_2
X_09500_ _09947_/A _09500_/B vssd1 vssd1 vccd1 vccd1 _09502_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10828__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07692_ _07752_/A _07691_/Y _07687_/Y vssd1 vssd1 vccd1 vccd1 _07703_/B sky130_fd_sc_hd__a21oi_1
X_06643_ reg1_val[27] _07049_/A vssd1 vssd1 vccd1 vccd1 _06643_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_78_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09431_ _12364_/A _08664_/A _09430_/Y vssd1 vssd1 vccd1 vccd1 _09432_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_87_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06574_ hold42/X vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__inv_2
X_09362_ _09362_/A _09362_/B vssd1 vssd1 vccd1 vccd1 _09364_/A sky130_fd_sc_hd__xnor2_4
X_08313_ _08313_/A _08313_/B vssd1 vssd1 vccd1 vccd1 _08316_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_11 reg1_val[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 reg1_val[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09293_ fanout65/X _07092_/Y _10245_/A1 fanout59/X vssd1 vssd1 vccd1 vccd1 _09294_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_44 instruction[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_33 reg2_val[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_55 reg2_val[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08244_ _09670_/A _08244_/B vssd1 vssd1 vccd1 vccd1 _08246_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10365__A _11398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08175_ _08177_/A _08177_/B vssd1 vssd1 vccd1 vccd1 _08175_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10213__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07126_ _07107_/X _12740_/B _07112_/B _07585_/B1 reg1_val[22] vssd1 vssd1 vccd1 vccd1
+ _07129_/C sky130_fd_sc_hd__o311a_1
XFILLER_0_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07057_ _07057_/A _07057_/B vssd1 vssd1 vccd1 vccd1 _07059_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06735__A3 _12719_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07959_ _07959_/A _07959_/B vssd1 vssd1 vccd1 vccd1 _07960_/B sky130_fd_sc_hd__nand2_1
X_10970_ _12087_/B _10970_/B vssd1 vssd1 vccd1 vccd1 _10972_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout51_A _07079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09629_ _09630_/A _09630_/B vssd1 vssd1 vccd1 vccd1 _09629_/X sky130_fd_sc_hd__and2_1
XANTENNA__07696__A1 _09669_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07696__B2 _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12640_ _12640_/A _12640_/B vssd1 vssd1 vccd1 vccd1 new_PC[27] sky130_fd_sc_hd__xnor2_4
XANTENNA__06737__B _07270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12571_ _12572_/A _12572_/B _12572_/C vssd1 vssd1 vccd1 vccd1 _12582_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_65_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11522_ _11522_/A _11522_/B vssd1 vssd1 vccd1 vccd1 _11524_/C sky130_fd_sc_hd__xor2_2
XANTENNA__12992__A2 _13000_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07849__A _08580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11453_ _11451_/Y _11453_/B vssd1 vssd1 vccd1 vccd1 _11454_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_18_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10404_ _10404_/A _10404_/B vssd1 vssd1 vccd1 vccd1 _10405_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11384_ _11385_/A _11385_/B vssd1 vssd1 vccd1 vccd1 _11479_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_104_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13123_ _13147_/A hold291/X vssd1 vssd1 vccd1 vccd1 _13365_/D sky130_fd_sc_hd__and2_1
XANTENNA__09070__B1 _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10335_ _10599_/A _08877_/B fanout6/X _10500_/A vssd1 vssd1 vccd1 vccd1 _10336_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10507__A1 _11779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10266_ _10265_/A _10265_/B _10267_/A vssd1 vssd1 vccd1 vccd1 _10266_/Y sky130_fd_sc_hd__o21ai_1
X_13054_ hold147/X _13094_/A2 _13101_/A2 hold150/X _13259_/A vssd1 vssd1 vccd1 vccd1
+ hold159/A sky130_fd_sc_hd__o221a_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10507__B2 _11764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12005_ _12218_/A _12001_/X _12004_/X vssd1 vssd1 vccd1 vccd1 dest_val[23] sky130_fd_sc_hd__o21ai_4
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09373__B2 _09146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10197_ _10197_/A _10197_/B vssd1 vssd1 vccd1 vccd1 _10198_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11483__A2 _07608_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12907_ _12905_/X _12907_/B vssd1 vssd1 vccd1 vccd1 _13120_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__12649__B _12650_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06647__B _06675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12838_ hold20/X _12862_/B vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__or2_1
XFILLER_0_75_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09428__A2 _12420_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12769_ _12767_/X _12769_/B vssd1 vssd1 vccd1 vccd1 _12780_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_17_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06663__A _12795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07759__A _08580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06662__A2 _06927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12196__B1 _12064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10746__B2 _08289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10746__A1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09980_ _09980_/A _09980_/B vssd1 vssd1 vccd1 vccd1 _09982_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07611__B2 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07611__A1 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08931_ _09779_/A _08931_/B vssd1 vssd1 vccd1 vccd1 _08933_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08862_ _09671_/A _08862_/B vssd1 vssd1 vccd1 vccd1 _08866_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__11171__A1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11171__B2 _11476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07914__A2 _07983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07813_ _07813_/A _07813_/B vssd1 vssd1 vccd1 vccd1 _07876_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09116__A1 _07830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08793_ _08793_/A _08793_/B _08793_/C vssd1 vssd1 vccd1 vccd1 _08794_/B sky130_fd_sc_hd__and3_1
X_07744_ _07749_/A _07749_/B _07733_/X vssd1 vssd1 vccd1 vccd1 _07816_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__09116__B2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11474__A2 _12158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07675_ _07676_/A _07676_/B vssd1 vssd1 vccd1 vccd1 _07675_/X sky130_fd_sc_hd__or2_1
X_06626_ instruction[38] _06675_/B vssd1 vssd1 vccd1 vccd1 _12708_/B sky130_fd_sc_hd__and2_4
X_09414_ _12064_/S _09413_/Y _09242_/B vssd1 vssd1 vccd1 vccd1 _09414_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_109_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13170__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12423__A1 _10159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12423__B2 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08627__B1 _08649_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09345_ _10234_/A2 fanout29/X _07274_/Y _07959_/B vssd1 vssd1 vccd1 vccd1 _09346_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12974__A2 _13257_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09276_ _09512_/B _09276_/B vssd1 vssd1 vccd1 vccd1 _09278_/C sky130_fd_sc_hd__or2_1
XFILLER_0_118_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08227_ _08227_/A _08227_/B vssd1 vssd1 vccd1 vccd1 _08278_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_105_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08158_ _08158_/A _08158_/B vssd1 vssd1 vccd1 vccd1 _08230_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07109_ reg1_val[18] reg1_val[19] _07109_/C vssd1 vssd1 vccd1 vccd1 _12740_/B sky130_fd_sc_hd__or3_4
X_08089_ _06992_/A fanout98/X fanout84/X _08613_/A vssd1 vssd1 vccd1 vccd1 _08090_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout99_A _07096_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10120_ _10120_/A _10120_/B vssd1 vssd1 vccd1 vccd1 _10121_/B sky130_fd_sc_hd__xnor2_4
X_10051_ _09993_/A _09993_/B _09994_/Y vssd1 vssd1 vccd1 vccd1 _10135_/A sky130_fd_sc_hd__a21bo_2
XFILLER_0_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10953_ _10954_/A _10954_/B vssd1 vssd1 vccd1 vccd1 _10953_/X sky130_fd_sc_hd__and2_1
XFILLER_0_97_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10673__B1 _11637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08330__A2 _09770_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10884_ _10882_/A _10882_/B _10885_/B vssd1 vssd1 vccd1 vccd1 _10884_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08963__A _10092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12623_ _12623_/A _12623_/B _12623_/C _12623_/D vssd1 vssd1 vccd1 vccd1 _12624_/B
+ sky130_fd_sc_hd__and4_2
XFILLER_0_109_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12554_ _12560_/B _12554_/B vssd1 vssd1 vccd1 vccd1 new_PC[13] sky130_fd_sc_hd__and2_4
XFILLER_0_66_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11505_ _11401_/A _11401_/B _11412_/A vssd1 vssd1 vccd1 vccd1 _11516_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12485_ reg1_val[4] curr_PC[4] _12520_/S vssd1 vssd1 vccd1 vccd1 _12487_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09794__A _09794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11436_ _11223_/Y _11330_/Y _11332_/B vssd1 vssd1 vccd1 vccd1 _11436_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_34_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11367_ _10159_/A _11249_/B _11366_/X vssd1 vssd1 vccd1 vccd1 _11367_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13106_ _13106_/A _13106_/B vssd1 vssd1 vccd1 vccd1 _13106_/X sky130_fd_sc_hd__xor2_1
X_10318_ curr_PC[7] _10448_/C vssd1 vssd1 vccd1 vccd1 _10318_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ _11298_/A _11298_/B vssd1 vssd1 vccd1 vccd1 _11302_/B sky130_fd_sc_hd__xor2_1
X_13037_ _13246_/A hold138/X vssd1 vssd1 vccd1 vccd1 hold139/A sky130_fd_sc_hd__and2_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08203__A _08454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10249_ _10249_/A _10249_/B _10249_/C vssd1 vssd1 vccd1 vccd1 _10383_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_28_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09649__A2 _07608_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08873__A _12336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09969__A _10092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07460_ _09944_/A _07460_/B vssd1 vssd1 vccd1 vccd1 _07540_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07391_ _07121_/Y fanout29/X _07282_/Y _07959_/B vssd1 vssd1 vccd1 vccd1 _07392_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09130_ _09130_/A _09130_/B vssd1 vssd1 vccd1 vccd1 _09143_/A sky130_fd_sc_hd__xor2_4
XANTENNA__07489__A _09922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09061_ _09357_/A _09061_/B vssd1 vssd1 vccd1 vccd1 _09063_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_32_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08012_ _08013_/A _08013_/B vssd1 vssd1 vccd1 vccd1 _08012_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_114_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12842__B _12862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07001__B _12644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout101_A _07088_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09585__B2 _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11392__A1 _12233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11392__B2 _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09963_ _09963_/A _09963_/B vssd1 vssd1 vccd1 vccd1 _09965_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08914_ _08914_/A _08914_/B vssd1 vssd1 vccd1 vccd1 _08917_/B sky130_fd_sc_hd__xor2_4
X_09894_ _09892_/Y _09893_/X _07117_/C _12422_/A vssd1 vssd1 vccd1 vccd1 _09894_/X
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _09661_/B2 fanout86/X fanout82/X fanout98/X vssd1 vssd1 vccd1 vccd1 _08846_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13165__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08776_ _08779_/A _08776_/B vssd1 vssd1 vccd1 vccd1 _11810_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_79_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07727_ _07751_/A _07751_/B vssd1 vssd1 vccd1 vccd1 _07806_/A sky130_fd_sc_hd__and2_1
XFILLER_0_94_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07658_ _07658_/A _07658_/B vssd1 vssd1 vccd1 vccd1 _07659_/B sky130_fd_sc_hd__xnor2_2
X_06609_ instruction[1] instruction[2] instruction[0] pred_val vssd1 vssd1 vccd1 vccd1
+ _06927_/B sky130_fd_sc_hd__and4bb_2
XFILLER_0_48_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07589_ _07589_/A _07589_/B _07589_/C vssd1 vssd1 vccd1 vccd1 _07591_/A sky130_fd_sc_hd__and3_1
XFILLER_0_48_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09328_ _09330_/A _09330_/B _09330_/C vssd1 vssd1 vccd1 vccd1 _09331_/A sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout14_A _12335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09812__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09259_ _11752_/S _09257_/X _09258_/X vssd1 vssd1 vccd1 vccd1 dest_val[0] sky130_fd_sc_hd__o21ai_4
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12270_ hold284/A _12270_/B vssd1 vssd1 vccd1 vccd1 _12324_/B sky130_fd_sc_hd__or2_1
XFILLER_0_105_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11221_ _11222_/A _11222_/B vssd1 vssd1 vccd1 vccd1 _11331_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_105_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11152_ _07270_/A _12422_/A _11151_/Y vssd1 vssd1 vccd1 vccd1 _11152_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10103_ _10104_/A _10104_/B vssd1 vssd1 vccd1 vccd1 _10105_/A sky130_fd_sc_hd__nand2_1
X_11083_ _11084_/A _11084_/B vssd1 vssd1 vccd1 vccd1 _11201_/A sky130_fd_sc_hd__nor2_1
X_10034_ _06898_/B _12420_/A0 _10033_/X vssd1 vssd1 vccd1 vccd1 _10034_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11985_ _11985_/A _11985_/B vssd1 vssd1 vccd1 vccd1 _11987_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_86_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10936_ _11159_/C _10935_/Y _10821_/A _10933_/X vssd1 vssd1 vccd1 vccd1 dest_val[12]
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_128_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10867_ _10868_/A _10868_/B vssd1 vssd1 vccd1 vccd1 _10990_/B sky130_fd_sc_hd__or2_1
XFILLER_0_39_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12606_ reg1_val[22] curr_PC[22] _12631_/S vssd1 vssd1 vccd1 vccd1 _12608_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_94_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09301__B _10476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06925__B _06926_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10798_ _10796_/Y _10797_/X _10674_/X _10679_/X vssd1 vssd1 vccd1 vccd1 _10798_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11071__B1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12537_ _12546_/A _12537_/B vssd1 vssd1 vccd1 vccd1 _12539_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_81_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12468_ _12469_/A _12469_/B vssd1 vssd1 vccd1 vccd1 _12476_/B sky130_fd_sc_hd__or2_1
XANTENNA__09728__S _09728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11419_ _11419_/A _11419_/B vssd1 vssd1 vccd1 vccd1 _11422_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_22_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06660__B _06783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10463__A _11182_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12399_ _12399_/A _12399_/B vssd1 vssd1 vccd1 vccd1 _12399_/X sky130_fd_sc_hd__and2_1
XFILLER_0_10_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06960_ _09233_/B instruction[5] _12438_/A _06960_/D vssd1 vssd1 vccd1 vccd1 _06960_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_39_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12323__B1 _11648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06891_ instruction[3] instruction[4] vssd1 vssd1 vccd1 vccd1 _06960_/D sky130_fd_sc_hd__nor2_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07772__A _08664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11294__A _12336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08630_ _08630_/A _08630_/B _08628_/Y vssd1 vssd1 vccd1 vccd1 _08638_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08561_ _08657_/B _08561_/A2 _08561_/B1 _08649_/A2 vssd1 vssd1 vccd1 vccd1 _08562_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08492_ _08495_/A _08495_/B vssd1 vssd1 vccd1 vccd1 _08492_/X sky130_fd_sc_hd__and2_1
X_07512_ _07515_/A _07515_/B vssd1 vssd1 vccd1 vccd1 _07512_/X sky130_fd_sc_hd__or2_1
Xfanout28 _07231_/X vssd1 vssd1 vccd1 vccd1 fanout28/X sky130_fd_sc_hd__buf_8
XFILLER_0_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout17 _12286_/A vssd1 vssd1 vccd1 vccd1 fanout17/X sky130_fd_sc_hd__buf_6
X_07443_ _07443_/A _07443_/B vssd1 vssd1 vccd1 vccd1 _07463_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_9_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout39 _07170_/Y vssd1 vssd1 vccd1 vccd1 _07554_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_29_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07374_ _07374_/A _07374_/B vssd1 vssd1 vccd1 vccd1 _07376_/A sky130_fd_sc_hd__or2_1
X_09113_ _08937_/A _08937_/B _08934_/A vssd1 vssd1 vccd1 vccd1 _09126_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09044_ _09044_/A _09044_/B vssd1 vssd1 vccd1 vccd1 _09147_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12064__S _12064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07018__C1 _06984_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12562__A0 _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10373__A _11179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09946_ _10479_/A _09946_/B vssd1 vssd1 vccd1 vccd1 _09947_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12865__A1 _07316_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09877_ _06898_/C _09876_/X _11637_/A vssd1 vssd1 vccd1 vccd1 _09877_/Y sky130_fd_sc_hd__a21oi_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08533__A2 _08561_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08828_ _08827_/B _08828_/B vssd1 vssd1 vccd1 vccd1 _08829_/B sky130_fd_sc_hd__and2b_1
X_08759_ _08759_/A _08759_/B _08759_/C vssd1 vssd1 vccd1 vccd1 _11345_/D sky130_fd_sc_hd__nand3_2
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _11770_/A _11770_/B vssd1 vssd1 vccd1 vccd1 _11774_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10628__B1 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _10974_/A _08877_/B fanout6/X _10871_/A vssd1 vssd1 vccd1 vccd1 _10722_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_83_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10548__A _10779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10652_ _10653_/B _10653_/A vssd1 vssd1 vccd1 vccd1 _10777_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_106_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10583_ _11093_/A _07362_/B fanout16/X _10974_/A vssd1 vssd1 vccd1 vccd1 _10584_/B
+ sky130_fd_sc_hd__o22a_1
X_13371_ _13392_/CLK _13371_/D vssd1 vssd1 vccd1 vccd1 hold279/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12322_ _12322_/A1 _12370_/B hold227/A vssd1 vssd1 vccd1 vccd1 _12322_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07857__A _10207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11379__A _11770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12253_ _06672_/D _12188_/X _12404_/S _06669_/Y vssd1 vssd1 vccd1 vccd1 _12253_/X
+ sky130_fd_sc_hd__o211a_1
X_11204_ _11204_/A _11204_/B vssd1 vssd1 vccd1 vccd1 _11219_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_50_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12184_ _12184_/A _12184_/B vssd1 vssd1 vccd1 vccd1 _12306_/B sky130_fd_sc_hd__and2_1
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11135_ _11135_/A _11135_/B vssd1 vssd1 vccd1 vccd1 _11137_/A sky130_fd_sc_hd__nand2_1
X_11066_ _11066_/A _11066_/B vssd1 vssd1 vccd1 vccd1 _11067_/B sky130_fd_sc_hd__or2_1
X_10017_ _09384_/X _09388_/X _10294_/S vssd1 vssd1 vccd1 vccd1 _10017_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11842__A _12050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11968_ _11968_/A _11968_/B vssd1 vssd1 vccd1 vccd1 _11968_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_86_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11899_ _06860_/A _11898_/X _09225_/Y vssd1 vssd1 vccd1 vccd1 _11899_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11831__A2 _09257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10919_ _12064_/S _10919_/B vssd1 vssd1 vccd1 vccd1 _10919_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_39_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11988__S _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07090_ _10243_/A _07091_/B vssd1 vssd1 vccd1 vccd1 _10350_/A sky130_fd_sc_hd__or2_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07263__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10193__A _11393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout229 _12412_/A vssd1 vssd1 vccd1 vccd1 _11820_/A sky130_fd_sc_hd__clkbuf_8
X_09800_ _09800_/A _09800_/B vssd1 vssd1 vccd1 vccd1 _09821_/A sky130_fd_sc_hd__and2_1
Xfanout207 _09670_/A vssd1 vssd1 vccd1 vccd1 _09947_/A sky130_fd_sc_hd__buf_12
Xfanout218 _07149_/A vssd1 vssd1 vccd1 vccd1 _09725_/S sky130_fd_sc_hd__clkbuf_8
X_07992_ _08065_/A _07992_/B _07992_/C vssd1 vssd1 vccd1 vccd1 _08065_/B sky130_fd_sc_hd__nand3_2
X_06943_ instruction[22] _06590_/X _06942_/X _06716_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[4]
+ sky130_fd_sc_hd__o211a_4
X_09731_ _09724_/X _09730_/X _11247_/A vssd1 vssd1 vccd1 vccd1 _09732_/B sky130_fd_sc_hd__mux2_2
XANTENNA__08598__A _09404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12847__A1 _11592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08515__A2 _08515_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13009__A _13019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06874_ _06874_/A _06874_/B vssd1 vssd1 vccd1 vccd1 _06874_/Y sky130_fd_sc_hd__nand2_1
X_09662_ _11381_/A _09662_/B vssd1 vssd1 vccd1 vccd1 _09664_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07723__B1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09593_ _09593_/A _09593_/B vssd1 vssd1 vccd1 vccd1 _09593_/X sky130_fd_sc_hd__or2_1
X_08613_ _08613_/A _08613_/B _08613_/C vssd1 vssd1 vccd1 vccd1 _08615_/C sky130_fd_sc_hd__or3_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout266_A _12796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08544_ _08554_/A _08554_/B _08537_/Y vssd1 vssd1 vccd1 vccd1 _08567_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11283__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09222__A _11813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08475_ _09670_/A _08475_/B vssd1 vssd1 vccd1 vccd1 _08480_/B sky130_fd_sc_hd__xnor2_2
X_07426_ _07426_/A _07426_/B vssd1 vssd1 vccd1 vccd1 _07428_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__11898__S _12359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07357_ reg1_val[26] reg1_val[27] _07357_/C vssd1 vssd1 vccd1 vccd1 _12779_/B sky130_fd_sc_hd__or3_4
XFILLER_0_45_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06581__A _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07288_ _07217_/Y fanout25/X _10500_/A _08112_/B vssd1 vssd1 vccd1 vccd1 _07289_/B
+ sky130_fd_sc_hd__o22a_1
X_09027_ _09027_/A _09027_/B vssd1 vssd1 vccd1 vccd1 _09029_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_103_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11338__A1 _10416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold250 hold297/A vssd1 vssd1 vccd1 vccd1 hold250/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 hold261/A vssd1 vssd1 vccd1 vccd1 hold261/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07006__A2 _12644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold283 hold283/A vssd1 vssd1 vccd1 vccd1 hold283/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 hold272/A vssd1 vssd1 vccd1 vccd1 hold272/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__11927__A _12096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold294 hold294/A vssd1 vssd1 vccd1 vccd1 hold294/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout81_A _07261_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09929_ _09797_/A _09797_/B _09800_/A vssd1 vssd1 vccd1 vccd1 _09933_/A sky130_fd_sc_hd__o21ai_1
X_12940_ hold36/X hold275/X vssd1 vssd1 vccd1 vccd1 _13178_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10849__B1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07714__B1 _07282_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12871_ _08974_/Y _12871_/A2 hold49/X _13246_/A vssd1 vssd1 vccd1 vccd1 _13296_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11822_ hold274/A _11822_/B vssd1 vssd1 vccd1 vccd1 _11910_/B sky130_fd_sc_hd__or2_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11274__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ _11567_/X _11626_/Y _11720_/B _11893_/A vssd1 vssd1 vccd1 vccd1 _11807_/A
+ sky130_fd_sc_hd__a31o_1
X_11684_ _11685_/B _11684_/B vssd1 vssd1 vccd1 vccd1 _11778_/B sky130_fd_sc_hd__and2b_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _10647_/A _10647_/B _10648_/Y vssd1 vssd1 vccd1 vccd1 _10774_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_83_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09219__B1 _11820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10635_ _10635_/A _10635_/B vssd1 vssd1 vccd1 vccd1 _10636_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_64_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12493__A _12665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13354_ _13354_/CLK _13354_/D vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10725__B _12428_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12305_ _12430_/B _12305_/B vssd1 vssd1 vccd1 vccd1 _12399_/A sky130_fd_sc_hd__xnor2_2
X_10566_ _11990_/A1 _10685_/B hold208/A vssd1 vssd1 vccd1 vccd1 _10566_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08442__B2 _08627_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08442__A1 _09669_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13285_ _13385_/CLK _13285_/D vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__dfxtp_1
X_10497_ _10498_/A _10498_/B vssd1 vssd1 vccd1 vccd1 _10634_/B sky130_fd_sc_hd__or2_1
XFILLER_0_87_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12236_ _12284_/B _12236_/B _12237_/B vssd1 vssd1 vccd1 vccd1 _12296_/A sky130_fd_sc_hd__and3_1
X_12167_ _12167_/A _12167_/B vssd1 vssd1 vccd1 vccd1 _12172_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10001__A1 _09862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11118_ _11118_/A _11118_/B vssd1 vssd1 vccd1 vccd1 _11333_/A sky130_fd_sc_hd__or2_2
XANTENNA__06756__A1 _06927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12098_ _12098_/A _12098_/B vssd1 vssd1 vccd1 vccd1 _12099_/B sky130_fd_sc_hd__or2_1
XANTENNA__12829__A1 _07232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11049_ _10821_/A _11046_/X _11047_/X _11048_/Y vssd1 vssd1 vccd1 vccd1 dest_val[13]
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_36_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07181__A1 _11134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06590_ _06911_/C _06911_/B instruction[2] vssd1 vssd1 vccd1 vccd1 _06590_/X sky130_fd_sc_hd__or3b_4
XANTENNA__06666__A _06723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13254__B2 _06577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08260_ _08315_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08286_/B sky130_fd_sc_hd__xor2_1
XANTENNA__07484__A2 _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07211_ _07212_/A _07212_/B _07212_/C vssd1 vssd1 vccd1 vccd1 _07213_/A sky130_fd_sc_hd__a21oi_2
X_08191_ _08641_/B _10595_/A1 _10338_/B2 _08627_/A2 vssd1 vssd1 vccd1 vccd1 _08192_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11568__B2 _11868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11568__A1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07142_ reg1_val[24] reg1_val[25] vssd1 vssd1 vccd1 vccd1 _07357_/C sky130_fd_sc_hd__or2_2
XFILLER_0_27_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07073_ _09947_/A _07073_/B _10243_/A vssd1 vssd1 vccd1 vccd1 _07073_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_2_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12850__B _12862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09217__A _09218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07975_ _07974_/B _07974_/C _07974_/A vssd1 vssd1 vccd1 vccd1 _07996_/B sky130_fd_sc_hd__o21ba_1
X_09714_ _09715_/A _09715_/B vssd1 vssd1 vccd1 vccd1 _09714_/X sky130_fd_sc_hd__or2_1
X_06926_ instruction[13] _06926_/B vssd1 vssd1 vccd1 vccd1 dest_pred[2] sky130_fd_sc_hd__and2_4
X_06857_ reg1_val[21] _06984_/B vssd1 vssd1 vccd1 vccd1 _06857_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_97_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09645_ _09646_/A _09646_/B vssd1 vssd1 vccd1 vccd1 _09782_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07960__A _09836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11482__A _12093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06788_ reg1_val[5] _06972_/C vssd1 vssd1 vccd1 vccd1 _06788_/Y sky130_fd_sc_hd__nand2_1
X_09576_ _09569_/X _09575_/X _11247_/A vssd1 vssd1 vccd1 vccd1 _09596_/B sky130_fd_sc_hd__mux2_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10059__B2 _12233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12453__C1 _12422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _08527_/A _08527_/B vssd1 vssd1 vccd1 vccd1 _08543_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08458_ _08502_/A _08458_/B vssd1 vssd1 vccd1 vccd1 _08485_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07409_ _07604_/A _07409_/B vssd1 vssd1 vccd1 vccd1 _07507_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10420_ _11630_/A _10420_/B _10420_/C vssd1 vssd1 vccd1 vccd1 _10420_/Y sky130_fd_sc_hd__nor3_1
X_08389_ _08540_/B _08561_/B1 _08576_/A2 _08515_/A2 vssd1 vssd1 vccd1 vccd1 _08390_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_116_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10351_ _10479_/A _10350_/Y _10349_/X vssd1 vssd1 vccd1 vccd1 _10353_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07200__A _10092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13070_ hold79/X _12805_/A _13250_/B _13345_/Q _13039_/A vssd1 vssd1 vccd1 vccd1
+ hold80/A sky130_fd_sc_hd__o221a_1
XFILLER_0_60_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10282_ _09713_/B _10278_/Y _10281_/Y vssd1 vssd1 vccd1 vccd1 _10283_/B sky130_fd_sc_hd__o21ai_4
X_12021_ _12021_/A _12021_/B vssd1 vssd1 vccd1 vccd1 _12022_/B sky130_fd_sc_hd__and2_1
XANTENNA__08031__A _08454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12923_ _13133_/A _13134_/A _13133_/B vssd1 vssd1 vccd1 vccd1 _13139_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__07163__A1 _07149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12854_ hold24/X _12862_/B vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__or2_1
XFILLER_0_96_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ _11014_/B _11801_/Y _11802_/Y _11804_/Y vssd1 vssd1 vccd1 vccd1 _11806_/B
+ sky130_fd_sc_hd__o211a_2
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ reg1_val[29] _12790_/B vssd1 vssd1 vccd1 vccd1 _12786_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_29_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11736_ _11646_/B _11826_/B _13317_/Q vssd1 vssd1 vccd1 vccd1 _11738_/A sky130_fd_sc_hd__a21oi_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11667_ _11668_/B _11667_/B vssd1 vssd1 vccd1 vccd1 _11783_/A sky130_fd_sc_hd__and2b_1
XANTENNA__10736__A _11582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11598_ _11490_/A _11490_/B _11487_/A vssd1 vssd1 vccd1 vccd1 _11598_/Y sky130_fd_sc_hd__a21oi_1
X_10618_ _10618_/A _10618_/B _10618_/C vssd1 vssd1 vccd1 vccd1 _10619_/B sky130_fd_sc_hd__and3_1
X_13406_ instruction[6] vssd1 vssd1 vccd1 vccd1 loadstore_size[1] sky130_fd_sc_hd__buf_12
XANTENNA__09612__B1 _07232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08415__B2 _08613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08415__A1 _06992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13337_ _13360_/CLK _13337_/D vssd1 vssd1 vccd1 vccd1 hold158/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10549_ _11809_/A _10549_/B _10581_/C vssd1 vssd1 vccd1 vccd1 _10549_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08966__A2 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11840__D_N _11567_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13268_ _13365_/CLK _13268_/D vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11567__A _12050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12670__B _12670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13199_ hold262/X _13198_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13199_/X sky130_fd_sc_hd__mux2_1
X_12219_ _12220_/B _12218_/Y _12631_/S _12215_/X vssd1 vssd1 vccd1 vccd1 dest_val[26]
+ sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_47_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07760_ _10595_/A1 _08484_/B _09479_/B1 _10338_/B2 vssd1 vssd1 vccd1 vccd1 _07761_/B
+ sky130_fd_sc_hd__o22a_1
X_06711_ reg2_val[18] _06783_/A _06724_/B1 _06710_/Y vssd1 vssd1 vccd1 vccd1 _07087_/A
+ sky130_fd_sc_hd__o2bb2a_4
XANTENNA__09679__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09430_ _12364_/A _08502_/A _08663_/A vssd1 vssd1 vccd1 vccd1 _09430_/Y sky130_fd_sc_hd__o21ai_1
X_07691_ _07752_/B vssd1 vssd1 vccd1 vccd1 _07691_/Y sky130_fd_sc_hd__inv_2
X_06642_ reg2_val[27] _06766_/B _06677_/B1 _06641_/Y vssd1 vssd1 vccd1 vccd1 _07049_/A
+ sky130_fd_sc_hd__o2bb2a_2
X_06573_ hold56/X vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__inv_2
X_09361_ _09361_/A _09361_/B vssd1 vssd1 vccd1 vccd1 _09362_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_87_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12986__B1 _13257_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08312_ _08347_/A _08347_/B _08301_/Y vssd1 vssd1 vccd1 vccd1 _08320_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__08103__B1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09292_ _09292_/A _09292_/B vssd1 vssd1 vccd1 vccd1 _09295_/B sky130_fd_sc_hd__xor2_1
XANTENNA_12 reg1_val[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09500__A _09947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 reg1_val[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08243_ _08641_/B _10338_/B2 _08457_/A2 _08627_/A2 vssd1 vssd1 vccd1 vccd1 _08244_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_45 instruction[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout229_A _12412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_34 reg2_val[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_56 wb_clk_i vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout131_A _07098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08174_ _08174_/A _08174_/B vssd1 vssd1 vccd1 vccd1 _08177_/B sky130_fd_sc_hd__xor2_2
X_07125_ _11584_/A vssd1 vssd1 vccd1 vccd1 _11484_/A sky130_fd_sc_hd__clkinv_4
XANTENNA__07020__A _07020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10213__B2 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10213__A1 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07056_ _07057_/A _07057_/B vssd1 vssd1 vccd1 vccd1 _07363_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_100_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07690__A _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07958_ _10092_/A _07958_/B vssd1 vssd1 vccd1 vccd1 _07962_/A sky130_fd_sc_hd__xnor2_1
X_06909_ _09234_/B _06909_/B vssd1 vssd1 vccd1 vccd1 dest_pred_val sky130_fd_sc_hd__xnor2_4
X_07889_ _07889_/A _07889_/B _07889_/C vssd1 vssd1 vccd1 vccd1 _08001_/A sky130_fd_sc_hd__or3_1
XANTENNA__13218__B2 _13223_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout44_A _07157_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09628_ _09834_/A _09628_/B vssd1 vssd1 vccd1 vccd1 _09630_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07696__A2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12426__C1 _12631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09559_ _11138_/A _10024_/B _09249_/Y vssd1 vssd1 vccd1 vccd1 _09560_/A sky130_fd_sc_hd__a21oi_2
X_12570_ _12639_/A _12570_/B vssd1 vssd1 vccd1 vccd1 _12572_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09410__A _12644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11521_ _11522_/A _11522_/B vssd1 vssd1 vccd1 vccd1 _11616_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__06656__B1 _06783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11452_ reg1_val[17] curr_PC[17] vssd1 vssd1 vccd1 vccd1 _11453_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11383_ _11582_/A _11383_/B vssd1 vssd1 vccd1 vccd1 _11385_/B sky130_fd_sc_hd__xnor2_1
X_10403_ _10401_/A _10401_/B _10404_/B vssd1 vssd1 vccd1 vccd1 _10403_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09070__A1 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10334_ _10275_/A _10275_/B _10273_/Y vssd1 vssd1 vccd1 vccd1 _10415_/A sky130_fd_sc_hd__a21boi_4
X_13122_ hold290/X _13254_/A2 _13121_/X _06577_/A vssd1 vssd1 vccd1 vccd1 hold291/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07081__B1 _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09070__B2 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10507__A2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10265_ _10265_/A _10265_/B vssd1 vssd1 vccd1 vccd1 _10267_/B sky130_fd_sc_hd__nor2_1
X_13053_ _10243_/A _12820_/B hold148/X vssd1 vssd1 vccd1 vccd1 hold149/A sky130_fd_sc_hd__a21boi_1
XANTENNA__07908__B1 _08613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12004_ _12631_/S _12004_/B _12079_/B vssd1 vssd1 vccd1 vccd1 _12004_/X sky130_fd_sc_hd__or3_1
X_10196_ _10197_/A _10197_/B vssd1 vssd1 vccd1 vccd1 _10198_/A sky130_fd_sc_hd__and2_1
XFILLER_0_17_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13209__B2 _13223_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12906_ hold256/X hold111/X vssd1 vssd1 vccd1 vccd1 _12907_/B sky130_fd_sc_hd__nand2b_1
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ _07269_/Y _12863_/A2 hold51/X _13249_/A vssd1 vssd1 vccd1 vccd1 _13279_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09833__B1 fanout72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12768_ reg1_val[26] _12790_/B vssd1 vssd1 vccd1 vccd1 _12769_/B sky130_fd_sc_hd__or2_1
XANTENNA__12665__B _12665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11719_ _11884_/A _11719_/B vssd1 vssd1 vccd1 vccd1 _11720_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_83_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06663__B _07147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12699_ _12699_/A _12699_/B _12699_/C vssd1 vssd1 vccd1 vccd1 _12700_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_127_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09597__C1 _09242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10746__A2 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07611__A2 _09669_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11297__A _11398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08930_ _07121_/Y _07417_/B fanout42/X _07134_/Y vssd1 vssd1 vccd1 vccd1 _08931_/B
+ sky130_fd_sc_hd__a22o_1
X_08861_ _07983_/A _07608_/Y _08859_/Y _12642_/A vssd1 vssd1 vccd1 vccd1 _08862_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11171__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08572__B1 _07282_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07812_ _07810_/A _07810_/B _07811_/Y vssd1 vssd1 vccd1 vccd1 _07876_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__09116__A2 _10599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08792_ _08772_/B _08772_/C _08779_/X _08791_/B vssd1 vssd1 vccd1 vccd1 _08793_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07743_ _07743_/A _07743_/B vssd1 vssd1 vccd1 vccd1 _07749_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__13017__A _13019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07674_ _07674_/A _07674_/B vssd1 vssd1 vccd1 vccd1 _07676_/B sky130_fd_sc_hd__xnor2_4
X_06625_ _06673_/A vssd1 vssd1 vccd1 vccd1 _06625_/Y sky130_fd_sc_hd__inv_2
X_09413_ _09413_/A _09413_/B vssd1 vssd1 vccd1 vccd1 _09413_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09824__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08627__A1 _09404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08627__B2 _08641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09344_ _09344_/A _09344_/B vssd1 vssd1 vccd1 vccd1 _09347_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_118_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09275_ _09274_/B _09275_/B vssd1 vssd1 vccd1 vccd1 _09276_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08226_ _08275_/A _08275_/B _08187_/X vssd1 vssd1 vccd1 vccd1 _08278_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08157_ _08157_/A _08157_/B vssd1 vssd1 vccd1 vccd1 _08158_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_15_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07108_ reg1_val[16] reg1_val[17] vssd1 vssd1 vccd1 vccd1 _07109_/C sky130_fd_sc_hd__or2_2
XFILLER_0_113_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10823__B _11050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08088_ _08088_/A _08088_/B vssd1 vssd1 vccd1 vccd1 _08119_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_113_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07039_ _08657_/B fanout59/X fanout57/X _08649_/A2 vssd1 vssd1 vccd1 vccd1 _07040_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10050_ _09998_/A _09998_/B _09996_/X vssd1 vssd1 vccd1 vccd1 _10136_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_11_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10370__B1 _10476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07118__A1 _11029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10952_ _11179_/A _10952_/B vssd1 vssd1 vccd1 vccd1 _10954_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_128_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10883_ _10741_/A _10741_/B _10740_/A vssd1 vssd1 vccd1 vccd1 _10885_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_85_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12622_ _12608_/B _12616_/B _12633_/A vssd1 vssd1 vccd1 vccd1 _12623_/D sky130_fd_sc_hd__o21ai_1
XFILLER_0_66_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12553_ _12553_/A _12553_/B _12553_/C vssd1 vssd1 vccd1 vccd1 _12554_/B sky130_fd_sc_hd__nand3_1
XANTENNA__06629__B1 _06766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11504_ _11504_/A _11504_/B vssd1 vssd1 vccd1 vccd1 _11518_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_109_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12484_ _12490_/B _12484_/B vssd1 vssd1 vccd1 vccd1 new_PC[3] sky130_fd_sc_hd__and2_4
XFILLER_0_80_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11435_ _11801_/A vssd1 vssd1 vccd1 vccd1 _11435_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11829__B _11829_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11366_ _09221_/Y _11262_/X _11364_/Y _11365_/X vssd1 vssd1 vccd1 vccd1 _11366_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07054__B1 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11297_ _11398_/A _11297_/B vssd1 vssd1 vccd1 vccd1 _11298_/B sky130_fd_sc_hd__xor2_1
X_13105_ _13147_/A hold304/X vssd1 vssd1 vccd1 vccd1 _13361_/D sky130_fd_sc_hd__and2_1
X_10317_ _12365_/A _10286_/Y _10287_/X _10316_/X _10285_/Y vssd1 vssd1 vccd1 vccd1
+ _10317_/X sky130_fd_sc_hd__a311o_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13036_ hold232/A _13248_/A2 _13248_/B1 hold137/X vssd1 vssd1 vccd1 vccd1 hold138/A
+ sky130_fd_sc_hd__a22o_1
X_10248_ _10247_/A _10247_/B _10247_/C vssd1 vssd1 vccd1 vccd1 _10249_/C sky130_fd_sc_hd__a21o_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10179_ _10179_/A _10179_/B vssd1 vssd1 vccd1 vccd1 _10179_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11580__A _11929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07390_ _10092_/A _07390_/B vssd1 vssd1 vccd1 vccd1 _07394_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09060_ _09060_/A _09060_/B _09060_/C vssd1 vssd1 vccd1 vccd1 _09061_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_114_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08011_ _08011_/A _08011_/B vssd1 vssd1 vccd1 vccd1 _08013_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_114_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12615__S _12638_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11916__B2 _09221_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09585__A2 _07149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11392__A2 _07131_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09962_ _09963_/A _09963_/B vssd1 vssd1 vccd1 vccd1 _10124_/A sky130_fd_sc_hd__and2_1
XFILLER_0_110_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08913_ _08914_/B _08914_/A vssd1 vssd1 vccd1 vccd1 _08913_/Y sky130_fd_sc_hd__nand2b_1
X_09893_ hold290/A _09425_/C _10170_/C _12416_/C1 vssd1 vssd1 vccd1 vccd1 _09893_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11755__A _12336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08844_ _08844_/A _08844_/B vssd1 vssd1 vccd1 vccd1 _08869_/A sky130_fd_sc_hd__xnor2_1
X_08775_ _08774_/A _08774_/B _11538_/B _11538_/C _08768_/Y vssd1 vssd1 vccd1 vccd1
+ _11809_/B sky130_fd_sc_hd__a2111o_1
X_07726_ _09836_/A _07726_/B vssd1 vssd1 vccd1 vccd1 _07751_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11852__B1 _08859_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07657_ _07658_/A _07658_/B vssd1 vssd1 vccd1 vccd1 _08904_/B sky130_fd_sc_hd__and2b_1
X_06608_ instruction[0] instruction[1] instruction[2] instruction[41] pred_val vssd1
+ vssd1 vccd1 vccd1 _12796_/A sky130_fd_sc_hd__o311a_4
XFILLER_0_94_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06584__A _12438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07588_ _07588_/A _11844_/A vssd1 vssd1 vccd1 vccd1 _07589_/C sky130_fd_sc_hd__or2_1
XFILLER_0_118_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09327_ _11497_/A _09327_/B vssd1 vssd1 vccd1 vccd1 _09330_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07284__B1 _07282_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09258_ curr_PC[0] _10821_/A vssd1 vssd1 vccd1 vccd1 _09258_/X sky130_fd_sc_hd__or2_1
XFILLER_0_106_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09189_ reg1_val[4] reg1_val[27] _09211_/S vssd1 vssd1 vccd1 vccd1 _09189_/X sky130_fd_sc_hd__mux2_1
X_08209_ _08269_/A _08269_/B vssd1 vssd1 vccd1 vccd1 _08270_/A sky130_fd_sc_hd__or2_1
XFILLER_0_120_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11220_ _11109_/A _11109_/B _11110_/Y vssd1 vssd1 vccd1 vccd1 _11222_/B sky130_fd_sc_hd__o21ai_2
X_11151_ _12421_/A1 _11150_/X _06738_/A vssd1 vssd1 vccd1 vccd1 _11151_/Y sky130_fd_sc_hd__a21oi_1
X_10102_ _10102_/A _10102_/B vssd1 vssd1 vccd1 vccd1 _10104_/B sky130_fd_sc_hd__xnor2_1
X_11082_ _11080_/X _11081_/Y _11179_/A vssd1 vssd1 vccd1 vccd1 _11084_/B sky130_fd_sc_hd__mux2_1
X_10033_ _06790_/A _12144_/A1 _09422_/B _06788_/Y _10032_/X vssd1 vssd1 vccd1 vccd1
+ _10033_/X sky130_fd_sc_hd__o221a_1
X_11984_ reg1_val[23] curr_PC[23] vssd1 vssd1 vccd1 vccd1 _11985_/B sky130_fd_sc_hd__or2_1
XANTENNA__11843__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10935_ curr_PC[12] _10821_/B _11752_/S vssd1 vssd1 vccd1 vccd1 _10935_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10866_ _10866_/A _10866_/B vssd1 vssd1 vccd1 vccd1 _10868_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12605_ _12611_/B _12605_/B vssd1 vssd1 vccd1 vccd1 new_PC[21] sky130_fd_sc_hd__xnor2_4
XFILLER_0_39_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11071__A1 _07013_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10797_ reg1_val[11] curr_PC[11] vssd1 vssd1 vccd1 vccd1 _10797_/X sky130_fd_sc_hd__or2_1
XFILLER_0_66_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09301__C _10476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07275__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11071__B2 _11779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12536_ _12696_/B _12536_/B vssd1 vssd1 vccd1 vccd1 _12537_/B sky130_fd_sc_hd__or2_1
XFILLER_0_26_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12467_ _12476_/A _12467_/B vssd1 vssd1 vccd1 vccd1 _12469_/B sky130_fd_sc_hd__nand2_1
X_11418_ _11416_/X _11418_/B vssd1 vssd1 vccd1 vccd1 _11419_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_1_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12398_ _12429_/B _12398_/B vssd1 vssd1 vccd1 vccd1 _12398_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11349_ _11349_/A _11349_/B vssd1 vssd1 vccd1 vccd1 _11349_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11126__A2 _11124_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13019_ _13019_/A hold220/X vssd1 vssd1 vccd1 vccd1 _13319_/D sky130_fd_sc_hd__and2_1
X_06890_ instruction[6] _06889_/Y _06881_/X vssd1 vssd1 vccd1 vccd1 _06890_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_55_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08868__B _08868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08560_ _08664_/A _08560_/B vssd1 vssd1 vccd1 vccd1 _08593_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10919__A _12064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07511_ _08334_/A _07511_/B vssd1 vssd1 vccd1 vccd1 _07515_/B sky130_fd_sc_hd__xnor2_1
X_08491_ _08491_/A _08491_/B vssd1 vssd1 vccd1 vccd1 _08495_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_92_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout18 _12009_/B vssd1 vssd1 vccd1 vccd1 _12335_/B sky130_fd_sc_hd__clkbuf_8
Xfanout29 fanout30/X vssd1 vssd1 vccd1 vccd1 fanout29/X sky130_fd_sc_hd__clkbuf_8
X_07442_ _07442_/A _07442_/B vssd1 vssd1 vccd1 vccd1 _07443_/B sky130_fd_sc_hd__and2_1
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07373_ _07373_/A _07373_/B vssd1 vssd1 vccd1 vccd1 _07374_/B sky130_fd_sc_hd__nor2_1
XANTENNA__13051__A2 _12820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09112_ _09112_/A _09112_/B vssd1 vssd1 vccd1 vccd1 _09128_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09043_ _09549_/A _08919_/X _09708_/A _09552_/B _09552_/A vssd1 vssd1 vccd1 vccd1
+ _09044_/B sky130_fd_sc_hd__o32a_1
XFILLER_0_102_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06851__B _07097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08124__A _10092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09945_ _10245_/A1 fanout17/X fanout14/X _10245_/B2 vssd1 vssd1 vccd1 vccd1 _09946_/B
+ sky130_fd_sc_hd__o22a_1
X_09876_ _12404_/S _06824_/X _09875_/Y vssd1 vssd1 vccd1 vccd1 _09876_/X sky130_fd_sc_hd__o21a_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07174__S _12093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _08828_/B _08827_/B vssd1 vssd1 vccd1 vccd1 _08829_/A sky130_fd_sc_hd__and2b_1
X_08758_ _08759_/B _08759_/C _08759_/A vssd1 vssd1 vccd1 vccd1 _11345_/C sky130_fd_sc_hd__a21o_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10628__A1 _12233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10628__B2 _08289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10829__A _11179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07709_ _07709_/A _07709_/B vssd1 vssd1 vccd1 vccd1 _07805_/B sky130_fd_sc_hd__xor2_1
X_08689_ _08689_/A _08689_/B vssd1 vssd1 vccd1 vccd1 _08766_/A sky130_fd_sc_hd__xnor2_4
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ _10720_/A _10720_/B vssd1 vssd1 vccd1 vccd1 _10741_/A sky130_fd_sc_hd__or2_1
XFILLER_0_67_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10548__B _10548_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ _10651_/A _10651_/B vssd1 vssd1 vccd1 vccd1 _10653_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12250__B1 _11892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13370_ _13398_/CLK _13370_/D vssd1 vssd1 vccd1 vccd1 hold294/A sky130_fd_sc_hd__dfxtp_1
X_10582_ _10530_/A _10530_/B _10531_/Y vssd1 vssd1 vccd1 vccd1 _10653_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12321_ hold224/A _12321_/B vssd1 vssd1 vccd1 vccd1 _12370_/B sky130_fd_sc_hd__or2_1
XFILLER_0_90_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12252_ _12306_/C _12250_/X _12251_/Y vssd1 vssd1 vccd1 vccd1 _12252_/X sky130_fd_sc_hd__o21a_1
X_11203_ _11204_/A _11204_/B vssd1 vssd1 vccd1 vccd1 _11203_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__10283__B _10283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12183_ _12299_/A _12183_/B vssd1 vssd1 vccd1 vccd1 _12306_/A sky130_fd_sc_hd__xnor2_2
X_11134_ _11134_/A curr_PC[14] vssd1 vssd1 vccd1 vccd1 _11135_/B sky130_fd_sc_hd__or2_1
X_11065_ _11066_/A _11066_/B vssd1 vssd1 vccd1 vccd1 _11067_/A sky130_fd_sc_hd__nand2_1
X_10016_ _11029_/S _10015_/Y _09251_/A vssd1 vssd1 vccd1 vccd1 _10016_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_0_116_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11967_ _11968_/B vssd1 vssd1 vccd1 vccd1 _11967_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06936__B _06944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10918_ _10915_/Y _10916_/X _10795_/X _10800_/A vssd1 vssd1 vccd1 vccd1 _10919_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_128_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11898_ _11896_/X _11897_/X _12359_/A vssd1 vssd1 vccd1 vccd1 _11898_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_73_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10849_ fanout36/X _10476_/B _10476_/C fanout34/X _12233_/B vssd1 vssd1 vccd1 vccd1
+ _10850_/B sky130_fd_sc_hd__o32a_1
XFILLER_0_109_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11044__A1 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12519_ _12525_/B _12519_/B vssd1 vssd1 vccd1 vccd1 new_PC[8] sky130_fd_sc_hd__and2_4
XANTENNA__10474__A _10748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10555__B1 _11637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08879__A _09936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout219 _10294_/S vssd1 vssd1 vccd1 vccd1 _10295_/S sky130_fd_sc_hd__buf_4
Xfanout208 _07004_/Y vssd1 vssd1 vccd1 vccd1 _09670_/A sky130_fd_sc_hd__buf_12
X_07991_ _07988_/A _07988_/B _07988_/C vssd1 vssd1 vccd1 vccd1 _07992_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06942_ instruction[29] _06944_/B vssd1 vssd1 vccd1 vccd1 _06942_/X sky130_fd_sc_hd__or2_1
X_09730_ _09726_/X _09729_/X _11138_/A vssd1 vssd1 vccd1 vccd1 _09730_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08598__B _08598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12847__A2 _12863_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10307__B1 _09422_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06873_ _06672_/D _06872_/X _06869_/X vssd1 vssd1 vccd1 vccd1 _06874_/B sky130_fd_sc_hd__a21o_1
X_09661_ fanout51/X _08199_/B fanout33/X _09661_/B2 vssd1 vssd1 vccd1 vccd1 _09662_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07723__A1 _08561_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07723__B2 _08561_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09592_ hold295/A _09425_/C _09590_/X _12416_/C1 vssd1 vssd1 vccd1 vccd1 _09593_/B
+ sky130_fd_sc_hd__a31o_1
X_08612_ _07121_/A _07121_/B _06992_/A vssd1 vssd1 vccd1 vccd1 _08615_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12848__B _12862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08543_ _08543_/A _08543_/B vssd1 vssd1 vccd1 vccd1 _08554_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11283__A1 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11283__B2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08474_ _08627_/A2 _08561_/A2 _09940_/B2 _08641_/B vssd1 vssd1 vccd1 vccd1 _08475_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_119_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13024__A2 _13171_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07425_ _07425_/A _07438_/A vssd1 vssd1 vccd1 vccd1 _07426_/B sky130_fd_sc_hd__nor2_2
XANTENNA__12232__B1 _12233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07356_ _07356_/A _07356_/B vssd1 vssd1 vccd1 vccd1 _07366_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07239__B1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07958__A _10092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07287_ _07287_/A _07287_/B vssd1 vssd1 vccd1 vccd1 _07373_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_5_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09026_ _08907_/A _08907_/B _08905_/Y vssd1 vssd1 vccd1 vccd1 _09027_/B sky130_fd_sc_hd__a21boi_4
XFILLER_0_103_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold262 hold262/A vssd1 vssd1 vccd1 vccd1 hold262/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 hold251/A vssd1 vssd1 vccd1 vccd1 hold251/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold240 hold240/A vssd1 vssd1 vccd1 vccd1 hold240/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold284 hold284/A vssd1 vssd1 vccd1 vccd1 hold284/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 hold273/A vssd1 vssd1 vccd1 vccd1 hold273/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11743__C1 _12421_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold295 hold295/A vssd1 vssd1 vccd1 vccd1 hold295/X sky130_fd_sc_hd__dlygate4sd3_1
X_09928_ _09928_/A _09928_/B vssd1 vssd1 vccd1 vccd1 _09984_/A sky130_fd_sc_hd__nor2_2
XANTENNA_fanout74_A fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10849__B2 _12233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10849__A1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09859_ _09860_/A _09860_/B vssd1 vssd1 vccd1 vccd1 _09859_/X sky130_fd_sc_hd__and2_1
XANTENNA__11943__A _12009_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12870_ hold48/X _12870_/B vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__or2_1
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _11820_/A _10695_/Y _11820_/Y _09242_/B vssd1 vssd1 vccd1 vccd1 _11821_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11274__A1 _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11274__B2 _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11752_ _11748_/X _11751_/Y _11752_/S vssd1 vssd1 vccd1 vccd1 dest_val[20] sky130_fd_sc_hd__mux2_8
XFILLER_0_28_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11683_ _12096_/A _11683_/B vssd1 vssd1 vccd1 vccd1 _11684_/B sky130_fd_sc_hd__xor2_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _11271_/A _11050_/A _11538_/A vssd1 vssd1 vccd1 vccd1 _10703_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10634_ _10634_/A _10634_/B _10634_/C vssd1 vssd1 vccd1 vccd1 _10635_/B sky130_fd_sc_hd__and3_1
XFILLER_0_125_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13353_ _13354_/CLK hold74/X vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08978__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12304_ _11719_/B _12043_/Y _12300_/X _12301_/Y _12303_/X vssd1 vssd1 vccd1 vccd1
+ _12305_/B sky130_fd_sc_hd__o311a_1
X_10565_ hold217/A _10565_/B vssd1 vssd1 vccd1 vccd1 _10685_/B sky130_fd_sc_hd__or2_1
XFILLER_0_51_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10785__B1 _12356_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08442__A2 _09770_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13284_ _13379_/CLK _13284_/D vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__dfxtp_1
X_10496_ _10634_/A _10496_/B vssd1 vssd1 vccd1 vccd1 _10498_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_51_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12235_ _12235_/A _12235_/B vssd1 vssd1 vccd1 vccd1 _12237_/B sky130_fd_sc_hd__xor2_1
XANTENNA__11734__C1 _06946_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12166_ _12167_/A _12167_/B vssd1 vssd1 vccd1 vccd1 _12239_/B sky130_fd_sc_hd__and2_1
X_11117_ _11117_/A _11117_/B _11117_/C vssd1 vssd1 vccd1 vccd1 _11118_/B sky130_fd_sc_hd__and3_1
XANTENNA__06756__A2 _06723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12097_ _12098_/A _12098_/B vssd1 vssd1 vccd1 vccd1 _12164_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09155__A0 _09218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11048_ curr_PC[13] _11159_/C _10821_/A vssd1 vssd1 vccd1 vccd1 _11048_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11853__A _12093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07181__A2 _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06666__B _12696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12999_ _13001_/A hold199/X vssd1 vssd1 vccd1 vccd1 _13309_/D sky130_fd_sc_hd__and2_1
XANTENNA__13254__A2 _13254_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13006__A2 _13171_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06682__A _06723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07210_ reg1_val[20] _07210_/B vssd1 vssd1 vccd1 vccd1 _07212_/C sky130_fd_sc_hd__xor2_2
X_08190_ _08564_/A _08190_/B vssd1 vssd1 vccd1 vccd1 _08193_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11568__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07141_ _11134_/A _11242_/A _07141_/C _07143_/A vssd1 vssd1 vccd1 vccd1 _08870_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_0_55_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06724__A2_N _06783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07072_ _07907_/B _07907_/C vssd1 vssd1 vccd1 vccd1 _07072_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_30_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07974_ _07974_/A _07974_/B _07974_/C vssd1 vssd1 vccd1 vccd1 _08064_/A sky130_fd_sc_hd__or3_1
X_09713_ _10137_/B _09713_/B vssd1 vssd1 vccd1 vccd1 _09715_/B sky130_fd_sc_hd__xnor2_2
X_06925_ instruction[12] _06926_/B vssd1 vssd1 vccd1 vccd1 dest_pred[1] sky130_fd_sc_hd__and2_4
XANTENNA__12150__C1 _12149_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06856_ _11636_/A _11632_/B _06855_/X vssd1 vssd1 vccd1 vccd1 _06856_/Y sky130_fd_sc_hd__a21oi_2
X_09644_ _09644_/A _09644_/B vssd1 vssd1 vccd1 vccd1 _09646_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_97_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06787_ reg1_val[5] _06972_/C vssd1 vssd1 vccd1 vccd1 _06790_/B sky130_fd_sc_hd__and2_1
X_09575_ _09571_/X _09574_/X _11138_/A vssd1 vssd1 vccd1 vccd1 _09575_/X sky130_fd_sc_hd__mux2_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10059__A2 _10476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08526_ _08545_/A _08545_/B vssd1 vssd1 vccd1 vccd1 _08550_/B sky130_fd_sc_hd__nor2_1
X_08457_ _06992_/A _08457_/A2 _08501_/B1 _08613_/A vssd1 vssd1 vccd1 vccd1 _08458_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12205__B1 _12205_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07408_ _09298_/B2 fanout57/X _08649_/A2 fanout63/X vssd1 vssd1 vccd1 vccd1 _07409_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_92_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08388_ _08580_/A _08388_/B vssd1 vssd1 vccd1 vccd1 _08420_/A sky130_fd_sc_hd__xnor2_1
X_07339_ _07340_/B vssd1 vssd1 vccd1 vccd1 _07339_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_103_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10350_ _10350_/A fanout8/X vssd1 vssd1 vccd1 vccd1 _10350_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_60_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07200__B _09667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10842__A _11929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10281_ _10001_/Y _10541_/A _10280_/Y vssd1 vssd1 vccd1 vccd1 _10281_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09009_ _09066_/C _09009_/B vssd1 vssd1 vccd1 vccd1 _09012_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_20_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13181__B2 _13223_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12020_ _12021_/A _12021_/B vssd1 vssd1 vccd1 vccd1 _12101_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_103_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12922_ hold46/X hold260/X vssd1 vssd1 vccd1 vccd1 _13133_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07699__B1 _09298_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07163__A2 _07959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12853_ _07013_/X _12863_/A2 hold63/X _13210_/A vssd1 vssd1 vccd1 vccd1 _13287_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11804_ _11621_/X _11966_/A _11803_/Y vssd1 vssd1 vccd1 vccd1 _11804_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ reg1_val[29] _12790_/B vssd1 vssd1 vccd1 vccd1 _12786_/A sky130_fd_sc_hd__or2_1
X_11735_ hold172/A _11735_/B vssd1 vssd1 vccd1 vccd1 _11826_/B sky130_fd_sc_hd__or2_1
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07598__A _11844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11666_ _11584_/A _07213_/A _08974_/Y _11665_/Y vssd1 vssd1 vccd1 vccd1 _11667_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_71_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13405_ instruction[5] vssd1 vssd1 vccd1 vccd1 loadstore_size[0] sky130_fd_sc_hd__buf_12
XFILLER_0_24_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11597_ _11503_/A _11503_/B _11502_/A vssd1 vssd1 vccd1 vccd1 _11603_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__12009__A _12009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10617_ _10618_/A _10618_/B _10618_/C vssd1 vssd1 vccd1 vccd1 _10619_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__09612__A1 _07554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09612__B2 _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08415__A2 _10338_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13336_ _13360_/CLK hold149/X vssd1 vssd1 vccd1 vccd1 hold147/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10548_ _10779_/A _10548_/B vssd1 vssd1 vccd1 vccd1 _10581_/C sky130_fd_sc_hd__xor2_4
XFILLER_0_24_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13267_ _13365_/CLK _13267_/D vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12218_ _12218_/A _12218_/B vssd1 vssd1 vccd1 vccd1 _12218_/Y sky130_fd_sc_hd__nand2_1
X_10479_ _10479_/A _10479_/B _10479_/C vssd1 vssd1 vccd1 vccd1 _10481_/A sky130_fd_sc_hd__nand3_1
XANTENNA__09318__A _09667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13198_ _13198_/A _13198_/B vssd1 vssd1 vccd1 vccd1 _13198_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__11567__B _11567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12149_ _12365_/A _12128_/Y _12129_/X _12148_/Y vssd1 vssd1 vccd1 vccd1 _12149_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09679__A1 _09934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06710_ _06723_/A _12655_/B vssd1 vssd1 vccd1 vccd1 _06710_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09679__B2 _09822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07690_ _10246_/A _07690_/B vssd1 vssd1 vccd1 vccd1 _07752_/B sky130_fd_sc_hd__xnor2_2
X_06641_ _06703_/A _12702_/B vssd1 vssd1 vccd1 vccd1 _06641_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06572_ hold5/X vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__inv_2
XANTENNA__08103__A1 _08561_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09360_ _09361_/A _09361_/B vssd1 vssd1 vccd1 vccd1 _09360_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_86_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09300__B1 _09669_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08311_ _08311_/A _08311_/B vssd1 vssd1 vccd1 vccd1 _08347_/B sky130_fd_sc_hd__xor2_2
XANTENNA__08103__B2 _08576_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09291_ _09292_/A _09292_/B vssd1 vssd1 vccd1 vccd1 _09467_/A sky130_fd_sc_hd__nor2_1
XANTENNA_13 reg1_val[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08242_ _08664_/A _08242_/B vssd1 vssd1 vccd1 vccd1 _08246_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_7_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_35 reg2_val[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_46 reg1_val[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_57 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_24 reg1_val[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07301__A _10749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout124_A _10209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09603__A1 _12365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08173_ _08120_/A _08120_/B _08118_/X vssd1 vssd1 vccd1 vccd1 _08174_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_27_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07020__B _07020_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10213__A2 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07124_ _07129_/A _07129_/B vssd1 vssd1 vccd1 vccd1 _11584_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_42_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07055_ _09947_/A _07055_/B vssd1 vssd1 vccd1 vccd1 _07057_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07957_ _08561_/B1 _08199_/B fanout33/X _08576_/A2 vssd1 vssd1 vccd1 vccd1 _07958_/B
+ sky130_fd_sc_hd__o22a_1
X_06908_ instruction[3] _06890_/X _06902_/X _06906_/Y _06904_/X vssd1 vssd1 vccd1
+ vccd1 _06909_/B sky130_fd_sc_hd__a221o_2
X_07888_ _07888_/A _07888_/B vssd1 vssd1 vccd1 vccd1 _07889_/C sky130_fd_sc_hd__or2_1
XANTENNA__13218__A2 _13223_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06839_ _10813_/A reg1_val[11] vssd1 vssd1 vccd1 vccd1 _06839_/X sky130_fd_sc_hd__and2b_1
X_09627_ fanout46/X _10871_/A _10974_/A _07830_/B vssd1 vssd1 vccd1 vccd1 _09628_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09558_ _10295_/S _09398_/X _09248_/B vssd1 vssd1 vccd1 vccd1 _10024_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08509_ _08527_/B vssd1 vssd1 vccd1 vccd1 _08509_/Y sky130_fd_sc_hd__inv_2
X_11520_ _11520_/A _11520_/B vssd1 vssd1 vccd1 vccd1 _11522_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_108_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09489_ fanout63/X fanout86/X fanout82/X fanout61/X vssd1 vssd1 vccd1 vccd1 _09490_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_108_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11451_ reg1_val[17] curr_PC[17] vssd1 vssd1 vccd1 vccd1 _11451_/Y sky130_fd_sc_hd__nor2_1
X_11382_ fanout26/X fanout12/X fanout8/X _07231_/X vssd1 vssd1 vccd1 vccd1 _11383_/B
+ sky130_fd_sc_hd__o22a_1
X_10402_ _10255_/A _10255_/C _10255_/B vssd1 vssd1 vccd1 vccd1 _10404_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_33_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13121_ hold256/X _13120_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13121_/X sky130_fd_sc_hd__mux2_1
X_10333_ _09868_/C _10331_/X _10332_/X _10330_/Y vssd1 vssd1 vccd1 vccd1 _10416_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_33_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07081__A1 _09943_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09070__A2 _07068_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07081__B2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10264_ _10089_/A _10089_/B _10087_/Y vssd1 vssd1 vccd1 vccd1 _10267_/A sky130_fd_sc_hd__o21ai_2
X_13052_ hold156/A _13094_/A2 _13101_/A2 hold147/X _13259_/A vssd1 vssd1 vccd1 vccd1
+ hold148/A sky130_fd_sc_hd__o221a_1
XANTENNA__07908__A1 _07080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08042__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12003_ curr_PC[22] curr_PC[23] _12003_/C vssd1 vssd1 vccd1 vccd1 _12079_/B sky130_fd_sc_hd__and3_1
X_10195_ _11582_/A _10195_/B vssd1 vssd1 vccd1 vccd1 _10197_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08030__B1 _09479_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08977__A _09672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11468__A1 _10159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13209__A2 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12905_ hold111/X hold256/X vssd1 vssd1 vccd1 vccd1 _12905_/X sky130_fd_sc_hd__and2b_1
XANTENNA__10140__A1 _09862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12836_ hold50/X _12862_/B vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__or2_1
XFILLER_0_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06944__B _06944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10747__A _11179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13123__A _13147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09833__A1 _07830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12767_ reg1_val[26] _12790_/B vssd1 vssd1 vccd1 vccd1 _12767_/X sky130_fd_sc_hd__and2_1
XANTENNA__09833__B2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11718_ _11884_/A _11719_/B vssd1 vssd1 vccd1 vccd1 _11841_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_84_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12698_ _12699_/A _12699_/B _12699_/C vssd1 vssd1 vccd1 vccd1 _12705_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_126_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11649_ hold264/A _11649_/B vssd1 vssd1 vccd1 vccd1 _11739_/B sky130_fd_sc_hd__or2_1
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13319_ _13373_/CLK _13319_/D vssd1 vssd1 vccd1 vccd1 hold219/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08860_ _08860_/A _08860_/B vssd1 vssd1 vccd1 vccd1 _08860_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08572__B2 _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07811_ _07820_/A _07820_/B vssd1 vssd1 vccd1 vccd1 _07811_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_74_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08791_ _08791_/A _08791_/B vssd1 vssd1 vccd1 vccd1 _08793_/B sky130_fd_sc_hd__or2_1
X_07742_ _07739_/B _07819_/B _07739_/A vssd1 vssd1 vccd1 vccd1 _07749_/A sky130_fd_sc_hd__o21ba_1
X_07673_ _07673_/A _07673_/B vssd1 vssd1 vccd1 vccd1 _07674_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_94_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06624_ _06622_/X _06624_/B vssd1 vssd1 vccd1 vccd1 _06673_/A sky130_fd_sc_hd__and2b_1
X_09412_ _09412_/A _09412_/B vssd1 vssd1 vccd1 vccd1 _09413_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12856__B _12870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09343_ _09343_/A _09343_/B vssd1 vssd1 vccd1 vccd1 _09344_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09824__B2 _09934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09824__A1 _07283_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08627__A2 _08627_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07835__B1 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08127__A _08664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09274_ _09275_/B _09274_/B vssd1 vssd1 vccd1 vccd1 _09512_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08225_ _08232_/A _08232_/B _08214_/X vssd1 vssd1 vccd1 vccd1 _08275_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_99_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09588__B1 _11637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08156_ _08156_/A _08156_/B vssd1 vssd1 vccd1 vccd1 _08157_/B sky130_fd_sc_hd__and2_1
XFILLER_0_16_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07107_ _11134_/A _11242_/A _07141_/C vssd1 vssd1 vccd1 vccd1 _07107_/X sky130_fd_sc_hd__or3_1
XANTENNA__10392__A _11284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08087_ _08087_/A _08185_/A vssd1 vssd1 vccd1 vccd1 _08120_/A sky130_fd_sc_hd__or2_1
XFILLER_0_30_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13136__B2 _06577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10823__C _11050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07038_ _07030_/A _07030_/B _09673_/A vssd1 vssd1 vccd1 vccd1 _07038_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_3_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10370__B2 _12233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ _08876_/A _12428_/B _12385_/B vssd1 vssd1 vccd1 vccd1 fanout6/A sky130_fd_sc_hd__o21a_1
XFILLER_0_98_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10951_ fanout75/X fanout12/X fanout8/A fanout78/X vssd1 vssd1 vccd1 vccd1 _10952_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12621_ _12621_/A _12621_/B _12621_/C _12621_/D vssd1 vssd1 vccd1 vccd1 _12623_/C
+ sky130_fd_sc_hd__or4_1
X_10882_ _10882_/A _10882_/B vssd1 vssd1 vccd1 vccd1 _10885_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_97_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11162__S _11752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09815__A1 _09302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12552_ _12553_/A _12553_/B _12553_/C vssd1 vssd1 vccd1 vccd1 _12560_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_93_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11503_ _11503_/A _11503_/B vssd1 vssd1 vccd1 vccd1 _11504_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_81_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12483_ _12483_/A _12483_/B _12483_/C vssd1 vssd1 vccd1 vccd1 _12484_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_80_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11434_ _11434_/A _11623_/B vssd1 vssd1 vccd1 vccd1 _11801_/A sky130_fd_sc_hd__and2_1
XFILLER_0_53_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11398__A _11398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07054__A1 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11365_ hold204/A _11646_/B _11461_/B _11648_/A vssd1 vssd1 vccd1 vccd1 _11365_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08251__B1 _09479_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07054__B2 _09669_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11296_ _07032_/Y _07171_/A fanout38/X _11946_/B vssd1 vssd1 vccd1 vccd1 _11297_/B
+ sky130_fd_sc_hd__a22o_1
X_10316_ _09225_/Y _10290_/X _10291_/Y _10315_/X vssd1 vssd1 vccd1 vccd1 _10316_/X
+ sky130_fd_sc_hd__a31o_1
X_13104_ _12804_/A hold303/X _13103_/X _13254_/A2 hold245/X vssd1 vssd1 vccd1 vccd1
+ hold304/A sky130_fd_sc_hd__a32o_1
XFILLER_0_0_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13035_ _13142_/A hold233/X vssd1 vssd1 vccd1 vccd1 hold234/A sky130_fd_sc_hd__and2_1
X_10247_ _10247_/A _10247_/B _10247_/C vssd1 vssd1 vccd1 vccd1 _10249_/B sky130_fd_sc_hd__nand3_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09751__B1 _09238_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10178_ _10176_/Y _10178_/B vssd1 vssd1 vccd1 vccd1 _10179_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_89_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09503__B1 _09673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12819_ _07121_/Y _13101_/B2 hold55/X _13147_/A vssd1 vssd1 vccd1 vccd1 _13270_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_56_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08010_ _08075_/A _08008_/X _07954_/Y vssd1 vssd1 vccd1 vccd1 _08013_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__07786__A _10207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09961_ _09961_/A _09961_/B vssd1 vssd1 vccd1 vccd1 _09963_/B sky130_fd_sc_hd__xor2_1
XANTENNA__13118__B2 _06577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12326__C1 _12376_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08912_ _08912_/A _08912_/B vssd1 vssd1 vccd1 vccd1 _08914_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_110_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12631__S _12631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09892_ _09425_/C _10170_/C hold290/A vssd1 vssd1 vccd1 vccd1 _09892_/Y sky130_fd_sc_hd__a21oi_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout191_A _12803_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08843_ _08844_/B vssd1 vssd1 vccd1 vccd1 _08843_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08410__A _08454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08774_ _08774_/A _08774_/B vssd1 vssd1 vccd1 vccd1 _11723_/A sky130_fd_sc_hd__and2_1
XANTENNA__07026__A _09672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07725_ _07166_/Y _07959_/B fanout29/X _07173_/Y vssd1 vssd1 vccd1 vccd1 _07726_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11852__A1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11852__B2 _07171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07656_ _08904_/A _07656_/B vssd1 vssd1 vccd1 vccd1 _07658_/B sky130_fd_sc_hd__nor2_1
X_06607_ instruction[0] instruction[2] instruction[1] pred_val vssd1 vssd1 vccd1 vccd1
+ _06607_/X sky130_fd_sc_hd__or4bb_1
XANTENNA__10387__A _11770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07587_ reg1_val[29] _07587_/B vssd1 vssd1 vccd1 vccd1 _07587_/Y sky130_fd_sc_hd__xnor2_1
X_09326_ _09677_/A _08877_/B fanout6/X _09472_/A vssd1 vssd1 vccd1 vccd1 _09327_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09257_ _12808_/A _09256_/X _09257_/S vssd1 vssd1 vccd1 vccd1 _09257_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_47_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07284__A1 _07959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08208_ _08208_/A _08208_/B vssd1 vssd1 vccd1 vccd1 _08269_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07284__B2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09188_ reg1_val[5] reg1_val[26] _09211_/S vssd1 vssd1 vccd1 vccd1 _09188_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_50_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08139_ _08580_/A _08139_/B vssd1 vssd1 vccd1 vccd1 _08217_/A sky130_fd_sc_hd__xnor2_1
X_11150_ _12420_/A0 _09422_/B _11150_/S vssd1 vssd1 vccd1 vccd1 _11150_/X sky130_fd_sc_hd__mux2_1
X_10101_ _10102_/B _10102_/A vssd1 vssd1 vccd1 vccd1 _10265_/B sky130_fd_sc_hd__and2b_1
XANTENNA__10850__A _11182_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11081_ _11081_/A fanout7/X vssd1 vssd1 vccd1 vccd1 _11081_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12541__S _12638_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10032_ _12416_/C1 _10030_/X _10031_/Y _09257_/S _06827_/B vssd1 vssd1 vccd1 vccd1
+ _10032_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_98_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_4_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13379_/CLK sky130_fd_sc_hd__clkbuf_8
X_11983_ reg1_val[23] curr_PC[23] vssd1 vssd1 vccd1 vccd1 _11985_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11843__A1 _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11843__B2 _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10934_ curr_PC[11] curr_PC[12] _10934_/C vssd1 vssd1 vccd1 vccd1 _11159_/C sky130_fd_sc_hd__and3_1
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10865_ _10866_/A _10866_/B vssd1 vssd1 vccd1 vccd1 _10990_/A sky130_fd_sc_hd__nand2_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12604_ _12611_/A _12600_/Y _12596_/A vssd1 vssd1 vccd1 vccd1 _12605_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_109_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12535_ _12696_/B _12536_/B vssd1 vssd1 vccd1 vccd1 _12546_/A sky130_fd_sc_hd__nand2_1
X_10796_ reg1_val[11] curr_PC[11] vssd1 vssd1 vccd1 vccd1 _10796_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_39_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07275__A1 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11071__A2 _07171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08472__B1 _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07275__B2 fanout72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12466_ _12645_/B _12466_/B vssd1 vssd1 vccd1 vccd1 _12467_/B sky130_fd_sc_hd__or2_1
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11417_ _11417_/A _11417_/B _11415_/Y vssd1 vssd1 vccd1 vccd1 _11418_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_112_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12017__A _12017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12397_ _12183_/B _12430_/B _12300_/C _12429_/A _12396_/X vssd1 vssd1 vccd1 vccd1
+ _12398_/B sky130_fd_sc_hd__o41a_1
X_11348_ _11349_/A _11349_/B vssd1 vssd1 vccd1 vccd1 _11348_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11279_ _11279_/A _11279_/B vssd1 vssd1 vccd1 vccd1 _11280_/B sky130_fd_sc_hd__or2_1
X_13018_ hold188/X _13171_/B2 _13209_/A2 hold219/X vssd1 vssd1 vccd1 vccd1 hold220/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12323__A2 _12447_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11591__A _11591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07510_ _08457_/A2 _08289_/B fanout75/X _10500_/A vssd1 vssd1 vccd1 vccd1 _07511_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11834__A1 _11637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08490_ _08470_/A _08470_/B _08489_/Y vssd1 vssd1 vccd1 vccd1 _08495_/A sky130_fd_sc_hd__a21bo_1
Xfanout19 _11497_/A vssd1 vssd1 vccd1 vccd1 _12087_/B sky130_fd_sc_hd__buf_6
XFILLER_0_76_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07441_ _07439_/Y _07562_/B _07436_/X vssd1 vssd1 vccd1 vccd1 _07495_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_91_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07372_ _07372_/A _07372_/B vssd1 vssd1 vccd1 vccd1 _07377_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_29_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09111_ _09111_/A _09111_/B vssd1 vssd1 vccd1 vccd1 _09112_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_115_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09042_ _09034_/A _09034_/B _08915_/X vssd1 vssd1 vccd1 vccd1 _09552_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout204_A _08658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06777__B1 _06776_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09944_ _09944_/A _09944_/B vssd1 vssd1 vccd1 vccd1 _09949_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06792__A3 _12665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09875_ _12404_/S _09875_/B vssd1 vssd1 vccd1 vccd1 _09875_/Y sky130_fd_sc_hd__nand2_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _08826_/A _08826_/B vssd1 vssd1 vccd1 vccd1 _08828_/B sky130_fd_sc_hd__xnor2_1
X_08757_ _08757_/A _08757_/B _08749_/C _08749_/A vssd1 vssd1 vccd1 vccd1 _08759_/C
+ sky130_fd_sc_hd__or4bb_2
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10628__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08688_ _08433_/B _08432_/Y _08753_/A _08403_/X vssd1 vssd1 vccd1 vccd1 _08761_/A
+ sky130_fd_sc_hd__a31o_2
X_07708_ _07708_/A _07708_/B vssd1 vssd1 vccd1 vccd1 _07805_/A sky130_fd_sc_hd__xor2_2
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07639_ _07639_/A _07639_/B vssd1 vssd1 vccd1 vccd1 _07640_/B sky130_fd_sc_hd__or2_1
X_10650_ _10651_/A _10651_/B vssd1 vssd1 vccd1 vccd1 _10777_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09309_ _09476_/B _09309_/B vssd1 vssd1 vccd1 vccd1 _09321_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_118_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10581_ _10581_/A _10581_/B _10581_/C _10453_/B vssd1 vssd1 vccd1 vccd1 _11271_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_0_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12320_ _12412_/A _12318_/X _12319_/X _06946_/X vssd1 vssd1 vccd1 vccd1 _12331_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12251_ _12306_/C _12250_/X _09150_/X vssd1 vssd1 vccd1 vccd1 _12251_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08206__B1 _10476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11202_ _11202_/A _11202_/B vssd1 vssd1 vccd1 vccd1 _11204_/B sky130_fd_sc_hd__and2_1
XFILLER_0_102_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09954__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12182_ _11890_/B _12043_/B _12302_/B _12181_/X vssd1 vssd1 vccd1 vccd1 _12183_/B
+ sky130_fd_sc_hd__a31oi_4
X_11133_ _11134_/A curr_PC[14] vssd1 vssd1 vccd1 vccd1 _11135_/A sky130_fd_sc_hd__nand2_1
X_11064_ _11582_/A _11064_/B vssd1 vssd1 vccd1 vccd1 _11066_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10316__A1 _09225_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ _11028_/S _09571_/X _11247_/C vssd1 vssd1 vccd1 vccd1 _10015_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11966_ _11966_/A _12114_/A vssd1 vssd1 vccd1 vccd1 _11968_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_86_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13018__B1 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10917_ _10795_/X _10800_/A _10915_/Y _10916_/X vssd1 vssd1 vccd1 vccd1 _10917_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11897_ _11814_/A _11811_/X _06857_/Y vssd1 vssd1 vccd1 vccd1 _11897_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_73_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10848_ _10848_/A _10848_/B vssd1 vssd1 vccd1 vccd1 _10868_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10779_ _10779_/A _10900_/A vssd1 vssd1 vccd1 vccd1 _11009_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_42_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08445__B1 _08561_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12518_ _12518_/A _12518_/B _12518_/C vssd1 vssd1 vccd1 vccd1 _12519_/B sky130_fd_sc_hd__nand3_1
XANTENNA__08870__D _12779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12449_ hold297/A _12414_/X _12449_/B1 vssd1 vssd1 vccd1 vccd1 _12449_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_42_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09945__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout209 _06961_/X vssd1 vssd1 vccd1 vccd1 _09257_/S sky130_fd_sc_hd__clkbuf_8
X_07990_ _08575_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _07992_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06941_ instruction[21] _06590_/X _06940_/X _06716_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[3]
+ sky130_fd_sc_hd__o211a_4
XFILLER_0_66_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09660_ _09794_/A _09660_/B vssd1 vssd1 vccd1 vccd1 _09664_/A sky130_fd_sc_hd__xnor2_1
X_06872_ _06672_/A _06871_/X _06870_/X vssd1 vssd1 vccd1 vccd1 _06872_/X sky130_fd_sc_hd__a21o_1
X_08611_ _08619_/A _08619_/B vssd1 vssd1 vccd1 vccd1 _08611_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07723__A2 _08112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09591_ _09425_/C _09590_/X hold295/A vssd1 vssd1 vccd1 vccd1 _09593_/A sky130_fd_sc_hd__a21oi_1
X_08542_ _08569_/A _08569_/B vssd1 vssd1 vccd1 vccd1 _08554_/A sky130_fd_sc_hd__and2b_1
XANTENNA__11283__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08473_ _08564_/A _08473_/B vssd1 vssd1 vccd1 vccd1 _08480_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_119_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout154_A _07015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07424_ _07437_/B _07424_/B vssd1 vssd1 vccd1 vccd1 _07438_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12864__B _12870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12232__A1 _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07355_ _07356_/A _07356_/B vssd1 vssd1 vccd1 vccd1 _07355_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_17_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07239__A1 _08112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07239__B2 _08501_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08987__A1 _12404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07286_ _07287_/A _07287_/B vssd1 vssd1 vccd1 vccd1 _07292_/B sky130_fd_sc_hd__and2_1
XANTENNA__11991__B1 _12205_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08135__A _08564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09025_ _09025_/A _09025_/B vssd1 vssd1 vccd1 vccd1 _09027_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold241 hold241/A vssd1 vssd1 vccd1 vccd1 hold241/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 hold230/A vssd1 vssd1 vccd1 vccd1 hold230/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 hold252/A vssd1 vssd1 vccd1 vccd1 hold252/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_40_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold274 hold274/A vssd1 vssd1 vccd1 vccd1 hold274/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 hold263/A vssd1 vssd1 vccd1 vccd1 hold263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 hold285/A vssd1 vssd1 vccd1 vccd1 hold285/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 hold296/A vssd1 vssd1 vccd1 vccd1 hold296/X sky130_fd_sc_hd__dlygate4sd3_1
X_09927_ _09926_/B _09927_/B vssd1 vssd1 vccd1 vccd1 _09928_/B sky130_fd_sc_hd__and2b_1
XANTENNA_fanout67_A fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10849__A2 _10476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09858_ _09858_/A _09858_/B vssd1 vssd1 vccd1 vccd1 _09860_/B sky130_fd_sc_hd__xnor2_2
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07714__A2 _12823_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09789_ _09790_/A _09790_/B vssd1 vssd1 vccd1 vccd1 _09789_/X sky130_fd_sc_hd__and2b_1
X_08809_ _08809_/A _08809_/B vssd1 vssd1 vccd1 vccd1 _08810_/B sky130_fd_sc_hd__or2_1
X_11820_ _11820_/A _11820_/B vssd1 vssd1 vccd1 vccd1 _11820_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_68_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11751_ _11837_/B _11751_/B vssd1 vssd1 vccd1 vccd1 _11751_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11274__A2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10702_ _11752_/S _10698_/X _10701_/X vssd1 vssd1 vccd1 vccd1 dest_val[10] sky130_fd_sc_hd__o21ai_4
X_11682_ _12169_/A fanout43/X fanout41/X _06998_/X vssd1 vssd1 vccd1 vccd1 _11683_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10633_ _10634_/A _10634_/B _10634_/C vssd1 vssd1 vccd1 vccd1 _10635_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__10234__B1 _07274_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10564_ _10561_/X _10563_/X _11820_/A vssd1 vssd1 vccd1 vccd1 _10564_/X sky130_fd_sc_hd__mux2_1
X_13352_ _13354_/CLK hold110/X vssd1 vssd1 vccd1 vccd1 hold108/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08978__A1 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12303_ _12180_/Y _12302_/Y _12300_/C vssd1 vssd1 vccd1 vccd1 _12303_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_36_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08045__A _08575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13283_ _13379_/CLK _13283_/D vssd1 vssd1 vccd1 vccd1 hold121/A sky130_fd_sc_hd__dfxtp_1
X_10495_ _10494_/B _10495_/B vssd1 vssd1 vccd1 vccd1 _10496_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__09575__S _11138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12234_ _12335_/B _12234_/B _12233_/X vssd1 vssd1 vccd1 vccd1 _12235_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_32_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12165_ _12239_/A _12165_/B vssd1 vssd1 vccd1 vccd1 _12167_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_31_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11116_ _11117_/A _11117_/B _11117_/C vssd1 vssd1 vccd1 vccd1 _11118_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__06756__A3 _12696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12096_ _12096_/A _12096_/B vssd1 vssd1 vccd1 vccd1 _12098_/B sky130_fd_sc_hd__xor2_1
X_11047_ curr_PC[13] _11159_/C vssd1 vssd1 vccd1 vccd1 _11047_/X sky130_fd_sc_hd__or2_1
X_12998_ hold185/X _13000_/A2 _13257_/A2 hold169/X vssd1 vssd1 vccd1 vccd1 hold199/A
+ sky130_fd_sc_hd__a22o_1
X_11949_ _11950_/A _11950_/B vssd1 vssd1 vccd1 vccd1 _12027_/B sky130_fd_sc_hd__and2b_1
XANTENNA__10473__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06963__A _12438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12684__B _12685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06682__B _12675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07140_ reg1_val[23] _12740_/B _07140_/C vssd1 vssd1 vccd1 vccd1 _07143_/A sky130_fd_sc_hd__or3_2
XFILLER_0_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09091__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07071_ _07907_/B _07907_/C vssd1 vssd1 vccd1 vccd1 _11764_/A sky130_fd_sc_hd__and2_4
XFILLER_0_112_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09712_ _09039_/B _09708_/X _09710_/X _09711_/X vssd1 vssd1 vccd1 vccd1 _09713_/B
+ sky130_fd_sc_hd__o211a_2
X_07973_ _07970_/A _07970_/B _07970_/C vssd1 vssd1 vccd1 vccd1 _07974_/C sky130_fd_sc_hd__a21oi_2
XFILLER_0_93_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06924_ instruction[11] _06926_/B vssd1 vssd1 vccd1 vccd1 dest_pred[0] sky130_fd_sc_hd__and2_4
X_06855_ reg1_val[19] _07078_/A vssd1 vssd1 vccd1 vccd1 _06855_/X sky130_fd_sc_hd__and2_1
X_09643_ _09644_/A _09644_/B vssd1 vssd1 vccd1 vccd1 _09782_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09514__A _11284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06857__B _06984_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09574_ _09572_/X _09573_/X _10295_/S vssd1 vssd1 vccd1 vccd1 _09574_/X sky130_fd_sc_hd__mux2_1
X_06786_ reg1_val[5] _06972_/C vssd1 vssd1 vccd1 vccd1 _06790_/A sky130_fd_sc_hd__nor2_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08525_ _08525_/A _08525_/B vssd1 vssd1 vccd1 vccd1 _08545_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10059__A3 _10476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08456_ _08575_/A _08456_/B vssd1 vssd1 vccd1 vccd1 _08485_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07407_ _09672_/A _07407_/B vssd1 vssd1 vccd1 vccd1 _07507_/A sky130_fd_sc_hd__xnor2_1
X_08387_ _08538_/A1 _08561_/A2 _09940_/B2 _08598_/B vssd1 vssd1 vccd1 vccd1 _08388_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08409__B1 _09479_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07338_ _10479_/A _07338_/B vssd1 vssd1 vccd1 vccd1 _07340_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_122_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09082__B1 _11198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07269_ _07270_/A _07270_/B vssd1 vssd1 vccd1 vccd1 _07269_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_61_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10280_ _10136_/A _10136_/B _10279_/X vssd1 vssd1 vccd1 vccd1 _10280_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09008_ _09008_/A _09008_/B vssd1 vssd1 vccd1 vccd1 _09009_/B sky130_fd_sc_hd__nor2_1
XANTENNA__13181__A2 _13223_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07396__B1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12921_ _13128_/A _13129_/A _13128_/B vssd1 vssd1 vccd1 vccd1 _13134_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__07699__A1 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07699__B2 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12852_ hold62/X _12862_/B vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__or2_1
X_11803_ _11617_/A _11710_/A _11710_/B vssd1 vssd1 vccd1 vccd1 _11803_/Y sky130_fd_sc_hd__a21boi_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _12787_/B _12783_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[28] sky130_fd_sc_hd__nor2_8
XANTENNA__06783__A _06783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11734_ _11820_/A _11732_/X _11733_/Y _06946_/X vssd1 vssd1 vccd1 vccd1 _11747_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07320__B1 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11665_ _07218_/X _08974_/Y _11584_/A vssd1 vssd1 vccd1 vccd1 _11665_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13404_ instruction[16] vssd1 vssd1 vccd1 vccd1 loadstore_dest[5] sky130_fd_sc_hd__buf_12
X_10616_ _10616_/A _10707_/A vssd1 vssd1 vccd1 vccd1 _10618_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11596_ _11504_/A _11504_/B _11493_/A vssd1 vssd1 vccd1 vccd1 _11609_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__12009__B _12009_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09612__A2 _10725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13335_ _13360_/CLK _13335_/D vssd1 vssd1 vccd1 vccd1 hold156/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10547_ _10003_/X _10541_/X _10543_/Y max_cap4/X _10546_/X vssd1 vssd1 vccd1 vccd1
+ _10548_/B sky130_fd_sc_hd__a221oi_4
XFILLER_0_122_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10478_ _10623_/A _10478_/B _10478_/C vssd1 vssd1 vccd1 vccd1 _10479_/C sky130_fd_sc_hd__nand3_1
X_13266_ _13365_/CLK _13266_/D vssd1 vssd1 vccd1 vccd1 hold154/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12217_ curr_PC[24] curr_PC[25] _12079_/B curr_PC[26] vssd1 vssd1 vccd1 vccd1 _12218_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13197_ _13210_/A hold263/X vssd1 vssd1 vccd1 vccd1 _13380_/D sky130_fd_sc_hd__and2_1
XFILLER_0_20_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12148_ _09242_/B _12135_/X _12147_/X vssd1 vssd1 vccd1 vccd1 _12148_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_47_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06958__A _06958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12079_ curr_PC[24] _12079_/B vssd1 vssd1 vccd1 vccd1 _12216_/C sky130_fd_sc_hd__and2_1
XANTENNA__09679__A2 _08877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12679__B _12680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06640_ instruction[37] _06675_/B vssd1 vssd1 vccd1 vccd1 _12702_/B sky130_fd_sc_hd__and2_4
XANTENNA__10694__B1 _10692_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08887__B1 _07238_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06571_ hold296/X vssd1 vssd1 vccd1 vccd1 _06571_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_59_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12986__A2 _13000_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09300__A1 _07608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08310_ _08306_/A _08306_/B _08309_/Y vssd1 vssd1 vccd1 vccd1 _08347_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__08103__A2 _08289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09290_ _10749_/A _09290_/B vssd1 vssd1 vccd1 vccd1 _09292_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_14 reg1_val[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08241_ _06992_/A fanout80/X fanout76/X _08613_/A vssd1 vssd1 vccd1 vccd1 _08242_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07311__B1 _08649_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_36 reg2_val[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_47 reg1_val[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 reg1_val[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_58 reg1_val[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08172_ _08172_/A _08172_/B vssd1 vssd1 vccd1 vccd1 _08174_/A sky130_fd_sc_hd__xor2_2
X_07123_ reg1_val[20] _07585_/B1 _07210_/B reg1_val[21] vssd1 vssd1 vccd1 vccd1 _07129_/B
+ sky130_fd_sc_hd__a211oi_4
XANTENNA_fanout117_A _07198_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07054_ fanout63/X _09301_/A fanout57/X _09669_/B2 vssd1 vssd1 vccd1 vccd1 _07055_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10154__S _12054_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07378__B1 _10240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07029__A _08502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07956_ _07956_/A _07956_/B vssd1 vssd1 vccd1 vccd1 _08006_/A sky130_fd_sc_hd__xnor2_2
X_06907_ _06949_/A instruction[4] vssd1 vssd1 vccd1 vccd1 _09234_/C sky130_fd_sc_hd__or2_2
X_07887_ _07853_/B _07887_/B vssd1 vssd1 vccd1 vccd1 _07888_/B sky130_fd_sc_hd__and2b_1
XANTENNA__08878__B1 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06838_ _10672_/A _06836_/Y _06837_/X vssd1 vssd1 vccd1 vccd1 _06838_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_0_69_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09626_ _11582_/A _09626_/B vssd1 vssd1 vccd1 vccd1 _09630_/A sky130_fd_sc_hd__xnor2_2
X_06769_ reg1_val[8] _07215_/A vssd1 vssd1 vccd1 vccd1 _06770_/B sky130_fd_sc_hd__nand2_1
X_09557_ _08664_/B _08715_/B _09557_/S vssd1 vssd1 vccd1 vccd1 _09557_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_93_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10437__B1 _11554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09488_ _09488_/A _09488_/B vssd1 vssd1 vccd1 vccd1 _09508_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08508_ _08658_/A _08508_/B vssd1 vssd1 vccd1 vccd1 _08527_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07302__B1 fanout72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08439_ _08465_/A _08465_/B vssd1 vssd1 vccd1 vccd1 _08467_/B sky130_fd_sc_hd__or2_1
XFILLER_0_93_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11450_ _11354_/A _11351_/Y _11353_/B vssd1 vssd1 vccd1 vccd1 _11454_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_80_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11381_ _11381_/A _11381_/B vssd1 vssd1 vccd1 vccd1 _11385_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10401_ _10401_/A _10401_/B vssd1 vssd1 vccd1 vccd1 _10404_/A sky130_fd_sc_hd__or2_1
XFILLER_0_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13120_ _13120_/A _13120_/B vssd1 vssd1 vccd1 vccd1 _13120_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__09419__A _12054_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10332_ _09044_/A _09044_/B _09863_/X _10331_/X vssd1 vssd1 vccd1 vccd1 _10332_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_33_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07081__A2 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13051_ _07073_/B _12820_/B hold157/X vssd1 vssd1 vccd1 vccd1 _13335_/D sky130_fd_sc_hd__a21boi_1
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12002_ curr_PC[22] _12003_/C curr_PC[23] vssd1 vssd1 vccd1 vccd1 _12004_/B sky130_fd_sc_hd__a21oi_1
X_10263_ _10118_/A _10118_/B _10119_/Y vssd1 vssd1 vccd1 vccd1 _10268_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__07908__A2 _07080_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ fanout62/X fanout28/X fanout26/X _11671_/A vssd1 vssd1 vccd1 vccd1 _10195_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08030__B2 _10221_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08030__A1 _08501_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12904_ _12902_/X _12904_/B vssd1 vssd1 vccd1 vccd1 _13124_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__07541__B1 _12823_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12835_ _07274_/Y _12863_/A2 hold107/X _13249_/A vssd1 vssd1 vccd1 vccd1 _13278_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09833__A2 _11093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12766_ _12766_/A _12770_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[25] sky130_fd_sc_hd__xnor2_4
X_11717_ _10904_/B _11334_/X _11713_/Y _11715_/X _11716_/Y vssd1 vssd1 vccd1 vccd1
+ _11719_/B sky130_fd_sc_hd__a311oi_4
XFILLER_0_84_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12697_ _12705_/A _12697_/B vssd1 vssd1 vccd1 vccd1 _12699_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11648_ _11648_/A _11648_/B _11648_/C vssd1 vssd1 vccd1 vccd1 _11657_/B sky130_fd_sc_hd__or3_1
XFILLER_0_52_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11579_ fanout45/X fanout17/X fanout14/X fanout47/X vssd1 vssd1 vccd1 vccd1 _11580_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09597__A1 _12064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13318_ _13373_/CLK hold190/X vssd1 vssd1 vccd1 vccd1 hold188/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13249_ _13249_/A hold176/X vssd1 vssd1 vccd1 vccd1 _13392_/D sky130_fd_sc_hd__and2_1
XANTENNA__11156__A1 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11156__B2 _10159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10903__A1 _10416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08572__A2 _07121_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07810_ _07810_/A _07810_/B vssd1 vssd1 vccd1 vccd1 _07820_/B sky130_fd_sc_hd__xor2_1
X_08790_ _08790_/A _08790_/B vssd1 vssd1 vccd1 vccd1 _08791_/B sky130_fd_sc_hd__or2_1
X_07741_ _07741_/A _07741_/B vssd1 vssd1 vccd1 vccd1 _07819_/B sky130_fd_sc_hd__or2_1
XANTENNA__11459__A2 _11995_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07672_ _07673_/A _07673_/B vssd1 vssd1 vccd1 vccd1 _07672_/X sky130_fd_sc_hd__and2_1
X_06623_ reg1_val[29] _08973_/A vssd1 vssd1 vccd1 vccd1 _06624_/B sky130_fd_sc_hd__or2_1
X_09411_ _12644_/A curr_PC[1] vssd1 vssd1 vccd1 vccd1 _09412_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09342_ _09343_/A _09343_/B vssd1 vssd1 vccd1 vccd1 _09344_/A sky130_fd_sc_hd__and2_1
XANTENNA__13081__A1 _11584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09824__A2 _08877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07312__A _07604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout234_A _09423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07835__B2 _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07835__A1 _09669_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09273_ _09779_/A _09273_/B vssd1 vssd1 vccd1 vccd1 _09274_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_74_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08224_ _08224_/A _08224_/B vssd1 vssd1 vccd1 vccd1 _08232_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_117_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11769__A _12093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08155_ _08155_/A _08155_/B vssd1 vssd1 vccd1 vccd1 _08158_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_99_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06870__B _06998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07106_ reg1_val[11] reg1_val[12] reg1_val[13] _07248_/B vssd1 vssd1 vccd1 vccd1
+ _07141_/C sky130_fd_sc_hd__or4_4
XFILLER_0_15_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08086_ _08087_/A _08086_/B _08086_/C vssd1 vssd1 vccd1 vccd1 _08185_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_101_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13136__A2 _13254_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07037_ _07031_/A _07031_/B _09673_/A vssd1 vssd1 vccd1 vccd1 _07037_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13195__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09760__A1 _12356_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10370__A2 _10476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08988_ _12438_/A _08985_/B _11844_/A reg1_val[30] _12795_/A vssd1 vssd1 vccd1 vccd1
+ _12385_/B sky130_fd_sc_hd__a2111o_1
XANTENNA__07771__B1 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07939_ _08014_/A _08014_/B vssd1 vssd1 vccd1 vccd1 _08015_/A sky130_fd_sc_hd__or2_1
X_10950_ _10950_/A _10950_/B vssd1 vssd1 vccd1 vccd1 _10954_/A sky130_fd_sc_hd__xnor2_2
X_10881_ _10756_/A _10756_/B _10754_/X vssd1 vssd1 vccd1 vccd1 _10886_/A sky130_fd_sc_hd__a21o_1
X_09609_ _09770_/B2 _07362_/B fanout16/X _07283_/X vssd1 vssd1 vccd1 vccd1 _09610_/B
+ sky130_fd_sc_hd__o22a_1
X_12620_ _12639_/A _12620_/B vssd1 vssd1 vccd1 vccd1 _12624_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_109_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12551_ _12560_/A _12551_/B vssd1 vssd1 vccd1 vccd1 _12553_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11502_ _11502_/A _11502_/B vssd1 vssd1 vccd1 vccd1 _11503_/B sky130_fd_sc_hd__nand2_1
X_12482_ _12483_/A _12483_/B _12483_/C vssd1 vssd1 vccd1 vccd1 _12490_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_65_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11679__A _12093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11433_ _11433_/A _11526_/A vssd1 vssd1 vccd1 vccd1 _11623_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_46_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11364_ _11646_/B _11461_/B hold204/A vssd1 vssd1 vccd1 vccd1 _11364_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07054__A2 _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08251__B2 _08561_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08251__A1 _08561_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08053__A _09341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11295_ _11298_/A vssd1 vssd1 vccd1 vccd1 _11295_/Y sky130_fd_sc_hd__inv_2
X_10315_ _12379_/B2 _10293_/X _10299_/X _09887_/X _10314_/X vssd1 vssd1 vccd1 vccd1
+ _10315_/X sky130_fd_sc_hd__a221o_1
X_13103_ hold11/X fanout2/X hold16/X vssd1 vssd1 vccd1 vccd1 _13103_/X sky130_fd_sc_hd__a21o_1
X_13034_ hold241/A _13248_/A2 _13248_/B1 hold232/X vssd1 vssd1 vccd1 vccd1 hold233/A
+ sky130_fd_sc_hd__a22o_1
X_10246_ _10246_/A _10246_/B vssd1 vssd1 vccd1 vccd1 _10247_/C sky130_fd_sc_hd__xor2_2
XANTENNA__09200__A0 _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07892__A _10092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_4_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10177_ reg1_val[6] curr_PC[6] vssd1 vssd1 vccd1 vccd1 _10178_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_28_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11310__A1 _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06677__A2_N _06766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12818_ hold54/X _12820_/B vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__or2_1
XANTENNA__09267__B1 _07238_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ reg1_val[22] _12755_/B vssd1 vssd1 vccd1 vccd1 _12751_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06971__A _07165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11589__A _11946_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10493__A _12224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11377__A1 _12050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09960_ _09960_/A _09960_/B vssd1 vssd1 vccd1 vccd1 _09961_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__13118__A2 _13254_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08911_ _08911_/A _08911_/B vssd1 vssd1 vccd1 vccd1 _08912_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_85_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09891_ hold256/A hold295/A hold235/A hold245/A vssd1 vssd1 vccd1 vccd1 _10170_/C
+ sky130_fd_sc_hd__or4_2
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08842_ _10479_/A _08842_/B vssd1 vssd1 vccd1 vccd1 _08844_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ _08772_/B _08772_/C _08779_/B vssd1 vssd1 vccd1 vccd1 _08774_/B sky130_fd_sc_hd__a21o_1
X_07724_ _09341_/A _07724_/B vssd1 vssd1 vccd1 vccd1 _07751_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07655_ _07655_/A _07655_/B _07655_/C vssd1 vssd1 vccd1 vccd1 _07656_/B sky130_fd_sc_hd__and3_1
X_06606_ instruction[0] instruction[2] instruction[1] pred_val vssd1 vssd1 vccd1 vccd1
+ _06606_/X sky130_fd_sc_hd__and4bb_1
XANTENNA__11852__A2 _07608_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07586_ reg1_val[29] _07587_/B vssd1 vssd1 vccd1 vccd1 _11844_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_48_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09325_ _09325_/A _11497_/A vssd1 vssd1 vccd1 vccd1 _09332_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_118_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10812__B1 _12416_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09256_ _09148_/Y _09151_/X _09255_/X vssd1 vssd1 vccd1 vccd1 _09256_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_47_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07284__A2 _12823_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11499__A _12096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08207_ _10207_/A _08207_/B vssd1 vssd1 vccd1 vccd1 _08269_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11368__A1 _06946_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09187_ _09185_/X _09186_/X _09403_/S vssd1 vssd1 vccd1 vccd1 _09187_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08138_ _08598_/B _10338_/B2 _08457_/A2 _08538_/A1 vssd1 vssd1 vccd1 vccd1 _08139_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10040__A1 _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08069_ _08068_/A _08079_/A vssd1 vssd1 vccd1 vccd1 _08170_/A sky130_fd_sc_hd__and2b_1
XANTENNA__11946__B _11946_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11080_ _11080_/A fanout7/X vssd1 vssd1 vccd1 vccd1 _11080_/X sky130_fd_sc_hd__or2_1
X_10100_ _10100_/A _10100_/B vssd1 vssd1 vccd1 vccd1 _10102_/B sky130_fd_sc_hd__xnor2_1
X_10031_ hold248/A _10031_/B vssd1 vssd1 vccd1 vccd1 _10031_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11982_ _06700_/A _11980_/X _11981_/Y vssd1 vssd1 vccd1 vccd1 _11982_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_105_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11843__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10933_ _10933_/A _10933_/B _10933_/C _10933_/D vssd1 vssd1 vccd1 vccd1 _10933_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10864_ _10864_/A _10864_/B vssd1 vssd1 vccd1 vccd1 _10866_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_85_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13045__A1 _09673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12603_ _12633_/A _12603_/B vssd1 vssd1 vccd1 vccd1 _12611_/B sky130_fd_sc_hd__xnor2_4
X_10795_ reg1_val[11] curr_PC[11] vssd1 vssd1 vccd1 vccd1 _10795_/X sky130_fd_sc_hd__and2_1
XFILLER_0_39_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12534_ reg1_val[11] curr_PC[11] _12638_/S vssd1 vssd1 vccd1 vccd1 _12536_/B sky130_fd_sc_hd__mux2_1
XANTENNA__08472__A1 _08515_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07275__A2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08472__B2 _08540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12465_ _12645_/B _12466_/B vssd1 vssd1 vccd1 vccd1 _12476_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07098__S _10479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11416_ _11417_/A _11417_/B _11415_/Y vssd1 vssd1 vccd1 vccd1 _11416_/X sky130_fd_sc_hd__o21ba_1
X_12396_ _12430_/B _12301_/Y _12429_/A _12395_/X vssd1 vssd1 vccd1 vccd1 _12396_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11347_ _06848_/X _11346_/X _11813_/S vssd1 vssd1 vccd1 vccd1 _11349_/B sky130_fd_sc_hd__mux2_1
XANTENNA__12308__B1 _09150_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12859__A1 _06998_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11278_ _11279_/A _11279_/B vssd1 vssd1 vccd1 vccd1 _11389_/A sky130_fd_sc_hd__nand2_1
X_13017_ _13019_/A hold189/X vssd1 vssd1 vccd1 vccd1 hold190/A sky130_fd_sc_hd__and2_1
X_10229_ _11844_/A _10229_/B vssd1 vssd1 vccd1 vccd1 _10233_/A sky130_fd_sc_hd__xnor2_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06966__A _12644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06685__B _07014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07440_ _07440_/A _07440_/B vssd1 vssd1 vccd1 vccd1 _07562_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_29_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07371_ _07371_/A _07371_/B vssd1 vssd1 vccd1 vccd1 _07372_/B sky130_fd_sc_hd__or2_1
XFILLER_0_72_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09110_ _09111_/A _09111_/B vssd1 vssd1 vccd1 vccd1 _09110_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_29_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09041_ _08807_/B _08807_/C _09549_/A _08920_/X _09708_/A vssd1 vssd1 vccd1 vccd1
+ _09044_/A sky130_fd_sc_hd__a2111o_1
XFILLER_0_17_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09943_ _09650_/A fanout13/X fanout8/X _09943_/B2 vssd1 vssd1 vccd1 vccd1 _09944_/B
+ sky130_fd_sc_hd__o22a_1
X_09874_ _06800_/Y _09743_/B _09743_/C _06802_/B vssd1 vssd1 vccd1 vccd1 _09875_/B
+ sky130_fd_sc_hd__o31ai_2
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08825_ _08825_/A _08825_/B vssd1 vssd1 vccd1 vccd1 _08826_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09479__B1 _09479_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08756_ _08434_/A _08434_/B _08755_/X vssd1 vssd1 vccd1 vccd1 _08759_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__06595__B _06944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08687_ _08757_/A _08687_/B _08687_/C vssd1 vssd1 vccd1 vccd1 _08753_/A sky130_fd_sc_hd__or3_2
X_07707_ _07709_/A _07709_/B vssd1 vssd1 vccd1 vccd1 _07707_/Y sky130_fd_sc_hd__nor2_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07638_ _07639_/A _07639_/B vssd1 vssd1 vccd1 vccd1 _08893_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_48_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07569_ _07679_/B _07679_/A vssd1 vssd1 vccd1 vccd1 _07569_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_118_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09398__S _09728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09308_ _09307_/B _09307_/C _09307_/A vssd1 vssd1 vccd1 vccd1 _09309_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout12_A fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09651__B1 _09944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10580_ _12471_/S _10452_/X _10579_/X vssd1 vssd1 vccd1 vccd1 dest_val[9] sky130_fd_sc_hd__o21a_4
XFILLER_0_35_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09239_ _09239_/A _09239_/B vssd1 vssd1 vccd1 vccd1 _09239_/X sky130_fd_sc_hd__or2_1
XFILLER_0_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12250_ _12050_/X _12306_/A _12306_/B _11892_/A vssd1 vssd1 vccd1 vccd1 _12250_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08206__A1 _08561_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08206__B2 _08576_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11201_ _11201_/A _11201_/B vssd1 vssd1 vccd1 vccd1 _11202_/B sky130_fd_sc_hd__nand2_1
X_12181_ _12044_/Y _12302_/B _12180_/Y vssd1 vssd1 vccd1 vccd1 _12181_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__10013__A1 _12438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09954__A1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09954__B2 _11868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11132_ _11131_/A _11131_/B _11131_/Y _09225_/Y vssd1 vssd1 vccd1 vccd1 _11157_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08331__A _08580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11063_ _12233_/B fanout26/X fanout17/X fanout28/X vssd1 vssd1 vccd1 vccd1 _11064_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09146__B _09146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10014_ _10014_/A _10014_/B vssd1 vssd1 vccd1 vccd1 _10014_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11965_ _11965_/A _12042_/A vssd1 vssd1 vccd1 vccd1 _12114_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_59_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10916_ reg1_val[12] curr_PC[12] vssd1 vssd1 vccd1 vccd1 _10916_/X sky130_fd_sc_hd__or2_1
X_11896_ _11814_/A _11812_/X _11829_/A vssd1 vssd1 vccd1 vccd1 _11896_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__06705__A_N _07078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09890__B1 _12205_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10847_ _12093_/A _10847_/B vssd1 vssd1 vccd1 vccd1 _10848_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_109_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10778_ _10778_/A _10778_/B vssd1 vssd1 vccd1 vccd1 _11008_/A sky130_fd_sc_hd__or2_4
XFILLER_0_54_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08445__B2 _08538_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08445__A1 _08598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12517_ _12518_/A _12518_/B _12518_/C vssd1 vssd1 vccd1 vccd1 _12525_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_42_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12448_ hold137/A _12448_/B vssd1 vssd1 vccd1 vccd1 _12448_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09945__A1 _10245_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12379_ _09221_/Y _09562_/Y _09596_/B _12379_/B2 _12378_/X vssd1 vssd1 vccd1 vccd1
+ _12380_/B sky130_fd_sc_hd__a221o_1
XANTENNA__09945__B2 _10245_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06940_ instruction[28] _06944_/B vssd1 vssd1 vccd1 vccd1 _06940_/X sky130_fd_sc_hd__or2_1
XFILLER_0_66_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06871_ reg1_val[24] _06995_/A vssd1 vssd1 vccd1 vccd1 _06871_/X sky130_fd_sc_hd__and2_1
XANTENNA__10307__A2 _12144_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08610_ _08610_/A _08610_/B vssd1 vssd1 vccd1 vccd1 _08619_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08381__B1 _10476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13257__B2 _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09590_ hold235/A hold245/A vssd1 vssd1 vccd1 vccd1 _09590_/X sky130_fd_sc_hd__or2_1
XFILLER_0_89_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08541_ _08564_/A _08541_/B vssd1 vssd1 vccd1 vccd1 _08569_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08472_ _08515_/A2 _08649_/B1 _09472_/A _08540_/B vssd1 vssd1 vccd1 vccd1 _08473_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_58_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07423_ _09922_/A _07423_/B vssd1 vssd1 vccd1 vccd1 _07424_/B sky130_fd_sc_hd__xor2_1
XANTENNA_fanout147_A _09943_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08416__A _08664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07354_ _07655_/B _07354_/B vssd1 vssd1 vccd1 vccd1 _07356_/B sky130_fd_sc_hd__and2_1
XANTENNA__07239__A2 _08457_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07285_ _09836_/A _07285_/B vssd1 vssd1 vccd1 vccd1 _07287_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09024_ _09024_/A _09024_/B vssd1 vssd1 vccd1 vccd1 _09025_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_26_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold220 hold220/A vssd1 vssd1 vccd1 vccd1 hold220/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 hold231/A vssd1 vssd1 vccd1 vccd1 hold231/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 hold242/A vssd1 vssd1 vccd1 vccd1 hold242/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 hold253/A vssd1 vssd1 vccd1 vccd1 hold253/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 hold264/A vssd1 vssd1 vccd1 vccd1 hold264/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 hold275/A vssd1 vssd1 vccd1 vccd1 hold275/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 hold286/A vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09247__A _10297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold297 hold297/A vssd1 vssd1 vccd1 vccd1 hold297/X sky130_fd_sc_hd__dlygate4sd3_1
X_09926_ _09927_/B _09926_/B vssd1 vssd1 vccd1 vccd1 _09928_/A sky130_fd_sc_hd__and2b_1
XANTENNA__07990__A _08575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10849__A3 _10476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09857_ _09858_/B _09858_/A vssd1 vssd1 vccd1 vccd1 _09857_/Y sky130_fd_sc_hd__nand2b_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09788_ _09788_/A _09788_/B vssd1 vssd1 vccd1 vccd1 _09790_/B sky130_fd_sc_hd__xor2_2
X_08808_ _08807_/B _08807_/C _08920_/B vssd1 vssd1 vccd1 vccd1 _08809_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__11259__A0 _12420_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08739_ _08739_/A _08739_/B vssd1 vssd1 vccd1 vccd1 _08739_/Y sky130_fd_sc_hd__nand2_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ curr_PC[19] _11749_/C curr_PC[20] vssd1 vssd1 vccd1 vccd1 _11751_/B sky130_fd_sc_hd__a21oi_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ _10821_/A _10934_/C _10701_/C vssd1 vssd1 vccd1 vccd1 _10701_/X sky130_fd_sc_hd__or3_2
X_11681_ _11681_/A _11681_/B vssd1 vssd1 vccd1 vccd1 _11685_/B sky130_fd_sc_hd__xor2_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10856__A _11582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10632_ _10709_/B _10632_/B vssd1 vssd1 vccd1 vccd1 _10634_/C sky130_fd_sc_hd__or2_1
XFILLER_0_64_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07230__A _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10234__A1 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10234__B2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13351_ _13354_/CLK _13351_/D vssd1 vssd1 vccd1 vccd1 hold123/A sky130_fd_sc_hd__dfxtp_1
X_10563_ _10157_/X _10562_/X _11029_/S vssd1 vssd1 vccd1 vccd1 _10563_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08978__A2 _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12302_ _12302_/A _12302_/B vssd1 vssd1 vccd1 vccd1 _12302_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_63_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10785__A2 _11050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13282_ _13373_/CLK _13282_/D vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__dfxtp_1
X_10494_ _10495_/B _10494_/B vssd1 vssd1 vccd1 vccd1 _10634_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_32_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11734__A1 _11820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12233_ _12233_/A _12233_/B _12335_/B _12233_/D vssd1 vssd1 vccd1 vccd1 _12233_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_32_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12164_ _12164_/A _12164_/B _12164_/C vssd1 vssd1 vccd1 vccd1 _12165_/B sky130_fd_sc_hd__and3_1
XFILLER_0_31_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12095_ fanout41/X _08859_/Y _08974_/Y fanout43/X vssd1 vssd1 vccd1 vccd1 _12096_/B
+ sky130_fd_sc_hd__a22o_1
X_11115_ _11115_/A _11115_/B vssd1 vssd1 vccd1 vccd1 _11117_/C sky130_fd_sc_hd__xor2_1
X_11046_ _11017_/X _11018_/Y _11045_/X _11016_/Y vssd1 vssd1 vccd1 vccd1 _11046_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_127_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11498__B1 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07405__A _09779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08115__A0 _09341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12998__B1 _13257_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12997_ _13001_/A hold186/X vssd1 vssd1 vccd1 vccd1 hold187/A sky130_fd_sc_hd__and2_1
X_11948_ _12027_/A _11948_/B vssd1 vssd1 vccd1 vccd1 _11950_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10473__A1 _10240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11879_ _11962_/B _11879_/B vssd1 vssd1 vccd1 vccd1 _11881_/C sky130_fd_sc_hd__nand2_1
XANTENNA__11670__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10473__B2 _10473_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13142__A _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09615__B1 _07238_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09091__A1 _09298_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07070_ _07070_/A _07070_/B vssd1 vssd1 vccd1 vccd1 _07907_/C sky130_fd_sc_hd__nand2_4
XFILLER_0_70_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12981__A _13001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09091__B2 _09298_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09711_ _09711_/A _10004_/A _09711_/C _10137_/A vssd1 vssd1 vccd1 vccd1 _09711_/X
+ sky130_fd_sc_hd__or4_1
X_07972_ _07972_/A _07972_/B vssd1 vssd1 vccd1 vccd1 _07974_/B sky130_fd_sc_hd__or2_1
X_06923_ instruction[2] instruction[1] pred_val instruction[0] vssd1 vssd1 vccd1 vccd1
+ _06926_/B sky130_fd_sc_hd__and4b_4
XANTENNA__12150__A1 _09149_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06854_ _11541_/A _06852_/X _06853_/X vssd1 vssd1 vccd1 vccd1 _11632_/B sky130_fd_sc_hd__a21o_1
X_09642_ _09522_/A _09522_/B _09519_/A vssd1 vssd1 vccd1 vccd1 _09644_/B sky130_fd_sc_hd__a21o_1
X_06785_ reg2_val[5] _06783_/A _12444_/B vssd1 vssd1 vccd1 vccd1 _06972_/C sky130_fd_sc_hd__a21o_2
X_09573_ _09187_/X _09212_/X _09728_/S vssd1 vssd1 vccd1 vccd1 _09573_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout264_A _12796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ _08524_/A _08524_/B vssd1 vssd1 vccd1 vccd1 _08525_/B sky130_fd_sc_hd__and2_1
XANTENNA__08106__B1 _09940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12453__A2 _07147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08455_ _08657_/B _10221_/B2 _09770_/B2 _08649_/A2 vssd1 vssd1 vccd1 vccd1 _08456_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12205__A2 _12447_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07406_ _06993_/A fanout65/X fanout59/X _08613_/A vssd1 vssd1 vccd1 vccd1 _07407_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08386_ _08397_/B _08397_/A vssd1 vssd1 vccd1 vccd1 _08399_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__08409__B2 _08649_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08409__A1 _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07337_ fanout53/X _10245_/B2 _10245_/A1 fanout51/X vssd1 vssd1 vccd1 vccd1 _07338_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09082__A1 _08199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07985__A _08664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09082__B2 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07268_ _11081_/A _11080_/A vssd1 vssd1 vccd1 vccd1 _07268_/Y sky130_fd_sc_hd__nand2_4
X_07199_ _10813_/A _07199_/B vssd1 vssd1 vccd1 vccd1 _07199_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_60_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09007_ _09008_/A _09008_/B vssd1 vssd1 vccd1 vccd1 _09066_/C sky130_fd_sc_hd__and2_1
XANTENNA__11300__A _12096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07396__B2 _07221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07396__A1 _07217_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12141__A1 _12447_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09909_ _09909_/A _09909_/B vssd1 vssd1 vccd1 vccd1 _09910_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09705__A _09707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_9_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12920_ hold18/X hold248/X vssd1 vssd1 vccd1 vccd1 _13128_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07699__A2 _09298_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12851_ _11779_/A _12863_/A2 hold35/X _13210_/A vssd1 vssd1 vccd1 vccd1 _13286_/D
+ sky130_fd_sc_hd__o211a_1
X_11802_ _11802_/A _11802_/B vssd1 vssd1 vccd1 vccd1 _11802_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_68_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12782_ _12782_/A _12782_/B _12782_/C vssd1 vssd1 vccd1 vccd1 _12783_/B sky130_fd_sc_hd__and3_2
XANTENNA__10586__A _11398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11733_ _11820_/A _11733_/B vssd1 vssd1 vccd1 vccd1 _11733_/Y sky130_fd_sc_hd__nand2_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11652__A0 _09228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07320__A1 _09669_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11664_ _11929_/A _11664_/B vssd1 vssd1 vccd1 vccd1 _11668_/B sky130_fd_sc_hd__xnor2_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07320__B2 _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11404__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13403_ instruction[15] vssd1 vssd1 vccd1 vccd1 loadstore_dest[4] sky130_fd_sc_hd__buf_12
X_10615_ _10748_/A _07298_/B fanout8/A _10614_/Y vssd1 vssd1 vccd1 vccd1 _10707_/A
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_64_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11595_ _11595_/A _11595_/B vssd1 vssd1 vccd1 vccd1 _11610_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_24_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13334_ _13360_/CLK hold2/X vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10546_ _10280_/Y _10780_/A _10545_/Y vssd1 vssd1 vccd1 vccd1 _10546_/X sky130_fd_sc_hd__a21o_2
XFILLER_0_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10477_ _10478_/B _10478_/C _10207_/A vssd1 vssd1 vccd1 vccd1 _10479_/B sky130_fd_sc_hd__a21o_1
X_13265_ _13360_/CLK hold12/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12216_ curr_PC[25] curr_PC[26] _12216_/C vssd1 vssd1 vccd1 vccd1 _12220_/B sky130_fd_sc_hd__and3_1
X_13196_ hold262/X _13223_/A2 _13195_/X _13223_/B2 vssd1 vssd1 vccd1 vccd1 hold263/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11567__D _11567_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12147_ _12141_/Y _12142_/X _12146_/Y _12139_/X vssd1 vssd1 vccd1 vccd1 _12147_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10391__B1 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12078_ curr_PC[24] _12079_/B vssd1 vssd1 vccd1 vccd1 _12078_/X sky130_fd_sc_hd__or2_1
X_11029_ _09560_/Y _11028_/X _11029_/S vssd1 vssd1 vccd1 vccd1 _11030_/B sky130_fd_sc_hd__mux2_1
XANTENNA__13137__A _13147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08887__A1 _07959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08887__B2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11891__B1 _12049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12695__B _12696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10446__A1 _09242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09300__A2 _07608_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07311__A1 fanout68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08240_ _08314_/A _08314_/B vssd1 vssd1 vccd1 vccd1 _08315_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07311__B2 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_37 reg2_val[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_15 reg1_val[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_48 reg1_val[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 reg1_val[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08171_ _08172_/A _08172_/B vssd1 vssd1 vccd1 vccd1 _08171_/X sky130_fd_sc_hd__and2_1
X_07122_ reg1_val[20] _07107_/X _12740_/B reg1_val[21] _07585_/B1 vssd1 vssd1 vccd1
+ vccd1 _07129_/A sky130_fd_sc_hd__o311a_2
XFILLER_0_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_59 reg1_val[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07053_ _08502_/A _07053_/B vssd1 vssd1 vccd1 vccd1 _07057_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_112_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12371__A1 _12447_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07378__A1 _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07378__B2 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07955_ _07955_/A _07955_/B vssd1 vssd1 vccd1 vccd1 _08075_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_128_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06906_ _09239_/A vssd1 vssd1 vccd1 vccd1 _06906_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08878__A1 _07172_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09625_ _11406_/A fanout28/X fanout26/X _11309_/A vssd1 vssd1 vccd1 vccd1 _09626_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_37_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07886_ _07885_/A _07885_/B _07885_/C vssd1 vssd1 vccd1 vccd1 _07889_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__08878__B2 _09325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06837_ _07233_/A reg1_val[10] vssd1 vssd1 vccd1 vccd1 _06837_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_78_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06768_ reg1_val[8] _07215_/A vssd1 vssd1 vccd1 vccd1 _06768_/Y sky130_fd_sc_hd__nor2_1
X_09556_ _10049_/A _09556_/B vssd1 vssd1 vccd1 vccd1 _09557_/S sky130_fd_sc_hd__nand2_1
X_06699_ reg1_val[21] _06984_/B vssd1 vssd1 vccd1 vccd1 _11814_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09487_ _10479_/A _09487_/B vssd1 vssd1 vccd1 vccd1 _09488_/B sky130_fd_sc_hd__xnor2_1
X_08507_ _07030_/Y _12823_/A1 _07282_/Y _07038_/X vssd1 vssd1 vccd1 vccd1 _08508_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07302__A1 _10871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07302__B2 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08438_ _08438_/A _08438_/B vssd1 vssd1 vccd1 vccd1 _08465_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08369_ _08664_/A _08369_/B vssd1 vssd1 vccd1 vccd1 _08375_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_18_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11380_ _11381_/A _11381_/B vssd1 vssd1 vccd1 vccd1 _11479_/A sky130_fd_sc_hd__and2_1
XFILLER_0_104_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10400_ _10204_/A _10204_/B _10202_/X vssd1 vssd1 vccd1 vccd1 _10405_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_33_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10331_ _10331_/A _10542_/A _10661_/A _10661_/B vssd1 vssd1 vccd1 vccd1 _10331_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_104_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11030__A _12412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10262_ _10128_/A _10128_/B _10126_/X vssd1 vssd1 vccd1 vccd1 _10270_/A sky130_fd_sc_hd__a21oi_2
X_13050_ hold1/X _13094_/A2 _13101_/A2 hold156/X _13259_/A vssd1 vssd1 vccd1 vccd1
+ hold157/A sky130_fd_sc_hd__o221a_1
X_12001_ _11973_/Y _11974_/X _11977_/X _12000_/X vssd1 vssd1 vccd1 vccd1 _12001_/X
+ sky130_fd_sc_hd__o211a_1
X_10193_ _11393_/A _10193_/B vssd1 vssd1 vccd1 vccd1 _10197_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08030__A2 _08484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12903_ hold290/A hold54/X vssd1 vssd1 vccd1 vccd1 _12904_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__12796__A _12796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12834_ hold106/X _12862_/B vssd1 vssd1 vccd1 vccd1 hold107/A sky130_fd_sc_hd__or2_1
XFILLER_0_69_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12765_ reg1_val[25] _12790_/B vssd1 vssd1 vccd1 vccd1 _12770_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_29_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11716_ _11716_/A _11716_/B vssd1 vssd1 vccd1 vccd1 _11716_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12696_ reg1_val[11] _12696_/B vssd1 vssd1 vccd1 vccd1 _12697_/B sky130_fd_sc_hd__or2_1
XFILLER_0_25_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11647_ _11646_/B _11735_/B hold172/A vssd1 vssd1 vccd1 vccd1 _11648_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11578_ _11578_/A _11578_/B vssd1 vssd1 vccd1 vccd1 _11595_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08514__A _10243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13317_ _13373_/CLK hold174/X vssd1 vssd1 vccd1 vccd1 _13317_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06960__C _12438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10529_ _10405_/A _10405_/B _10403_/X vssd1 vssd1 vccd1 vccd1 _10530_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__06804__B1 _06803_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13248_ hold297/X _13248_/A2 _13247_/Y _13248_/B1 hold175/X vssd1 vssd1 vccd1 vccd1
+ hold176/A sky130_fd_sc_hd__a32o_1
XFILLER_0_58_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13179_ _13179_/A _13179_/B vssd1 vssd1 vccd1 vccd1 _13179_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__10364__B1 _07262_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06969__A _12438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06688__B _12665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07740_ _07557_/B _07557_/C _07557_/D _07558_/A vssd1 vssd1 vccd1 vccd1 _07741_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11864__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07671_ _07671_/A _07671_/B vssd1 vssd1 vccd1 vccd1 _07673_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_90_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06622_ reg1_val[29] _08973_/A vssd1 vssd1 vccd1 vccd1 _06622_/X sky130_fd_sc_hd__and2_1
X_09410_ _12644_/A curr_PC[1] vssd1 vssd1 vccd1 vccd1 _09412_/A sky130_fd_sc_hd__or2_1
XFILLER_0_90_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09341_ _09341_/A _09341_/B vssd1 vssd1 vccd1 vccd1 _09343_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12813__C1 _13147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07835__A2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09272_ _07417_/B _12823_/A1 _07282_/Y fanout42/X vssd1 vssd1 vccd1 vccd1 _09273_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11919__A1 _12446_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08223_ _08283_/A _08283_/B _08219_/X vssd1 vssd1 vccd1 vccd1 _08232_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_15_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout227_A _07117_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08154_ _08213_/A _08213_/B _08143_/X vssd1 vssd1 vccd1 vccd1 _08162_/B sky130_fd_sc_hd__a21o_1
X_07105_ reg1_val[8] reg1_val[9] reg1_val[10] _07105_/D vssd1 vssd1 vccd1 vccd1 _07248_/B
+ sky130_fd_sc_hd__or4_2
X_08085_ _08085_/A _08085_/B vssd1 vssd1 vccd1 vccd1 _08086_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07036_ _07036_/A _07036_/B vssd1 vssd1 vccd1 vccd1 _11946_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_3_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06879__A _12795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10370__A3 _10476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ _12404_/S _08985_/Y reg1_val[31] vssd1 vssd1 vccd1 vccd1 _12009_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__07771__B2 _06993_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07771__A1 _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10107__B1 _07274_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07938_ _07938_/A _07938_/B vssd1 vssd1 vccd1 vccd1 _08014_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07206__C _12359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07869_ _07869_/A _07869_/B vssd1 vssd1 vccd1 vccd1 _07951_/B sky130_fd_sc_hd__xnor2_1
X_10880_ _10742_/A _10742_/B _10759_/A vssd1 vssd1 vccd1 vccd1 _10890_/A sky130_fd_sc_hd__o21a_1
X_09608_ _09508_/A _09508_/B _09506_/Y vssd1 vssd1 vccd1 vccd1 _09623_/A sky130_fd_sc_hd__a21o_2
X_09539_ _09539_/A _09539_/B vssd1 vssd1 vccd1 vccd1 _09540_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_109_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09815__A3 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12550_ _12708_/B _12550_/B vssd1 vssd1 vccd1 vccd1 _12551_/B sky130_fd_sc_hd__or2_1
XFILLER_0_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11501_ _11500_/B _11501_/B vssd1 vssd1 vccd1 vccd1 _11502_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_108_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12481_ _12490_/A _12481_/B vssd1 vssd1 vccd1 vccd1 _12483_/C sky130_fd_sc_hd__nand2_1
XANTENNA__12555__S _12638_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11432_ _11430_/Y _11432_/B vssd1 vssd1 vccd1 vccd1 _11618_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07039__B1 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08334__A _08334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11363_ hold182/A _11363_/B vssd1 vssd1 vccd1 vccd1 _11461_/B sky130_fd_sc_hd__or2_1
X_13102_ hold16/X hold11/X fanout2/X vssd1 vssd1 vccd1 vccd1 hold303/A sky130_fd_sc_hd__nand3_1
XFILLER_0_34_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08251__A2 _08484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11294_ _12336_/A _11294_/B vssd1 vssd1 vccd1 vccd1 _11298_/A sky130_fd_sc_hd__xnor2_1
X_10314_ _12064_/S _12446_/C1 _10313_/Y _10308_/Y vssd1 vssd1 vccd1 vccd1 _10314_/X
+ sky130_fd_sc_hd__a31o_1
X_13033_ _13246_/A hold242/X vssd1 vssd1 vccd1 vccd1 _13326_/D sky130_fd_sc_hd__and2_1
XANTENNA__10803__S _11029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10245_ _10245_/A1 fanout13/X fanout8/X _10245_/B2 vssd1 vssd1 vccd1 vccd1 _10246_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10176_ reg1_val[6] curr_PC[6] vssd1 vssd1 vccd1 vccd1 _10176_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_100_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout190 _13248_/B1 vssd1 vssd1 vccd1 vccd1 _13223_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_88_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09503__A2 _12158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11310__A2 _12017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12817_ _07134_/Y _12805_/Y hold112/X _13147_/A vssd1 vssd1 vccd1 vccd1 _13269_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13063__A2 _12826_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09267__A1 _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09267__B2 _07554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12748_ _12760_/B _12748_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[21] sky130_fd_sc_hd__xor2_4
XFILLER_0_72_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12679_ reg1_val[8] _12680_/B vssd1 vssd1 vccd1 vccd1 _12679_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_114_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06971__B _07172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11377__A2 _11567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08244__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10585__B1 _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09890_ hold300/A _10049_/A _10166_/C _12205_/B1 vssd1 vssd1 vccd1 vccd1 _09890_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08910_ _08911_/B _08911_/A vssd1 vssd1 vccd1 vccd1 _08910_/Y sky130_fd_sc_hd__nand2b_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08841_ fanout63/X _10245_/B2 _10245_/A1 fanout61/X vssd1 vssd1 vccd1 vccd1 _08842_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ _08779_/B _08772_/B _08772_/C vssd1 vssd1 vccd1 vccd1 _08774_/A sky130_fd_sc_hd__nand3_1
XANTENNA__10949__A _11182_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07723_ _08561_/A2 _08112_/B fanout25/X _08561_/B1 vssd1 vssd1 vccd1 vccd1 _07724_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07654_ _07655_/A _07655_/B _07655_/C vssd1 vssd1 vccd1 vccd1 _08904_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06605_ _06949_/A _06605_/B vssd1 vssd1 vccd1 vccd1 is_store sky130_fd_sc_hd__nor2_8
XFILLER_0_125_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07585_ reg1_val[28] _08870_/C _12779_/B _07585_/B1 vssd1 vssd1 vccd1 vccd1 _07587_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09324_ _09324_/A _09324_/B vssd1 vssd1 vccd1 vccd1 _09335_/A sky130_fd_sc_hd__xnor2_2
X_09255_ _09233_/B instruction[5] _06889_/Y _06960_/D _09254_/X vssd1 vssd1 vccd1
+ vccd1 _09255_/X sky130_fd_sc_hd__a41o_1
XFILLER_0_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12014__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08206_ _08561_/B1 _08411_/B _10476_/A _08576_/A2 vssd1 vssd1 vccd1 vccd1 _08207_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_71_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09186_ reg1_val[6] reg1_val[25] _09211_/S vssd1 vssd1 vccd1 vccd1 _09186_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08137_ _09670_/A _08137_/B vssd1 vssd1 vccd1 vccd1 _08140_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10040__A2 _12446_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07993__A _09836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08068_ _08068_/A _08068_/B _08068_/C vssd1 vssd1 vccd1 vccd1 _08079_/A sky130_fd_sc_hd__or3_1
X_07019_ _07020_/A _07020_/B vssd1 vssd1 vccd1 vccd1 _07019_/X sky130_fd_sc_hd__and2_2
XFILLER_0_3_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11946__C _11946_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10030_ hold248/A _10031_/B vssd1 vssd1 vccd1 vccd1 _10030_/X sky130_fd_sc_hd__and2_1
XANTENNA__11828__B1 _11648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11981_ _06700_/A _11980_/X _09225_/Y vssd1 vssd1 vccd1 vccd1 _11981_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10932_ _09221_/Y _10914_/X _10920_/X _12446_/C1 _10931_/X vssd1 vssd1 vccd1 vccd1
+ _10933_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_98_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07233__A _07233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10863_ _10864_/A _10864_/B vssd1 vssd1 vccd1 vccd1 _10980_/C sky130_fd_sc_hd__or2_1
XANTENNA__13045__A2 _12820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12602_ reg1_val[21] curr_PC[21] _12631_/S vssd1 vssd1 vccd1 vccd1 _12603_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_94_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12253__B1 _12404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11056__A1 _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10794_ _06753_/Y _10792_/Y _10793_/Y vssd1 vssd1 vccd1 vccd1 _10818_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12533_ _12539_/B _12533_/B vssd1 vssd1 vccd1 vccd1 new_PC[10] sky130_fd_sc_hd__and2_4
XFILLER_0_81_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06791__B _06810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08472__A2 _08649_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12464_ _12644_/A curr_PC[1] _12471_/S vssd1 vssd1 vccd1 vccd1 _12466_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_34_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11415_ _11295_/Y _11298_/B _11303_/A vssd1 vssd1 vccd1 vccd1 _11415_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12395_ _12298_/A _12348_/A _12348_/B vssd1 vssd1 vccd1 vccd1 _12395_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__10567__B1 _12205_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11346_ _11239_/A _11237_/X _11259_/S vssd1 vssd1 vccd1 vccd1 _11346_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_61_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11277_ _11584_/A _11277_/B vssd1 vssd1 vccd1 vccd1 _11279_/B sky130_fd_sc_hd__xnor2_1
X_13016_ _13317_/Q _13171_/B2 _13209_/A2 hold188/X vssd1 vssd1 vccd1 vccd1 hold189/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10228_ _07232_/X _07596_/A _07596_/B _07360_/X _10725_/A vssd1 vssd1 vccd1 vccd1
+ _10229_/B sky130_fd_sc_hd__a32o_1
X_10159_ _10159_/A _10159_/B vssd1 vssd1 vccd1 vccd1 _10159_/Y sky130_fd_sc_hd__nor2_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07143__A _07143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08239__A _08334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07370_ _07370_/A _07370_/B vssd1 vssd1 vccd1 vccd1 _07571_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09040_ _09040_/A _09040_/B _09040_/C _09040_/D vssd1 vssd1 vccd1 vccd1 _10321_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_115_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09942_ _09942_/A _09942_/B vssd1 vssd1 vccd1 vccd1 _09963_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_40_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12224__A _12224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout294_A _12359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09873_ _10049_/A _08720_/A _08720_/B _10788_/A _09872_/Y vssd1 vssd1 vccd1 vccd1
+ _09873_/Y sky130_fd_sc_hd__a311oi_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _09922_/A _08824_/B vssd1 vssd1 vccd1 vccd1 _08825_/B sky130_fd_sc_hd__xor2_1
X_08755_ _08434_/A _08434_/B _08686_/B vssd1 vssd1 vccd1 vccd1 _08755_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09479__A1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09479__B2 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07706_ _07706_/A _07706_/B vssd1 vssd1 vccd1 vccd1 _07709_/B sky130_fd_sc_hd__xnor2_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ _08687_/B _08686_/B vssd1 vssd1 vccd1 vccd1 _08757_/B sky130_fd_sc_hd__or2_1
XANTENNA__08149__A _10207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07053__A _08502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07637_ _09922_/A _07637_/B vssd1 vssd1 vccd1 vccd1 _07639_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_36_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07568_ _07568_/A _07568_/B vssd1 vssd1 vccd1 vccd1 _07679_/B sky130_fd_sc_hd__xnor2_2
X_09307_ _09307_/A _09307_/B _09307_/C vssd1 vssd1 vccd1 vccd1 _09476_/B sky130_fd_sc_hd__and3_1
XFILLER_0_0_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11994__C1 _12376_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07499_ _07402_/A _07402_/B _07401_/A vssd1 vssd1 vccd1 vccd1 _07501_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_8_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09238_ _09239_/A _09239_/B vssd1 vssd1 vccd1 vccd1 _09238_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_51_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09169_ reg1_val[8] reg1_val[23] _09180_/S vssd1 vssd1 vccd1 vccd1 _09169_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08206__A2 _08411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11200_ _11201_/A _11201_/B vssd1 vssd1 vccd1 vccd1 _11202_/A sky130_fd_sc_hd__or2_1
X_12180_ _12041_/A _12110_/Y _12112_/B vssd1 vssd1 vccd1 vccd1 _12180_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09954__A2 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11131_ _11131_/A _11131_/B vssd1 vssd1 vccd1 vccd1 _11131_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_31_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11062_ _11393_/A _11062_/B vssd1 vssd1 vccd1 vccd1 _11066_/A sky130_fd_sc_hd__xnor2_1
X_10013_ _12438_/A _06826_/Y _10012_/Y vssd1 vssd1 vccd1 vccd1 _10014_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__10721__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11964_ _11964_/A _11964_/B vssd1 vssd1 vccd1 vccd1 _12113_/A sky130_fd_sc_hd__nand2_2
XANTENNA__13018__A2 _13171_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10915_ reg1_val[12] curr_PC[12] vssd1 vssd1 vccd1 vccd1 _10915_/Y sky130_fd_sc_hd__nand2_1
X_11895_ _08784_/B _11893_/X _11894_/Y vssd1 vssd1 vccd1 vccd1 _11895_/X sky130_fd_sc_hd__o21a_2
X_10846_ _11764_/A _07171_/A fanout38/X _11592_/A vssd1 vssd1 vccd1 vccd1 _10847_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12226__B1 fanout8/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08558__A_N _08564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10777_ _10777_/A _10777_/B _10777_/C vssd1 vssd1 vccd1 vccd1 _10778_/B sky130_fd_sc_hd__and3_1
XFILLER_0_82_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08445__A2 _08561_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12516_ _12525_/A _12516_/B vssd1 vssd1 vccd1 vccd1 _12518_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12447_ hold232/A _12417_/X _12447_/B1 vssd1 vssd1 vccd1 vccd1 _12448_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09945__A2 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12378_ _06622_/X _11995_/B _12377_/Y _06624_/B _12422_/A vssd1 vssd1 vccd1 vccd1
+ _12378_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_50_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11329_ _11329_/A _11329_/B vssd1 vssd1 vccd1 vccd1 _11331_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12979__A _13001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06870_ reg1_val[25] _06998_/A vssd1 vssd1 vccd1 vccd1 _06870_/X sky130_fd_sc_hd__and2_1
XANTENNA__06977__A _11038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08381__A1 _08649_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08381__B2 _09404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13257__A2 _13257_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08540_ _09404_/S _08540_/B vssd1 vssd1 vccd1 vccd1 _08541_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_82_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08471_ _08471_/A _08471_/B vssd1 vssd1 vccd1 vccd1 _08483_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_106_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07422_ _07554_/B _07173_/Y _07175_/A _07148_/Y vssd1 vssd1 vccd1 vccd1 _07423_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07353_ _07353_/A _07353_/B vssd1 vssd1 vccd1 vccd1 _07354_/B sky130_fd_sc_hd__or2_1
XFILLER_0_127_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07284_ _07959_/B _12823_/A1 _07282_/Y fanout29/X vssd1 vssd1 vccd1 vccd1 _07285_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11991__A2 _12447_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09023_ _09024_/A _09024_/B vssd1 vssd1 vccd1 vccd1 _09023_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_26_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold210 hold210/A vssd1 vssd1 vccd1 vccd1 hold210/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 hold232/A vssd1 vssd1 vccd1 vccd1 hold232/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11743__A2 _09422_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold243 hold301/A vssd1 vssd1 vccd1 vccd1 hold243/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 hold221/A vssd1 vssd1 vccd1 vccd1 hold221/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold287 hold287/A vssd1 vssd1 vccd1 vccd1 hold287/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 hold276/A vssd1 vssd1 vccd1 vccd1 hold276/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold254 hold254/A vssd1 vssd1 vccd1 vccd1 hold254/X sky130_fd_sc_hd__buf_1
Xhold265 hold265/A vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10951__B1 fanout8/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold298 hold298/A vssd1 vssd1 vccd1 vccd1 hold298/X sky130_fd_sc_hd__dlygate4sd3_1
X_09925_ _09925_/A _09925_/B vssd1 vssd1 vccd1 vccd1 _09927_/B sky130_fd_sc_hd__xnor2_1
X_09856_ _09856_/A _09856_/B vssd1 vssd1 vccd1 vccd1 _09858_/B sky130_fd_sc_hd__xnor2_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08807_ _08920_/B _08807_/B _08807_/C vssd1 vssd1 vccd1 vccd1 _08809_/A sky130_fd_sc_hd__and3_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ _09655_/B _09658_/B _09655_/A vssd1 vssd1 vccd1 vccd1 _09788_/B sky130_fd_sc_hd__o21ba_1
X_06999_ _06993_/A fanout68/X _06993_/Y fanout65/X vssd1 vssd1 vccd1 vccd1 _07000_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11259__A1 _09422_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08738_ _10668_/C _10668_/D _08737_/B _08737_/A _10668_/B vssd1 vssd1 vccd1 vccd1
+ _08744_/A sky130_fd_sc_hd__a221o_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08669_ _08714_/A _08717_/A _08668_/Y _08666_/B vssd1 vssd1 vccd1 vccd1 _08719_/B
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10700_ curr_PC[9] _10699_/C curr_PC[10] vssd1 vssd1 vccd1 vccd1 _10701_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__09872__A1 _10049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11680_ _11681_/A _11681_/B vssd1 vssd1 vccd1 vccd1 _11778_/A sky130_fd_sc_hd__and2b_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07511__A _08334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10631_ _10631_/A _10631_/B vssd1 vssd1 vccd1 vccd1 _10632_/B sky130_fd_sc_hd__and2_1
XFILLER_0_118_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10234__A2 _10234_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13350_ _13354_/CLK hold91/X vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__dfxtp_1
X_10562_ _09392_/X _09406_/X _11028_/S vssd1 vssd1 vccd1 vccd1 _10562_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_11_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13281_ _13373_/CLK _13281_/D vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__dfxtp_1
X_12301_ _12178_/A _12242_/Y _12244_/B vssd1 vssd1 vccd1 vccd1 _12301_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10493_ _12224_/A _10493_/B vssd1 vssd1 vccd1 vccd1 _10494_/B sky130_fd_sc_hd__xor2_1
X_12232_ _12233_/A _12233_/D _12233_/B vssd1 vssd1 vccd1 vccd1 _12234_/B sky130_fd_sc_hd__o21a_1
XANTENNA__08342__A _08342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12163_ _12164_/A _12164_/B _12164_/C vssd1 vssd1 vccd1 vccd1 _12239_/A sky130_fd_sc_hd__a21oi_1
X_12094_ _12164_/A _12094_/B vssd1 vssd1 vccd1 vccd1 _12098_/A sky130_fd_sc_hd__and2_1
X_11114_ _11115_/B _11115_/A vssd1 vssd1 vccd1 vccd1 _11224_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__11498__A1 _07032_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11045_ _09225_/Y _11021_/X _11022_/Y _11031_/X _11044_/Y vssd1 vssd1 vccd1 vccd1
+ _11045_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_127_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11498__B2 _11946_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12447__B1 _12447_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12996_ hold213/A _13000_/A2 _13257_/A2 hold185/X vssd1 vssd1 vccd1 vccd1 hold186/A
+ sky130_fd_sc_hd__a22o_1
X_11947_ fanout58/X _12009_/B _11945_/Y vssd1 vssd1 vccd1 vccd1 _11948_/B sky130_fd_sc_hd__o21a_1
XANTENNA__09312__B1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11670__B2 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11878_ _11878_/A _11878_/B _11878_/C vssd1 vssd1 vccd1 vccd1 _11879_/B sky130_fd_sc_hd__or3_1
XANTENNA__11670__A1 _11868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10473__A2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10829_ _11179_/A _10829_/B vssd1 vssd1 vccd1 vccd1 _10834_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_67_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09615__B2 _07417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09615__A1 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07140__B _12740_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09091__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11186__B1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08252__A _08454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07971_ _07927_/B _07971_/B vssd1 vssd1 vccd1 vccd1 _07972_/B sky130_fd_sc_hd__and2b_1
X_06922_ hold160/A _12803_/B vssd1 vssd1 vccd1 vccd1 busy sky130_fd_sc_hd__nor2_8
XANTENNA__10006__B _10006_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09710_ _09370_/X _09546_/X _09547_/X vssd1 vssd1 vccd1 vccd1 _09710_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09083__A _10092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06853_ reg1_val[18] _07087_/A vssd1 vssd1 vccd1 vccd1 _06853_/X sky130_fd_sc_hd__and2_1
X_09641_ _09485_/B _09488_/B _09485_/A vssd1 vssd1 vccd1 vccd1 _09644_/A sky130_fd_sc_hd__o21bai_2
X_06784_ reg2_val[5] _06783_/A _12444_/B vssd1 vssd1 vccd1 vccd1 _06827_/B sky130_fd_sc_hd__a21oi_2
X_09572_ _09205_/X _09209_/X _09727_/S vssd1 vssd1 vccd1 vccd1 _09572_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09303__B1 _09302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08523_ _08553_/A _08523_/B vssd1 vssd1 vccd1 vccd1 _08545_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08106__A1 _08561_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08106__B2 _08411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout257_A hold191/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12453__A3 _11995_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11661__A1 _11752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08454_ _08454_/A _08454_/B vssd1 vssd1 vccd1 vccd1 _08460_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07405_ _09779_/A _07411_/B vssd1 vssd1 vccd1 vccd1 _07428_/A sky130_fd_sc_hd__and2_1
X_08385_ _08383_/Y _08408_/B _08380_/X vssd1 vssd1 vccd1 vccd1 _08397_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__08409__A2 _08484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07336_ _07336_/A _07336_/B vssd1 vssd1 vccd1 vccd1 _07340_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_61_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09082__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07267_ _09794_/A _07267_/B vssd1 vssd1 vccd1 vccd1 _11080_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09006_ _09836_/A _09006_/B vssd1 vssd1 vccd1 vccd1 _09008_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13166__B2 _13171_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07198_ _10813_/A _07199_/B vssd1 vssd1 vccd1 vccd1 _07198_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__07396__A2 _08112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12412__A _12412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09908_ _11752_/S _09906_/Y _09907_/X _09905_/X vssd1 vssd1 vccd1 vccd1 dest_val[4]
+ sky130_fd_sc_hd__a31o_4
XANTENNA_fanout72_A _10974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09705__B _09707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09839_ _09960_/A _09841_/B vssd1 vssd1 vccd1 vccd1 _09842_/A sky130_fd_sc_hd__nand2_1
X_12850_ hold34/X _12862_/B vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__or2_1
XANTENNA__06845__A_N _07270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11801_ _11801_/A _11802_/B vssd1 vssd1 vccd1 vccd1 _11801_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_68_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _12782_/B _12782_/C _12782_/A vssd1 vssd1 vccd1 vccd1 _12787_/B sky130_fd_sc_hd__a21oi_2
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11732_ _11732_/A _11732_/B vssd1 vssd1 vccd1 vccd1 _11732_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_96_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11652__A1 _09422_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07320__A2 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07856__B1 _10476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11663_ fanout45/X fanout14/X fanout12/X fanout47/X vssd1 vssd1 vccd1 vccd1 _11664_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11404__A1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11404__B2 _11671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13402_ instruction[14] vssd1 vssd1 vccd1 vccd1 loadstore_dest[3] sky130_fd_sc_hd__buf_12
X_10614_ _10240_/A fanout7/X _10748_/A vssd1 vssd1 vccd1 vccd1 _10614_/Y sky130_fd_sc_hd__o21ai_1
X_11594_ _11594_/A _11594_/B vssd1 vssd1 vccd1 vccd1 _11595_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13333_ _13360_/CLK _13333_/D vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10545_ _10415_/A _10415_/B _10544_/X vssd1 vssd1 vccd1 vccd1 _10545_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13264_ _13296_/CLK _13264_/D vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfxtp_1
X_10476_ _10476_/A _10476_/B _10476_/C vssd1 vssd1 vccd1 vccd1 _10478_/C sky130_fd_sc_hd__or3_1
XFILLER_0_51_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13195_ hold264/A _13194_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13195_/X sky130_fd_sc_hd__mux2_1
X_12215_ _12215_/A _12215_/B _12215_/C _12214_/X vssd1 vssd1 vccd1 vccd1 _12215_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_32_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12146_ _12379_/B2 _10165_/X _12145_/X vssd1 vssd1 vccd1 vccd1 _12146_/Y sky130_fd_sc_hd__a21boi_1
XANTENNA__10391__B2 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10391__A1 _11868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12077_ _12051_/Y _12052_/X _12056_/X _12076_/X vssd1 vssd1 vccd1 vccd1 _12077_/X
+ sky130_fd_sc_hd__a211o_1
X_11028_ _10020_/B _10023_/Y _11028_/S vssd1 vssd1 vccd1 vccd1 _11028_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07416__A _09834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11891__A1 _11892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08887__A2 _07232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12979_ _13001_/A hold238/X vssd1 vssd1 vccd1 vccd1 _13299_/D sky130_fd_sc_hd__and2_1
XFILLER_0_87_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07311__A2 _08657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_38 reg2_val[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_27 reg2_val[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_16 reg1_val[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08170_ _08170_/A _08170_/B vssd1 vssd1 vccd1 vccd1 _08172_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_27_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_49 reg1_val[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07121_ _07121_/A _07121_/B vssd1 vssd1 vccd1 vccd1 _07121_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_15_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07052_ fanout68/X _08613_/A fanout56/X _06993_/A vssd1 vssd1 vccd1 vccd1 _07053_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09772__B1 _10725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07378__A2 _10473_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07954_ _07955_/A _07955_/B vssd1 vssd1 vccd1 vccd1 _07954_/Y sky130_fd_sc_hd__nand2_1
X_06905_ instruction[3] instruction[4] vssd1 vssd1 vccd1 vccd1 _09239_/A sky130_fd_sc_hd__nand2_4
X_07885_ _07885_/A _07885_/B _07885_/C vssd1 vssd1 vccd1 vccd1 _07889_/A sky130_fd_sc_hd__and3_1
X_06836_ _06896_/C _06834_/X _06835_/X vssd1 vssd1 vccd1 vccd1 _06836_/Y sky130_fd_sc_hd__a21oi_1
X_09624_ _09624_/A _09624_/B vssd1 vssd1 vccd1 vccd1 _09638_/A sky130_fd_sc_hd__or2_1
XANTENNA__08878__A2 _07362_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06767_ _06815_/A _06817_/B1 _12685_/B _06766_/X vssd1 vssd1 vccd1 vccd1 _07215_/A
+ sky130_fd_sc_hd__a31o_4
X_09555_ _09555_/A _10321_/C vssd1 vssd1 vccd1 vccd1 _09555_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06698_ reg1_val[21] _06698_/B vssd1 vssd1 vccd1 vccd1 _06698_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_78_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10437__A2 _11829_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09486_ fanout68/X _10245_/B2 _10245_/A1 fanout65/X vssd1 vssd1 vccd1 vccd1 _09487_/B
+ sky130_fd_sc_hd__o22a_1
X_08506_ _08506_/A _08506_/B vssd1 vssd1 vccd1 vccd1 _08527_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07302__A2 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08437_ _08437_/A _08437_/B vssd1 vssd1 vccd1 vccd1 _08465_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08368_ _06992_/A _10595_/A1 _10338_/B2 _08613_/A vssd1 vssd1 vccd1 vccd1 _08369_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08299_ _08575_/A _08299_/B vssd1 vssd1 vccd1 vccd1 _08349_/B sky130_fd_sc_hd__xnor2_4
X_07319_ _09672_/A _07319_/B vssd1 vssd1 vccd1 vccd1 _07323_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__10070__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10330_ _10143_/A _10329_/Y _10328_/Y vssd1 vssd1 vccd1 vccd1 _10330_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_104_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10261_ _10121_/A _10121_/B _10105_/A vssd1 vssd1 vccd1 vccd1 _10272_/A sky130_fd_sc_hd__a21bo_2
X_12000_ _09242_/B _11988_/X _11999_/X _11982_/X vssd1 vssd1 vccd1 vccd1 _12000_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11570__B1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10192_ _11406_/A fanout47/X fanout45/X _11309_/A vssd1 vssd1 vccd1 vccd1 _10193_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09515__B1 _10338_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12902_ hold54/X hold290/A vssd1 vssd1 vccd1 vccd1 _12902_/X sky130_fd_sc_hd__and2b_1
XANTENNA__09451__A _09922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07541__A2 _10337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12833_ _07195_/X _12863_/A2 hold95/X _13162_/A vssd1 vssd1 vccd1 vccd1 _13277_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06794__B _07117_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12764_ _12764_/A _12770_/A vssd1 vssd1 vccd1 vccd1 _12766_/A sky130_fd_sc_hd__nand2_2
X_11715_ _11529_/X _11885_/A _11714_/X vssd1 vssd1 vccd1 vccd1 _11715_/X sky130_fd_sc_hd__a21o_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ reg1_val[11] _12696_/B vssd1 vssd1 vccd1 vccd1 _12705_/A sky130_fd_sc_hd__nand2_1
X_11646_ hold172/A _11646_/B _11735_/B vssd1 vssd1 vccd1 vccd1 _11648_/B sky130_fd_sc_hd__and3_1
XFILLER_0_83_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11577_ _11578_/A _11578_/B vssd1 vssd1 vccd1 vccd1 _11689_/B sky130_fd_sc_hd__nand2b_1
X_13316_ _13316_/CLK _13316_/D vssd1 vssd1 vccd1 vccd1 hold172/A sky130_fd_sc_hd__dfxtp_1
X_10528_ _10528_/A _10528_/B vssd1 vssd1 vccd1 vccd1 _10530_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10061__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13247_ _12973_/A _13247_/B vssd1 vssd1 vccd1 vccd1 _13247_/Y sky130_fd_sc_hd__nand2b_1
X_10459_ _11284_/A _10459_/B vssd1 vssd1 vccd1 vccd1 _10461_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09754__B1 _12420_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13178_ _13178_/A _13178_/B vssd1 vssd1 vccd1 vccd1 _13179_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10364__B2 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10364__A1 _07171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09626__A _11582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06969__B _07147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12129_ _12364_/A _12129_/B _12129_/C vssd1 vssd1 vccd1 vccd1 _12129_/X sky130_fd_sc_hd__or3_1
XFILLER_0_74_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12987__A _13001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11864__B2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11864__A1 _12009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06985__A _07036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07670_ _07671_/B _07671_/A vssd1 vssd1 vccd1 vccd1 _07670_/Y sky130_fd_sc_hd__nand2b_1
X_06621_ _06619_/Y _06724_/B1 _06766_/B reg2_val[29] vssd1 vssd1 vccd1 vccd1 _08973_/A
+ sky130_fd_sc_hd__a2bb2o_2
X_09340_ _08112_/B _11198_/A _11093_/A fanout25/X vssd1 vssd1 vccd1 vccd1 _09341_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_75_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09271_ _09512_/A _09271_/B vssd1 vssd1 vccd1 vccd1 _09275_/B sky130_fd_sc_hd__or2_1
XFILLER_0_117_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08222_ _08222_/A _08222_/B vssd1 vssd1 vccd1 vccd1 _08283_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12227__A _12336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout122_A _08334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08153_ _08153_/A _08153_/B vssd1 vssd1 vccd1 vccd1 _08213_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07104_ _07104_/A _07104_/B vssd1 vssd1 vccd1 vccd1 _07244_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_16_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08084_ _08083_/A _08083_/B _08083_/C vssd1 vssd1 vccd1 vccd1 _08086_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07035_ _07036_/A _07036_/B vssd1 vssd1 vccd1 vccd1 _07035_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_43_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10970__A _12087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06690__A_N _07016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06879__B _07147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ _12404_/S _08985_/Y reg1_val[31] vssd1 vssd1 vccd1 vccd1 _12428_/B sky130_fd_sc_hd__o21a_4
XFILLER_0_11_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07771__A2 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07937_ _07937_/A _07937_/B vssd1 vssd1 vccd1 vccd1 _08014_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10107__A1 _07171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10107__B2 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11855__B2 _11929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07868_ _07868_/A _07868_/B vssd1 vssd1 vccd1 vccd1 _07951_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06819_ _12644_/A _09728_/S vssd1 vssd1 vccd1 vccd1 _06819_/X sky130_fd_sc_hd__and2_1
X_09607_ _09540_/A _09540_/B _09541_/Y vssd1 vssd1 vccd1 vccd1 _09704_/A sky130_fd_sc_hd__a21bo_2
X_07799_ _07823_/A _07823_/B vssd1 vssd1 vccd1 vccd1 _07869_/A sky130_fd_sc_hd__and2_1
XFILLER_0_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09538_ _09538_/A _09538_/B vssd1 vssd1 vccd1 vccd1 _09539_/B sky130_fd_sc_hd__xor2_2
XANTENNA_fanout35_A _07192_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11500_ _11501_/B _11500_/B vssd1 vssd1 vccd1 vccd1 _11502_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_109_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12280__A1 _12335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09469_ _09469_/A _09469_/B vssd1 vssd1 vccd1 vccd1 _09471_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout1_A fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12480_ _12655_/B _12480_/B vssd1 vssd1 vccd1 vccd1 _12481_/B sky130_fd_sc_hd__or2_1
XANTENNA__08615__A _09672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11431_ _11431_/A _11431_/B _11431_/C vssd1 vssd1 vccd1 vccd1 _11432_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_108_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08236__B1 _10476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07039__B2 _08649_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07039__A1 _08657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11362_ _06728_/B _11360_/Y _11361_/X _11359_/Y vssd1 vssd1 vccd1 vccd1 _11362_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11240__C1 _09225_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10313_ _10313_/A _10313_/B vssd1 vssd1 vccd1 vccd1 _10313_/Y sky130_fd_sc_hd__xnor2_1
X_13101_ hold16/X _13101_/A2 _11946_/C _13101_/B2 _13100_/Y vssd1 vssd1 vccd1 vccd1
+ hold17/A sky130_fd_sc_hd__o221a_1
XANTENNA__06798__B1 _06797_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11293_ _11671_/A fanout23/X fanout15/X fanout52/X vssd1 vssd1 vccd1 vccd1 _11294_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_104_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13032_ hold227/X _13248_/A2 _13248_/B1 hold241/X vssd1 vssd1 vccd1 vccd1 hold242/A
+ sky130_fd_sc_hd__a22o_1
X_10244_ _10243_/B _10243_/C _10243_/A vssd1 vssd1 vccd1 vccd1 _10247_/B sky130_fd_sc_hd__a21o_1
X_10175_ _10039_/A _10036_/Y _10038_/B vssd1 vssd1 vccd1 vccd1 _10179_/A sky130_fd_sc_hd__o21a_1
Xfanout191 _12803_/B vssd1 vssd1 vccd1 vccd1 _13248_/B1 sky130_fd_sc_hd__buf_4
XFILLER_0_89_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout180 _10246_/A vssd1 vssd1 vccd1 vccd1 _08564_/A sky130_fd_sc_hd__buf_12
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12816_ hold111/X _12816_/B vssd1 vssd1 vccd1 vccd1 hold112/A sky130_fd_sc_hd__or2_1
XFILLER_0_96_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09267__A2 _10337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12747_ reg1_val[20] _12755_/B _12743_/A vssd1 vssd1 vccd1 vccd1 _12748_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_29_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12678_ _12677_/A _12674_/Y _12676_/B vssd1 vssd1 vccd1 vccd1 _12682_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_127_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06971__C _07149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11629_ _11630_/A _11630_/B _11630_/C vssd1 vssd1 vccd1 vccd1 _11631_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_108_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10585__A1 _10944_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10585__B2 _07097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06699__B _06984_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11534__B1 _11567_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07202__A1 _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08840_ _08840_/A _08840_/B vssd1 vssd1 vccd1 vccd1 _08844_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_20_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _08765_/A _08765_/B _08769_/A _08766_/A vssd1 vssd1 vccd1 vccd1 _08772_/C
+ sky130_fd_sc_hd__a211o_1
X_07722_ _07728_/A _07728_/B vssd1 vssd1 vccd1 vccd1 _07722_/X sky130_fd_sc_hd__and2_1
XFILLER_0_95_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07653_ _08833_/A _07653_/B vssd1 vssd1 vccd1 vccd1 _07655_/C sky130_fd_sc_hd__or2_1
XANTENNA__07604__A _07604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06604_ instruction[3] _06605_/B vssd1 vssd1 vccd1 vccd1 is_load sky130_fd_sc_hd__nor2_8
XFILLER_0_88_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07584_ _07584_/A _07584_/B vssd1 vssd1 vccd1 vccd1 _07589_/B sky130_fd_sc_hd__xor2_1
X_09323_ _09323_/A vssd1 vssd1 vccd1 vccd1 _09463_/B sky130_fd_sc_hd__inv_2
XANTENNA__10965__A _11770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09254_ _09234_/B _06881_/X _06906_/Y _09220_/X _09253_/X vssd1 vssd1 vccd1 vccd1
+ _09254_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_35_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12014__A1 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12014__B2 _12233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09185_ reg1_val[7] reg1_val[24] _09211_/S vssd1 vssd1 vccd1 vccd1 _09185_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08205_ _08334_/A _08205_/B vssd1 vssd1 vccd1 vccd1 _08208_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08136_ _08627_/A2 _10595_/A1 fanout72/X _08641_/B vssd1 vssd1 vccd1 vccd1 _08137_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10576__B2 _12379_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10576__A1 _09221_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09430__A2 _08502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08067_ _08064_/A _08064_/C _08064_/B vssd1 vssd1 vccd1 vccd1 _08068_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07018_ _07215_/B _07070_/A _07070_/B _06984_/B vssd1 vssd1 vccd1 vccd1 _07020_/B
+ sky130_fd_sc_hd__a211o_2
XANTENNA__10328__A1 _10276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09266__A _09936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06952__B1 _06783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ _08969_/A _08969_/B vssd1 vssd1 vccd1 vccd1 _08970_/B sky130_fd_sc_hd__nand2_1
X_11980_ _11813_/S _11979_/X _11978_/X vssd1 vssd1 vccd1 vccd1 _11980_/X sky130_fd_sc_hd__a21o_1
X_10931_ _10922_/X _10923_/Y _11643_/B _12379_/B2 _10929_/X vssd1 vssd1 vccd1 vccd1
+ _10931_/X sky130_fd_sc_hd__a221o_1
XANTENNA__07514__A _10207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10862_ _12017_/A _10862_/B vssd1 vssd1 vccd1 vccd1 _10864_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _12611_/A _12601_/B vssd1 vssd1 vccd1 vccd1 new_PC[20] sky130_fd_sc_hd__xnor2_4
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10793_ _06753_/Y _10792_/Y _09225_/Y vssd1 vssd1 vccd1 vccd1 _10793_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__08457__B1 _08501_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12532_ _12532_/A _12532_/B _12532_/C vssd1 vssd1 vccd1 vccd1 _12533_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_93_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12005__A1 _12218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12463_ _12469_/A _12463_/B vssd1 vssd1 vccd1 vccd1 new_PC[0] sky130_fd_sc_hd__and2_4
X_11414_ _11308_/A _11308_/B _11311_/A vssd1 vssd1 vccd1 vccd1 _11419_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_81_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12394_ _12394_/A _12394_/B vssd1 vssd1 vccd1 vccd1 _12429_/B sky130_fd_sc_hd__or2_1
XFILLER_0_1_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11345_ _11809_/A _11345_/B _11345_/C _11345_/D vssd1 vssd1 vccd1 vccd1 _11345_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11276_ _07051_/X fanout30/X _07316_/Y fanout32/X vssd1 vssd1 vccd1 vccd1 _11277_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_120_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13015_ _13019_/A hold173/X vssd1 vssd1 vccd1 vccd1 hold174/A sky130_fd_sc_hd__and2_1
X_10227_ _10395_/B _10227_/B vssd1 vssd1 vccd1 vccd1 _10255_/A sky130_fd_sc_hd__or2_1
XANTENNA__10115__A _11393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
X_10158_ _11247_/A _10157_/X _09251_/A vssd1 vssd1 vccd1 vccd1 _10159_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10089_ _10089_/A _10089_/B vssd1 vssd1 vccd1 vccd1 _10104_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07143__B _07357_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10007__B1 _12356_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06777__A3 _12675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09941_ _11497_/A _09941_/B vssd1 vssd1 vccd1 vccd1 _09942_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09872_ _10049_/A _08720_/A _08720_/B vssd1 vssd1 vccd1 vccd1 _09872_/Y sky130_fd_sc_hd__a21oi_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _07121_/Y _07175_/A _07282_/Y _07554_/B vssd1 vssd1 vccd1 vccd1 _08824_/B
+ sky130_fd_sc_hd__a22o_1
X_08754_ _08753_/A _08753_/B _08751_/C _08751_/B _08751_/A vssd1 vssd1 vccd1 vccd1
+ _11345_/B sky130_fd_sc_hd__a2111o_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09479__A2 _10473_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07705_ _07705_/A _07705_/B vssd1 vssd1 vccd1 vccd1 _07709_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07334__A _09944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11286__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08685_ _08745_/A _08745_/B _08492_/X _08686_/B vssd1 vssd1 vccd1 vccd1 _08687_/C
+ sky130_fd_sc_hd__a211oi_1
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07636_ _07121_/Y _07554_/B _07175_/A _07134_/Y vssd1 vssd1 vccd1 vccd1 _07637_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07567_ _07748_/A _07748_/B _07564_/Y vssd1 vssd1 vccd1 vccd1 _07679_/A sky130_fd_sc_hd__o21ai_2
X_09306_ _09672_/A _09306_/B _09306_/C vssd1 vssd1 vccd1 vccd1 _09307_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09237_ _09239_/B _09237_/B vssd1 vssd1 vccd1 vccd1 _09237_/X sky130_fd_sc_hd__or2_1
XFILLER_0_63_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07498_ _07374_/A _07374_/B _07376_/B _07377_/B _07377_/A vssd1 vssd1 vccd1 vccd1
+ _07501_/A sky130_fd_sc_hd__o32a_2
XFILLER_0_29_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09168_ _09160_/X _09167_/X _10294_/S vssd1 vssd1 vccd1 vccd1 _09168_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09099_ _09099_/A _09099_/B vssd1 vssd1 vccd1 vccd1 _09100_/B sky130_fd_sc_hd__or2_1
X_08119_ _08119_/A _08119_/B vssd1 vssd1 vccd1 vccd1 _08120_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_102_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11130_ _06844_/Y _11129_/Y _11813_/S vssd1 vssd1 vccd1 vccd1 _11131_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07509__A _08454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11061_ _12009_/A fanout47/X fanout45/X fanout58/X vssd1 vssd1 vccd1 vccd1 _11062_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11973__B _12049_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10721__A1 _10974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10012_ _12438_/A _10012_/B vssd1 vssd1 vccd1 vccd1 _10012_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10721__B2 _10871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11963_ _11963_/A vssd1 vssd1 vccd1 vccd1 _11964_/B sky130_fd_sc_hd__inv_2
XFILLER_0_98_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10914_ _09740_/X _10913_/X _11029_/S vssd1 vssd1 vccd1 vccd1 _10914_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11894_ _08784_/B _11893_/X _10788_/A vssd1 vssd1 vccd1 vccd1 _11894_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07350__B1 _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10845_ _10845_/A _10845_/B vssd1 vssd1 vccd1 vccd1 _10848_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12226__B2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12226__A1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09890__A2 _10049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10776_ _10777_/A _10777_/B _10777_/C vssd1 vssd1 vccd1 vccd1 _10776_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_82_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12515_ _12680_/B _12515_/B vssd1 vssd1 vccd1 vccd1 _12516_/B sky130_fd_sc_hd__or2_1
XFILLER_0_81_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12446_ _12445_/A _12445_/B _12445_/Y _12446_/C1 vssd1 vssd1 vccd1 vccd1 _12446_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11737__B1 _11648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12377_ _06622_/X _12420_/A0 _12421_/A1 vssd1 vssd1 vccd1 vccd1 _12377_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__08602__B1 _08580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11328_ _11329_/A _11329_/B vssd1 vssd1 vccd1 vccd1 _11431_/B sky130_fd_sc_hd__or2_1
XFILLER_0_120_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11259_ _12420_/A0 _09422_/B _11259_/S vssd1 vssd1 vccd1 vccd1 _11259_/X sky130_fd_sc_hd__mux2_1
XANTENNA__06977__B _07195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08381__A2 _08411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12995__A _13001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06993__A _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08470_ _08470_/A _08470_/B vssd1 vssd1 vccd1 vccd1 _08496_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07421_ _07425_/A _07421_/B vssd1 vssd1 vccd1 vccd1 _07437_/B sky130_fd_sc_hd__or2_1
XFILLER_0_73_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07352_ _07353_/A _07353_/B vssd1 vssd1 vccd1 vccd1 _07655_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_128_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11976__B1 _10788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07283_ _07283_/A _07283_/B vssd1 vssd1 vccd1 vccd1 _07283_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_5_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08841__B1 _10245_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09809__A _11182_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09022_ _09022_/A _09022_/B vssd1 vssd1 vccd1 vccd1 _09024_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_31_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_3_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13309_/CLK sky130_fd_sc_hd__clkbuf_8
Xhold200 hold200/A vssd1 vssd1 vccd1 vccd1 hold200/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 hold211/A vssd1 vssd1 vccd1 vccd1 hold211/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold233 hold233/A vssd1 vssd1 vccd1 vccd1 hold233/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 hold222/A vssd1 vssd1 vccd1 vccd1 hold222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 hold244/A vssd1 vssd1 vccd1 vccd1 hold244/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout202_A _10243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07329__A _10479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold277 hold277/A vssd1 vssd1 vccd1 vccd1 hold277/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 hold266/A vssd1 vssd1 vccd1 vccd1 hold266/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 hold255/A vssd1 vssd1 vccd1 vccd1 hold255/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10951__A1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold288 hold288/A vssd1 vssd1 vccd1 vccd1 hold288/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10951__B2 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold299 hold67/A vssd1 vssd1 vccd1 vccd1 hold299/X sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ _09788_/A _09788_/B _09789_/X vssd1 vssd1 vccd1 vccd1 _09925_/B sky130_fd_sc_hd__o21bai_2
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12153__B1 _12631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09855_ _09697_/A _09697_/B _09695_/Y vssd1 vssd1 vccd1 vccd1 _09856_/B sky130_fd_sc_hd__a21boi_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08806_ _08799_/B _08799_/C _08805_/A _08805_/B vssd1 vssd1 vccd1 vccd1 _08807_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06998_ _06998_/A _06998_/B vssd1 vssd1 vccd1 vccd1 _06998_/X sky130_fd_sc_hd__xor2_4
X_09786_ _09633_/A _09633_/B _09629_/X vssd1 vssd1 vccd1 vccd1 _09788_/A sky130_fd_sc_hd__a21oi_2
X_08737_ _08737_/A _08737_/B vssd1 vssd1 vccd1 vccd1 _08737_/Y sky130_fd_sc_hd__nand2_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08668_ _08668_/A vssd1 vssd1 vccd1 vccd1 _08668_/Y sky130_fd_sc_hd__inv_2
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12208__A1 _12421_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07619_ _09944_/A _07619_/B vssd1 vssd1 vccd1 vccd1 _07620_/B sky130_fd_sc_hd__xnor2_2
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10630_ _10631_/A _10631_/B vssd1 vssd1 vccd1 vccd1 _10709_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_76_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08599_ _08627_/A2 _08649_/B1 _09472_/A _08641_/B vssd1 vssd1 vccd1 vccd1 _08600_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10561_ _10561_/A _10561_/B vssd1 vssd1 vccd1 vccd1 _10561_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_64_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13280_ _13373_/CLK _13280_/D vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__dfxtp_1
X_12300_ _12300_/A _12300_/B _12300_/C vssd1 vssd1 vccd1 vccd1 _12300_/X sky130_fd_sc_hd__or3_1
X_10492_ fanout43/X _07262_/X _07269_/Y fanout41/X vssd1 vssd1 vccd1 vccd1 _10493_/B
+ sky130_fd_sc_hd__a22o_1
X_12231_ _12284_/B _12236_/B vssd1 vssd1 vccd1 vccd1 _12237_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_121_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12162_ _12235_/A _12162_/B vssd1 vssd1 vccd1 vccd1 _12164_/C sky130_fd_sc_hd__nor2_1
X_11113_ _11113_/A _11113_/B vssd1 vssd1 vccd1 vccd1 _11115_/B sky130_fd_sc_hd__xnor2_1
X_12093_ _12093_/A _12093_/B vssd1 vssd1 vccd1 vccd1 _12094_/B sky130_fd_sc_hd__nand2_1
X_11044_ _09222_/Y _11030_/B _11043_/X vssd1 vssd1 vccd1 vccd1 _11044_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11498__A2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06797__B _06810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12995_ _13001_/A hold214/X vssd1 vssd1 vccd1 vccd1 _13307_/D sky130_fd_sc_hd__and2_1
X_11946_ _11945_/Y _11946_/B _11946_/C vssd1 vssd1 vccd1 vccd1 _12027_/A sky130_fd_sc_hd__and3b_1
XANTENNA__10458__B1 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12998__A2 _13000_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09312__B2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09312__A1 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11877_ _11878_/A _11878_/B _11878_/C vssd1 vssd1 vccd1 vccd1 _11962_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__11670__A2 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10828_ fanout75/X fanout14/X fanout12/X fanout78/X vssd1 vssd1 vccd1 vccd1 _10829_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09615__A2 _10337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09076__B1 _10245_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10759_ _10759_/A _10759_/B vssd1 vssd1 vccd1 vccd1 _10772_/A sky130_fd_sc_hd__and2_1
XFILLER_0_82_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08823__B1 _07282_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11186__A1 _07051_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11186__B2 _12169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12429_ _12429_/A _12429_/B vssd1 vssd1 vccd1 vccd1 _12430_/C sky130_fd_sc_hd__or2_1
XFILLER_0_112_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07149__A _07149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12135__A0 _10159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07970_ _07970_/A _07970_/B _07970_/C vssd1 vssd1 vccd1 vccd1 _07974_/A sky130_fd_sc_hd__and3_1
XFILLER_0_120_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06988__A _06998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06921_ _12805_/A _12804_/B vssd1 vssd1 vccd1 vccd1 _06921_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_93_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09551__A1 _09371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06852_ _11449_/A _06850_/Y _06851_/X vssd1 vssd1 vccd1 vccd1 _06852_/X sky130_fd_sc_hd__a21o_1
X_09640_ _09498_/A _09498_/B _09495_/A vssd1 vssd1 vccd1 vccd1 _09646_/A sky130_fd_sc_hd__o21a_1
X_06783_ _06783_/A _06783_/B _12670_/B vssd1 vssd1 vccd1 vccd1 _12412_/A sky130_fd_sc_hd__or3b_4
XFILLER_0_93_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09571_ _09434_/X _09570_/X _10297_/S vssd1 vssd1 vccd1 vccd1 _09571_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08522_ _08522_/A _08522_/B vssd1 vssd1 vccd1 vccd1 _08550_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08106__A2 _10476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08453_ _08649_/B1 _08484_/B _09479_/B1 _09404_/S vssd1 vssd1 vccd1 vccd1 _08454_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07612__A _09947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11134__A _11134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07404_ _07404_/A _07404_/B vssd1 vssd1 vccd1 vccd1 _07411_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_9_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08384_ _08384_/A _08384_/B vssd1 vssd1 vccd1 vccd1 _08408_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_45_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07335_ _07336_/A _07336_/B vssd1 vssd1 vccd1 vccd1 _07335_/Y sky130_fd_sc_hd__nor2_1
X_07266_ _10623_/A _07267_/B vssd1 vssd1 vccd1 vccd1 _11081_/A sky130_fd_sc_hd__or2_2
XFILLER_0_73_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13166__A2 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09005_ _10725_/A _07959_/B fanout29/X _07232_/X vssd1 vssd1 vccd1 vccd1 _09006_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08443__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07197_ _07233_/A _07133_/A _06974_/B _06978_/C _07215_/B vssd1 vssd1 vccd1 vccd1
+ _07199_/B sky130_fd_sc_hd__o41a_4
XFILLER_0_60_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12126__B1 _11637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09907_ curr_PC[4] _10045_/C vssd1 vssd1 vccd1 vccd1 _09907_/X sky130_fd_sc_hd__or2_1
XANTENNA__12412__B _12412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10688__A0 _09228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11309__A _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout65_A _06997_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06628__A2_N _06766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09838_ _09838_/A _09838_/B vssd1 vssd1 vccd1 vccd1 _09841_/B sky130_fd_sc_hd__or2_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09769_ _09676_/A _09676_/B _09674_/Y vssd1 vssd1 vccd1 vccd1 _09784_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_96_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11800_ _11800_/A _11966_/A vssd1 vssd1 vccd1 vccd1 _11802_/B sky130_fd_sc_hd__and2_1
XFILLER_0_95_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12780_ _12780_/A _12780_/B _12780_/C vssd1 vssd1 vccd1 vccd1 _12782_/C sky130_fd_sc_hd__or3_1
XANTENNA__07522__A _08564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11731_ _11642_/A _11642_/B _11640_/A vssd1 vssd1 vccd1 vccd1 _11732_/B sky130_fd_sc_hd__o21a_1
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07856__A1 _08501_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07856__B2 _10221_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _11567_/X _11626_/Y _11893_/A vssd1 vssd1 vccd1 vccd1 _11720_/A sky130_fd_sc_hd__a21o_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11404__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11593_ _11593_/A _11593_/B vssd1 vssd1 vccd1 vccd1 _11594_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_107_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10613_ _10514_/A _10514_/B _10511_/A vssd1 vssd1 vccd1 vccd1 _10616_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12574__S _12638_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13401_ instruction[13] vssd1 vssd1 vccd1 vccd1 loadstore_dest[2] sky130_fd_sc_hd__buf_12
X_10544_ _10276_/A _10276_/B _10415_/A _10415_/B vssd1 vssd1 vccd1 vccd1 _10544_/X
+ sky130_fd_sc_hd__o22a_1
X_13332_ _13360_/CLK hold41/X vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09449__A _09936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10475_ _07608_/A _07608_/B _08411_/B vssd1 vssd1 vccd1 vccd1 _10478_/B sky130_fd_sc_hd__a21o_1
X_13263_ _13396_/CLK hold69/X vssd1 vssd1 vccd1 vccd1 hold191/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13194_ _13194_/A _13194_/B vssd1 vssd1 vccd1 vccd1 _13194_/Y sky130_fd_sc_hd__xnor2_1
X_12214_ _08800_/Y _12212_/X _12213_/Y vssd1 vssd1 vccd1 vccd1 _12214_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_20_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12145_ _06998_/A _09257_/S _09222_/Y _10159_/B _12144_/X vssd1 vssd1 vccd1 vccd1
+ _12145_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_20_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10391__A2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12076_ _06946_/X _12064_/X _12075_/Y _12058_/Y vssd1 vssd1 vccd1 vccd1 _12076_/X
+ sky130_fd_sc_hd__a211o_1
X_11027_ _11027_/A _11027_/B vssd1 vssd1 vccd1 vccd1 _11027_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_99_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13093__A1 _12224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12978_ hold301/X _13000_/A2 _13257_/A2 hold237/X vssd1 vssd1 vccd1 vccd1 hold238/A
+ sky130_fd_sc_hd__a22o_1
X_11929_ _11929_/A _11929_/B vssd1 vssd1 vccd1 vccd1 _11933_/B sky130_fd_sc_hd__xor2_1
XANTENNA__10851__B1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_28 reg2_val[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_39 reg2_val[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_17 reg1_val[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10603__B1 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07120_ _07121_/A _07121_/B vssd1 vssd1 vccd1 vccd1 _07120_/X sky130_fd_sc_hd__and2_1
XFILLER_0_6_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07051_ _07215_/B _07045_/X _08973_/D _07049_/Y vssd1 vssd1 vccd1 vccd1 _07051_/X
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_42_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12356__B1 _12356_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09772__A1 _07554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09772__B2 _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09094__A _09302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07607__A _07608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07953_ _07953_/A _07953_/B vssd1 vssd1 vccd1 vccd1 _07955_/B sky130_fd_sc_hd__xnor2_4
X_06904_ instruction[6] _06902_/X _06903_/Y _06960_/D vssd1 vssd1 vccd1 vccd1 _06904_/X
+ sky130_fd_sc_hd__o211a_1
X_07884_ _07937_/A _07884_/B vssd1 vssd1 vccd1 vccd1 _07885_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_97_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06835_ reg1_val[9] _07238_/A vssd1 vssd1 vccd1 vccd1 _06835_/X sky130_fd_sc_hd__and2_1
XANTENNA__09822__A _09822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09623_ _09623_/A _09623_/B vssd1 vssd1 vccd1 vccd1 _09690_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_78_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06766_ reg2_val[8] _06766_/B vssd1 vssd1 vccd1 vccd1 _06766_/X sky130_fd_sc_hd__and2_1
X_09554_ _10137_/A _09554_/B vssd1 vssd1 vccd1 vccd1 _10321_/C sky130_fd_sc_hd__xor2_4
X_06697_ reg1_val[21] _06698_/B vssd1 vssd1 vccd1 vccd1 _11829_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09485_ _09485_/A _09485_/B vssd1 vssd1 vccd1 vccd1 _09488_/A sky130_fd_sc_hd__nor2_1
X_08505_ _08506_/A _08506_/B vssd1 vssd1 vccd1 vccd1 _08505_/X sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_4_13_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08436_ _08436_/A _08436_/B vssd1 vssd1 vccd1 vccd1 _08437_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_108_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08367_ _08367_/A _08367_/B vssd1 vssd1 vccd1 vccd1 _08397_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_116_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07318_ _06993_/Y fanout56/X fanout17/X _06993_/A vssd1 vssd1 vccd1 vccd1 _07319_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_116_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08298_ _08657_/B _10595_/A1 _10338_/B2 _08649_/A2 vssd1 vssd1 vccd1 vccd1 _08299_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_6_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10070__A1 _10245_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10070__B2 _10245_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07249_ reg1_val[11] _07249_/B vssd1 vssd1 vccd1 vccd1 _10060_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_33_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10260_ _10260_/A _10260_/B vssd1 vssd1 vccd1 vccd1 _10274_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__11570__B2 _12169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11570__A1 _07051_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ _10056_/A _10055_/B _10053_/X vssd1 vssd1 vccd1 vccd1 _10203_/A sky130_fd_sc_hd__a21o_2
XANTENNA__09515__A1 _07830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09515__B2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12901_ hold248/X hold18/X vssd1 vssd1 vccd1 vccd1 _13128_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__09732__A _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12569__S _12638_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ hold94/X _12862_/B vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__or2_1
XFILLER_0_69_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12763_ _12763_/A _12763_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[24] sky130_fd_sc_hd__xnor2_4
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _11523_/Y _11615_/Y _11617_/B vssd1 vssd1 vccd1 vccd1 _11714_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12694_ _12699_/B _12694_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[10] sky130_fd_sc_hd__and2_4
X_11645_ hold180/A _11645_/B vssd1 vssd1 vccd1 vccd1 _11735_/B sky130_fd_sc_hd__or2_1
XFILLER_0_37_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11576_ _12096_/A _11576_/B vssd1 vssd1 vccd1 vccd1 _11578_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_4_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13315_ _13316_/CLK _13315_/D vssd1 vssd1 vccd1 vccd1 hold180/A sky130_fd_sc_hd__dfxtp_1
X_10527_ _10527_/A _10527_/B vssd1 vssd1 vccd1 vccd1 _10528_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10061__A1 _12009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10061__B2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13246_ _13246_/A hold251/X vssd1 vssd1 vccd1 vccd1 _13391_/D sky130_fd_sc_hd__and2_1
X_10458_ fanout58/X fanout28/X fanout26/X _11868_/A vssd1 vssd1 vccd1 vccd1 _10459_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13177_ _13210_/A _13177_/B vssd1 vssd1 vccd1 vccd1 _13376_/D sky130_fd_sc_hd__and2_1
XANTENNA__10364__A2 _07256_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11561__A1 _09242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10389_ _10389_/A _10389_/B vssd1 vssd1 vccd1 vccd1 _10390_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_20_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12128_ _12364_/A _12129_/C _12129_/B vssd1 vssd1 vccd1 vccd1 _12128_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12059_ _11987_/A _11987_/B _11985_/A vssd1 vssd1 vccd1 vccd1 _12063_/A sky130_fd_sc_hd__o21a_1
XANTENNA__11864__A2 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06985__B _07014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06620_ reg2_val[29] _06766_/B _06724_/B1 _06619_/Y vssd1 vssd1 vccd1 vccd1 _06866_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10788__A _10788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06740__A1 _06927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12274__C1 _12631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12813__A1 _07173_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09270_ _09269_/B _09270_/B vssd1 vssd1 vccd1 vccd1 _09271_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_117_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08221_ _08221_/A _08221_/B vssd1 vssd1 vccd1 vccd1 _08283_/A sky130_fd_sc_hd__and2_1
XANTENNA__12508__A _12675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08152_ _08150_/A _08150_/B _08221_/A vssd1 vssd1 vccd1 vccd1 _08213_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_15_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10052__A1 _09302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07103_ _07443_/A _07375_/B vssd1 vssd1 vccd1 vccd1 _07104_/B sky130_fd_sc_hd__nand2_1
X_08083_ _08083_/A _08083_/B _08083_/C vssd1 vssd1 vccd1 vccd1 _08087_/A sky130_fd_sc_hd__and3_1
XFILLER_0_31_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07034_ _07014_/A _06987_/A _06986_/C _07094_/B vssd1 vssd1 vccd1 vccd1 _07036_/B
+ sky130_fd_sc_hd__a31oi_4
XANTENNA__12329__B1 _12319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout115_A _07217_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08985_ reg1_val[30] _08985_/B vssd1 vssd1 vccd1 vccd1 _08985_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07936_ _07936_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07938_/B sky130_fd_sc_hd__xor2_1
XANTENNA__10107__A2 _07269_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07508__B1 _09479_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11855__A2 _12158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07867_ _07867_/A _07867_/B vssd1 vssd1 vccd1 vccd1 _07868_/B sky130_fd_sc_hd__xor2_2
XANTENNA__13057__A1 _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06818_ _06992_/A _09419_/B vssd1 vssd1 vccd1 vccd1 _09418_/B sky130_fd_sc_hd__nand2_1
X_09606_ _09545_/A _09545_/B _09543_/X vssd1 vssd1 vccd1 vccd1 _09707_/A sky130_fd_sc_hd__a21oi_4
X_07798_ _09836_/A _07798_/B vssd1 vssd1 vccd1 vccd1 _07823_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11068__B1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12265__C1 _12446_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06749_ reg2_val[11] _06810_/B vssd1 vssd1 vccd1 vccd1 _06749_/X sky130_fd_sc_hd__and2_1
XANTENNA__07072__A _07907_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09537_ _09538_/A _09538_/B vssd1 vssd1 vccd1 vccd1 _09537_/X sky130_fd_sc_hd__and2_1
XFILLER_0_66_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout28_A _07231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09468_ _09467_/A _09467_/B _09469_/A vssd1 vssd1 vccd1 vccd1 _09621_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09399_ _09396_/X _09398_/X _10295_/S vssd1 vssd1 vccd1 vccd1 _09399_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08419_ _08452_/A _08452_/B vssd1 vssd1 vccd1 vccd1 _08423_/A sky130_fd_sc_hd__or2_2
X_11430_ _11431_/A _11431_/B _11431_/C vssd1 vssd1 vccd1 vccd1 _11430_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_80_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07039__A2 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08236__B2 _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08236__A1 _08576_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11361_ _06727_/B _12422_/A _11995_/B _06726_/X vssd1 vssd1 vccd1 vccd1 _11361_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10043__A1 _12365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10312_ _10310_/Y _10312_/B vssd1 vssd1 vccd1 vccd1 _10313_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13100_ _06571_/Y _06577_/A rst vssd1 vssd1 vccd1 vccd1 _13100_/Y sky130_fd_sc_hd__a21oi_1
X_11292_ _11417_/B _11292_/B vssd1 vssd1 vccd1 vccd1 _11304_/A sky130_fd_sc_hd__or2_1
X_13031_ _13162_/A hold228/X vssd1 vssd1 vccd1 vccd1 _13325_/D sky130_fd_sc_hd__and2_1
X_10243_ _10243_/A _10243_/B _10243_/C vssd1 vssd1 vccd1 vccd1 _10247_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_100_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10174_ _06781_/A _11554_/A _11829_/B _10155_/A _10173_/X vssd1 vssd1 vccd1 vccd1
+ _10174_/X sky130_fd_sc_hd__a221o_1
XANTENNA__07247__A _10207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout192 _12416_/C1 vssd1 vssd1 vccd1 vccd1 _12376_/C1 sky130_fd_sc_hd__buf_4
Xfanout170 _12871_/A2 vssd1 vssd1 vccd1 vccd1 _12863_/A2 sky130_fd_sc_hd__buf_4
Xfanout181 _10246_/A vssd1 vssd1 vccd1 vccd1 _10479_/A sky130_fd_sc_hd__buf_12
XFILLER_0_89_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12815_ _07166_/Y _13101_/B2 hold93/X _13147_/A vssd1 vssd1 vccd1 vccd1 _13268_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ _12744_/Y _12746_/B vssd1 vssd1 vccd1 vccd1 _12760_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12677_ _12677_/A _12677_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[7] sky130_fd_sc_hd__xor2_4
XANTENNA__06971__D _07959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11628_ _11893_/A _11567_/X _11626_/Y _12356_/B1 vssd1 vssd1 vccd1 vccd1 _11628_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_0_25_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10585__A2 _07171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11559_ hold180/A _11646_/B _11645_/B _11648_/A vssd1 vssd1 vccd1 vccd1 _11559_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_80_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07986__B1 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08541__A _08564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13229_ _13229_/A _13229_/B vssd1 vssd1 vccd1 vccd1 _13230_/B sky130_fd_sc_hd__nand2_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08770_ _08276_/Y _08326_/Y _08279_/Y vssd1 vssd1 vccd1 vccd1 _08772_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_79_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07721_ _07721_/A _07721_/B vssd1 vssd1 vccd1 vccd1 _07728_/B sky130_fd_sc_hd__xor2_1
X_07652_ _07652_/A _07652_/B vssd1 vssd1 vccd1 vccd1 _07653_/B sky130_fd_sc_hd__and2_1
XFILLER_0_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06603_ instruction[0] instruction[1] instruction[2] pred_val vssd1 vssd1 vccd1 vccd1
+ _06605_/B sky130_fd_sc_hd__or4bb_4
XFILLER_0_94_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07583_ _09341_/A _07583_/B vssd1 vssd1 vccd1 vccd1 _07584_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09322_ _09324_/A _09324_/B vssd1 vssd1 vccd1 vccd1 _09323_/A sky130_fd_sc_hd__and2_1
X_09253_ _09216_/X _09221_/Y _09252_/Y _12379_/B2 _09241_/X vssd1 vssd1 vccd1 vccd1
+ _09253_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12014__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09184_ _09168_/X _09183_/X _11246_/S vssd1 vssd1 vccd1 vccd1 _09184_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08204_ _09472_/A _08289_/B fanout75/X _08649_/B1 vssd1 vssd1 vccd1 vccd1 _08205_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08135_ _08564_/A _08135_/B vssd1 vssd1 vccd1 vccd1 _08140_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07977__B1 fanout72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09547__A _09548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08066_ _08066_/A _08066_/B vssd1 vssd1 vccd1 vccd1 _08068_/B sky130_fd_sc_hd__nand2_1
X_07017_ _07016_/A _06987_/A _06969_/Y _06698_/B vssd1 vssd1 vccd1 vccd1 _07020_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_12_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07067__A _09947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10328__A2 _10276_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08968_ _08969_/A _08969_/B vssd1 vssd1 vccd1 vccd1 _09064_/B sky130_fd_sc_hd__or2_1
XANTENNA__11828__A2 _11990_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07919_ _07915_/Y _07917_/X _07918_/A vssd1 vssd1 vccd1 vccd1 _07929_/B sky130_fd_sc_hd__a21oi_2
X_08899_ _08899_/A _08899_/B vssd1 vssd1 vccd1 vccd1 _08900_/B sky130_fd_sc_hd__nor2_2
X_10930_ _11247_/A _09730_/X _09251_/A vssd1 vssd1 vccd1 vccd1 _11643_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_98_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12600_ _12601_/B vssd1 vssd1 vccd1 vccd1 _12600_/Y sky130_fd_sc_hd__inv_2
X_10861_ _11093_/A fanout10/X fanout5/X _10974_/A vssd1 vssd1 vccd1 vccd1 _10862_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10792_ _12054_/S _06838_/Y _10791_/Y vssd1 vssd1 vccd1 vccd1 _10792_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__08457__A1 _06992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08457__B2 _08613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12531_ _12532_/A _12532_/B _12532_/C vssd1 vssd1 vccd1 vccd1 _12539_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12462_ _12642_/B _12462_/B vssd1 vssd1 vccd1 vccd1 _12463_/B sky130_fd_sc_hd__or2_1
XFILLER_0_54_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11413_ _11304_/A _11304_/B _11312_/X vssd1 vssd1 vccd1 vccd1 _11424_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__10016__A1 _11029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12393_ _12391_/A _12391_/B _12391_/C vssd1 vssd1 vccd1 vccd1 _12394_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__10567__A2 _11990_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11344_ _11809_/A _11345_/B _11345_/C _11345_/D vssd1 vssd1 vccd1 vccd1 _11344_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11275_ _11929_/A _11275_/B vssd1 vssd1 vccd1 vccd1 _11279_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13014_ hold172/X _13171_/B2 _13209_/A2 _13317_/Q vssd1 vssd1 vccd1 vccd1 hold173/A
+ sky130_fd_sc_hd__a22o_1
X_10226_ _10225_/A _11946_/C _10225_/C vssd1 vssd1 vccd1 vccd1 _10227_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
X_10157_ _11028_/S _09399_/X _11247_/C vssd1 vssd1 vccd1 vccd1 _10157_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10088_ _10088_/A _10088_/B vssd1 vssd1 vccd1 vccd1 _10089_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09893__B1 _12416_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12729_ _12729_/A _12739_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[17] sky130_fd_sc_hd__xnor2_4
XFILLER_0_29_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12492__S _12520_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09940_ _07221_/X _08877_/B fanout6/X _09940_/B2 vssd1 vssd1 vccd1 vccd1 _09941_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_111_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09871_ _09766_/X _09909_/B _09870_/Y vssd1 vssd1 vccd1 vccd1 _09871_/Y sky130_fd_sc_hd__a21oi_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12521__A _12685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ _08822_/A _08822_/B vssd1 vssd1 vccd1 vccd1 _08825_/A sky130_fd_sc_hd__nor2_1
X_08753_ _08753_/A _08753_/B vssd1 vssd1 vccd1 vccd1 _08753_/X sky130_fd_sc_hd__and2_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08136__B1 fanout72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07704_ _07804_/A _07804_/B _07693_/X vssd1 vssd1 vccd1 vccd1 _07731_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08684_ _08681_/A _08681_/B _08681_/C _08741_/B _08682_/Y vssd1 vssd1 vccd1 vccd1
+ _08745_/B sky130_fd_sc_hd__a41o_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07635_ _08893_/A _07635_/B vssd1 vssd1 vccd1 vccd1 _07639_/A sky130_fd_sc_hd__and2_1
X_07566_ _07566_/A _07566_/B vssd1 vssd1 vccd1 vccd1 _07748_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08446__A _08580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09305_ _09306_/B _09306_/C _09672_/A vssd1 vssd1 vccd1 vccd1 _09307_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09236_ _09239_/B _09237_/B vssd1 vssd1 vccd1 vccd1 _09236_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07497_ _07414_/A _07414_/B _07426_/B _07429_/A vssd1 vssd1 vccd1 vccd1 _07502_/A
+ sky130_fd_sc_hd__o31ai_4
XFILLER_0_8_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09167_ _09163_/X _09166_/X _09727_/S vssd1 vssd1 vccd1 vccd1 _09167_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_50_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09098_ _09099_/A _09099_/B vssd1 vssd1 vccd1 vccd1 _09330_/B sky130_fd_sc_hd__nand2_1
X_08118_ _08119_/B _08119_/A vssd1 vssd1 vccd1 vccd1 _08118_/X sky130_fd_sc_hd__and2b_1
X_08049_ _10092_/A _08049_/B vssd1 vssd1 vccd1 vccd1 _08051_/B sky130_fd_sc_hd__xnor2_1
X_11060_ _11060_/A _11060_/B vssd1 vssd1 vccd1 vccd1 _11100_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10011_ _06796_/A _09875_/B _06796_/B vssd1 vssd1 vccd1 vccd1 _10012_/B sky130_fd_sc_hd__a21boi_1
XANTENNA__10721__A2 _08877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07525__A _09944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11962_ _11962_/A _11962_/B _11962_/C vssd1 vssd1 vccd1 vccd1 _11963_/A sky130_fd_sc_hd__and3_1
XFILLER_0_86_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11682__B1 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10913_ _09882_/X _09884_/X _11246_/S vssd1 vssd1 vccd1 vccd1 _10913_/X sky130_fd_sc_hd__mux2_1
X_11893_ _11893_/A _11893_/B vssd1 vssd1 vccd1 vccd1 _11893_/X sky130_fd_sc_hd__or2_1
XANTENNA__07350__A1 _07134_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10844_ _10844_/A _10844_/B vssd1 vssd1 vccd1 vccd1 _10845_/B sky130_fd_sc_hd__nor2_1
XANTENNA__12226__A2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09627__B1 _10974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07350__B2 _07166_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12514_ _12680_/B _12515_/B vssd1 vssd1 vccd1 vccd1 _12525_/A sky130_fd_sc_hd__nand2_1
X_10775_ _10777_/A _10777_/B _10777_/C vssd1 vssd1 vccd1 vccd1 _10778_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12445_ _12445_/A _12445_/B vssd1 vssd1 vccd1 vccd1 _12445_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_34_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12376_ hold258/A _12449_/B1 _12414_/B _12375_/Y _12376_/C1 vssd1 vssd1 vccd1 vccd1
+ _12376_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_105_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08602__A1 _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11327_ _11215_/A _11215_/B _11216_/Y vssd1 vssd1 vccd1 vccd1 _11329_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_50_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11258_ _11258_/A _11258_/B vssd1 vssd1 vccd1 vccd1 _11258_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09915__A _12224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11189_ _11189_/A _11189_/B vssd1 vssd1 vccd1 vccd1 _11190_/B sky130_fd_sc_hd__nor2_1
X_10209_ _10209_/A _10209_/B vssd1 vssd1 vccd1 vccd1 _10211_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10173__B1 _11995_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09650__A _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06993__B _12644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07420_ _07420_/A _07420_/B vssd1 vssd1 vccd1 vccd1 _07421_/B sky130_fd_sc_hd__and2_1
XFILLER_0_119_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10228__B2 _10725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10228__A1 _07232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07351_ _09922_/A _07351_/B vssd1 vssd1 vccd1 vccd1 _07353_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_122_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07282_ _07283_/A _07283_/B vssd1 vssd1 vccd1 vccd1 _07282_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08841__A1 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08841__B2 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09021_ _08883_/A _08883_/B _08881_/X vssd1 vssd1 vccd1 vccd1 _09024_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_13_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold201 hold201/A vssd1 vssd1 vccd1 vccd1 hold201/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold234 hold234/A vssd1 vssd1 vccd1 vccd1 hold234/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 hold212/A vssd1 vssd1 vccd1 vccd1 hold212/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 hold223/A vssd1 vssd1 vccd1 vccd1 hold223/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold267 hold267/A vssd1 vssd1 vccd1 vccd1 hold267/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 hold278/A vssd1 vssd1 vccd1 vccd1 hold278/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10951__A2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold245 hold245/A vssd1 vssd1 vccd1 vccd1 hold245/X sky130_fd_sc_hd__buf_1
Xhold256 hold256/A vssd1 vssd1 vccd1 vccd1 hold256/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_111_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold289 hold289/A vssd1 vssd1 vccd1 vccd1 hold289/X sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ _09923_/A _09923_/B vssd1 vssd1 vccd1 vccd1 _09925_/A sky130_fd_sc_hd__xor2_1
XANTENNA__09825__A _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09854_ _09854_/A _09854_/B vssd1 vssd1 vccd1 vccd1 _09856_/A sky130_fd_sc_hd__xnor2_2
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10703__A2 _11050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08805_ _08805_/A _08805_/B vssd1 vssd1 vccd1 vccd1 _08805_/X sky130_fd_sc_hd__or2_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07345__A _09779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06997_ _06998_/A _06998_/B vssd1 vssd1 vccd1 vccd1 _06997_/Y sky130_fd_sc_hd__xnor2_2
X_09785_ _09668_/A _09668_/B _09665_/A vssd1 vssd1 vccd1 vccd1 _09790_/A sky130_fd_sc_hd__o21a_1
X_08736_ _08681_/B _08681_/C _08681_/A vssd1 vssd1 vccd1 vccd1 _08737_/B sky130_fd_sc_hd__a21o_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08667_ _08658_/A _08661_/A _08667_/S vssd1 vssd1 vccd1 vccd1 _08668_/A sky130_fd_sc_hd__mux2_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09609__B1 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07618_ fanout57/X _09943_/B2 _09650_/A fanout63/X vssd1 vssd1 vccd1 vccd1 _07619_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07080__A _07080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08598_ _09404_/S _08598_/B vssd1 vssd1 vccd1 vccd1 _08609_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_76_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07549_ _07708_/A _07708_/B vssd1 vssd1 vccd1 vccd1 _07556_/C sky130_fd_sc_hd__and2_1
XANTENNA_fanout10_A _08877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10560_ _10558_/Y _10560_/B vssd1 vssd1 vccd1 vccd1 _10561_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_36_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10491_ _12087_/B _10491_/B vssd1 vssd1 vccd1 vccd1 _10495_/B sky130_fd_sc_hd__xnor2_1
X_09219_ _09413_/A _09218_/X _11820_/A vssd1 vssd1 vccd1 vccd1 _09219_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_8_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12230_ _12230_/A _12230_/B vssd1 vssd1 vccd1 vccd1 _12236_/B sky130_fd_sc_hd__or2_1
XFILLER_0_17_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12161_ _12160_/B _12161_/B vssd1 vssd1 vccd1 vccd1 _12162_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_31_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11112_ _11113_/A _11113_/B vssd1 vssd1 vccd1 vccd1 _11224_/A sky130_fd_sc_hd__nand2_1
X_12092_ _12093_/A _12093_/B vssd1 vssd1 vccd1 vccd1 _12164_/A sky130_fd_sc_hd__or2_1
XANTENNA__12144__A1 _12144_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11043_ _11033_/Y _11034_/X _11042_/Y _10159_/A _11041_/X vssd1 vssd1 vccd1 vccd1
+ _11043_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12994_ hold208/X _13000_/A2 _13257_/A2 hold213/X vssd1 vssd1 vccd1 vccd1 hold214/A
+ sky130_fd_sc_hd__a22o_1
X_11945_ _12336_/A _11945_/B vssd1 vssd1 vccd1 vccd1 _11945_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__10458__B2 _11868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10458__A1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09312__A2 _08199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11876_ _11876_/A _11876_/B vssd1 vssd1 vccd1 vccd1 _11878_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10827_ _10715_/A _10715_/B _10720_/A vssd1 vssd1 vccd1 vccd1 _10836_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09076__B2 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09076__A1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10758_ _10758_/A _10758_/B vssd1 vssd1 vccd1 vccd1 _10759_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08823__A1 _07121_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08823__B2 _07554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12336__A _12336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12428_ fanout7/X _12428_/B vssd1 vssd1 vccd1 vccd1 _12433_/A sky130_fd_sc_hd__nand2_1
X_10689_ _12421_/A1 _10688_/X _06759_/A vssd1 vssd1 vccd1 vccd1 _10689_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11186__A2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12383__A1 _12336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12359_ _12359_/A _12359_/B vssd1 vssd1 vccd1 vccd1 _12359_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_23_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06920_ _12804_/A _12805_/B vssd1 vssd1 vccd1 vccd1 _12803_/B sky130_fd_sc_hd__nor2_4
XANTENNA__07165__A _07165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06851_ reg1_val[17] _07097_/A vssd1 vssd1 vccd1 vccd1 _06851_/X sky130_fd_sc_hd__and2_1
XANTENNA__09551__A2 _09371_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11894__B1 _10788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06782_ _06582_/Y _06610_/X _06613_/Y _12670_/B _06927_/A vssd1 vssd1 vccd1 vccd1
+ _06782_/X sky130_fd_sc_hd__o2111a_2
X_09570_ _09190_/X _09194_/X _09725_/S vssd1 vssd1 vccd1 vccd1 _09570_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_89_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08521_ _08521_/A _08521_/B _08521_/C vssd1 vssd1 vccd1 vccd1 _08683_/A sky130_fd_sc_hd__and3_1
XFILLER_0_77_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08452_ _08452_/A _08452_/B vssd1 vssd1 vccd1 vccd1 _08460_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07403_ _07430_/A _07430_/B vssd1 vssd1 vccd1 vccd1 _07403_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout145_A _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08383_ _08408_/A vssd1 vssd1 vccd1 vccd1 _08383_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12071__A0 _11995_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07334_ _09944_/A _07334_/B vssd1 vssd1 vccd1 vccd1 _07336_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_18_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07265_ reg1_val[14] _07265_/B vssd1 vssd1 vccd1 vccd1 _07267_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09004_ _09341_/A _09004_/B vssd1 vssd1 vccd1 vccd1 _09008_/A sky130_fd_sc_hd__xnor2_1
X_07196_ _07133_/A _06974_/B _06978_/C _07215_/B vssd1 vssd1 vccd1 vccd1 _07233_/B
+ sky130_fd_sc_hd__o31a_4
XFILLER_0_41_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09906_ curr_PC[4] _10045_/C vssd1 vssd1 vccd1 vccd1 _09906_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_6_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11309__B _12017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09837_ _09838_/A _09838_/B vssd1 vssd1 vccd1 vccd1 _09960_/A sky130_fd_sc_hd__nand2_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09768_ _09699_/A _09699_/B _09700_/Y vssd1 vssd1 vccd1 vccd1 _09861_/A sky130_fd_sc_hd__o21ai_4
XANTENNA_fanout58_A _07035_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08719_ _08719_/A _08719_/B vssd1 vssd1 vccd1 vccd1 _08720_/B sky130_fd_sc_hd__xor2_2
XANTENNA__09290__A _10749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11730_ _11730_/A _11730_/B vssd1 vssd1 vccd1 vccd1 _11732_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _09699_/A _09699_/B vssd1 vssd1 vccd1 vccd1 _09701_/B sky130_fd_sc_hd__xnor2_2
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07856__A2 _08411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11661_ _11752_/S _11658_/X _11660_/Y vssd1 vssd1 vccd1 vccd1 dest_val[19] sky130_fd_sc_hd__o21ai_4
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11592_ _11592_/A _12428_/B vssd1 vssd1 vccd1 vccd1 _11593_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_107_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10612_ _10612_/A _10612_/B vssd1 vssd1 vccd1 vccd1 _10620_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07069__B1 _07016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13400_ instruction[12] vssd1 vssd1 vccd1 vccd1 loadstore_dest[1] sky130_fd_sc_hd__buf_12
XFILLER_0_9_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13331_ _13360_/CLK _13331_/D vssd1 vssd1 vccd1 vccd1 hold165/A sky130_fd_sc_hd__dfxtp_1
X_10543_ _09375_/A _09375_/B _10542_/X vssd1 vssd1 vccd1 vccd1 _10543_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_9_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13262_ hold160/X _12803_/C _13142_/A vssd1 vssd1 vccd1 vccd1 hold161/A sky130_fd_sc_hd__o21a_1
X_10474_ _10748_/A _10474_/B vssd1 vssd1 vccd1 vccd1 _10482_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_122_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13193_ _13193_/A _13193_/B vssd1 vssd1 vccd1 vccd1 _13194_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09230__A1 _12144_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12213_ _08800_/Y _12212_/X _12365_/A vssd1 vssd1 vccd1 vccd1 _12213_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_102_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12144_ _12144_/A1 _12143_/X _06652_/B vssd1 vssd1 vccd1 vccd1 _12144_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_102_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06601__B _06944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12075_ _12066_/Y _12067_/X _12070_/X _12074_/Y vssd1 vssd1 vccd1 vccd1 _12075_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_47_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11026_ reg1_val[12] curr_PC[12] _10917_/X vssd1 vssd1 vccd1 vccd1 _11027_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09404__S _09404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11628__B1 _12356_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07713__A _10207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12825__C1 _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13093__A2 _13101_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12977_ _13001_/A hold244/X vssd1 vssd1 vccd1 vccd1 _13298_/D sky130_fd_sc_hd__and2_1
X_11928_ _11929_/A _11929_/B vssd1 vssd1 vccd1 vccd1 _12012_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10851__B2 _11946_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11859_ _11860_/A _11860_/B vssd1 vssd1 vccd1 vccd1 _11861_/A sky130_fd_sc_hd__or2_1
XANTENNA__10851__A1 _07032_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_29 reg2_val[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_18 reg1_val[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10603__B2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10603__A1 _12009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07050_ _07215_/B _07045_/X _08973_/D _07049_/Y vssd1 vssd1 vccd1 vccd1 _07050_/Y
+ sky130_fd_sc_hd__a31oi_2
XFILLER_0_12_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07480__B1 _09298_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09772__A2 _10234_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10906__A2 _11050_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07607__B _07608_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07952_ _07952_/A _07952_/B vssd1 vssd1 vccd1 vccd1 _07955_/A sky130_fd_sc_hd__nor2_2
X_06903_ instruction[6] _06963_/B vssd1 vssd1 vccd1 vccd1 _06903_/Y sky130_fd_sc_hd__nand2_1
X_07883_ _07883_/A _07883_/B vssd1 vssd1 vccd1 vccd1 _07884_/B sky130_fd_sc_hd__and2_1
X_06834_ _10423_/A _06832_/X _06833_/X vssd1 vssd1 vccd1 vccd1 _06834_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09822__B _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09622_ _09622_/A _09622_/B vssd1 vssd1 vccd1 vccd1 _09623_/B sky130_fd_sc_hd__nor2_2
X_09553_ _10138_/A _10138_/B _09551_/X _09552_/X vssd1 vssd1 vccd1 vccd1 _09554_/B
+ sky130_fd_sc_hd__o211a_4
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06765_ _06763_/Y _06765_/B vssd1 vssd1 vccd1 vccd1 _06896_/C sky130_fd_sc_hd__nand2b_1
X_08504_ _09670_/A _08504_/B vssd1 vssd1 vccd1 vccd1 _08506_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12831__A2 _12863_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06696_ _06694_/Y _06724_/B1 _06766_/B reg2_val[21] vssd1 vssd1 vccd1 vccd1 _06698_/B
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_77_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09484_ _09484_/A _09484_/B vssd1 vssd1 vccd1 vccd1 _09485_/B sky130_fd_sc_hd__and2_1
XFILLER_0_93_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08435_ _08435_/A _08435_/B vssd1 vssd1 vccd1 vccd1 _08467_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11799__B _11884_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08366_ _08400_/A _08400_/B vssd1 vssd1 vccd1 vccd1 _08403_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07317_ _10476_/B _10476_/C vssd1 vssd1 vccd1 vccd1 _12286_/A sky130_fd_sc_hd__or2_2
XFILLER_0_46_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08454__A _08454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08297_ _08297_/A _08297_/B vssd1 vssd1 vccd1 vccd1 _08349_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_6_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10070__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07248_ _07248_/A _07248_/B vssd1 vssd1 vccd1 vccd1 _07249_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_33_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07179_ _07162_/A _07162_/B _07372_/A vssd1 vssd1 vccd1 vccd1 _07242_/A sky130_fd_sc_hd__a21bo_2
X_10190_ _10077_/A _10077_/B _10068_/Y vssd1 vssd1 vccd1 vccd1 _10204_/A sky130_fd_sc_hd__a21bo_2
XANTENNA__07223__B1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11570__A2 _07171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08971__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09515__A2 _10595_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12900_ hold260/X hold46/X vssd1 vssd1 vccd1 vccd1 _13133_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__09732__B _09732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12831_ _07199_/X _12863_/A2 hold86/X _13246_/A vssd1 vssd1 vccd1 vccd1 _13276_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13075__A2 _12826_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12762_ _12763_/A _12763_/B vssd1 vssd1 vccd1 vccd1 _12770_/A sky130_fd_sc_hd__nand2b_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _11716_/B vssd1 vssd1 vccd1 vccd1 _11713_/Y sky130_fd_sc_hd__inv_2
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _12693_/A _12693_/B _12693_/C vssd1 vssd1 vccd1 vccd1 _12694_/B sky130_fd_sc_hd__nand3_1
X_11644_ _12064_/S _11642_/Y _11643_/Y _09242_/B vssd1 vssd1 vccd1 vccd1 _11657_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_84_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11575_ _06998_/X fanout43/X fanout41/X _07032_/Y vssd1 vssd1 vccd1 vccd1 _11576_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13314_ _13316_/CLK hold179/X vssd1 vssd1 vccd1 vccd1 hold177/A sky130_fd_sc_hd__dfxtp_1
X_10526_ _10525_/A _10525_/B _10527_/A vssd1 vssd1 vccd1 vccd1 _10526_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10061__A2 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06804__A3 _12655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13245_ hold250/X _13248_/B1 _13244_/X _13248_/A2 vssd1 vssd1 vccd1 vccd1 hold251/A
+ sky130_fd_sc_hd__a22o_1
X_10457_ _11179_/A _10457_/B vssd1 vssd1 vccd1 vccd1 _10461_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10306__A2_N _12422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09754__A2 _12144_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13176_ hold275/X _13223_/A2 _13175_/X _13223_/B2 vssd1 vssd1 vccd1 vccd1 _13177_/B
+ sky130_fd_sc_hd__a22o_1
X_10388_ _10389_/A _10389_/B vssd1 vssd1 vccd1 vccd1 _10390_/A sky130_fd_sc_hd__and2_1
XANTENNA__08962__B1 _11093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ _06672_/A _12125_/X _12126_/Y vssd1 vssd1 vccd1 vccd1 _12127_/X sky130_fd_sc_hd__o21a_1
X_12058_ _10049_/A _08795_/A _08795_/B _10788_/A _12057_/Y vssd1 vssd1 vccd1 vccd1
+ _12058_/Y sky130_fd_sc_hd__a311oi_4
X_11009_ _11009_/A _11229_/A vssd1 vssd1 vccd1 vccd1 _11009_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__06689__A2_N _06810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08539__A _08580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12274__B1 _09422_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12813__A2 _13101_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08220_ _08220_/A _08220_/B vssd1 vssd1 vccd1 vccd1 _08221_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08151_ _08220_/A _08220_/B vssd1 vssd1 vccd1 vccd1 _08221_/A sky130_fd_sc_hd__or2_1
XFILLER_0_15_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07102_ _07102_/A _07102_/B vssd1 vssd1 vccd1 vccd1 _07375_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08082_ _08082_/A _08082_/B vssd1 vssd1 vccd1 vccd1 _08083_/C sky130_fd_sc_hd__and2_1
XFILLER_0_31_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07033_ _06995_/A _06994_/X _06995_/Y _06987_/Y vssd1 vssd1 vccd1 vccd1 _07033_/X
+ sky130_fd_sc_hd__a22o_2
XANTENNA__12329__B2 _09221_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12329__A1 _12379_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout108_A _07283_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07220__A3 _07117_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08984_ _08984_/A _08984_/B vssd1 vssd1 vccd1 vccd1 _09000_/A sky130_fd_sc_hd__xnor2_2
X_07935_ _07935_/A _07935_/B vssd1 vssd1 vccd1 vccd1 _07938_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07508__A1 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07508__B2 fanout72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10512__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09605_ _09765_/A _09765_/B _10321_/C _10049_/A vssd1 vssd1 vccd1 vccd1 _09715_/A
+ sky130_fd_sc_hd__o31ai_1
XFILLER_0_3_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07866_ _07866_/A _07866_/B vssd1 vssd1 vccd1 vccd1 _07868_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06817_ reg2_val[0] _06766_/B _06817_/B1 _06815_/X vssd1 vssd1 vccd1 vccd1 _06817_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13057__A2 _12826_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07797_ _07173_/Y _07959_/B fanout29/X _07148_/Y vssd1 vssd1 vccd1 vccd1 _07798_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11068__A1 _12169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11068__B2 _06998_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06748_ _10927_/S _06748_/B vssd1 vssd1 vccd1 vccd1 _06897_/D sky130_fd_sc_hd__or2_2
XANTENNA__07072__B _07907_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09536_ _09351_/A _09351_/B _09349_/Y vssd1 vssd1 vccd1 vccd1 _09538_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_109_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09467_ _09467_/A _09467_/B vssd1 vssd1 vccd1 vccd1 _09469_/B sky130_fd_sc_hd__nor2_1
X_06679_ reg1_val[23] _07036_/A vssd1 vssd1 vccd1 vccd1 _06680_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_19_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08418_ _08575_/A _08418_/B vssd1 vssd1 vccd1 vccd1 _08452_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09398_ _09244_/X _09397_/X _09728_/S vssd1 vssd1 vccd1 vccd1 _09398_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08236__A2 _08411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08349_ _08349_/A _08349_/B vssd1 vssd1 vccd1 vccd1 _08351_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_19_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11360_ _06726_/X _12420_/A0 _12421_/A1 vssd1 vssd1 vccd1 vccd1 _11360_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07444__B1 _10240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10311_ reg1_val[7] curr_PC[7] vssd1 vssd1 vccd1 vccd1 _10312_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07995__A1 _09836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11291_ _11291_/A _11291_/B vssd1 vssd1 vccd1 vccd1 _11292_/B sky130_fd_sc_hd__and2_1
X_13030_ hold224/X _13248_/A2 _13248_/B1 hold227/X vssd1 vssd1 vccd1 vccd1 hold228/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10242_ _10749_/A _10242_/B _10242_/C vssd1 vssd1 vccd1 vccd1 _10243_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_100_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10173_ _07283_/A _12422_/A _11995_/B _06779_/X _10172_/Y vssd1 vssd1 vccd1 vccd1
+ _10173_/X sky130_fd_sc_hd__a221o_1
XANTENNA__09743__A _12438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout171 _12805_/Y vssd1 vssd1 vccd1 vccd1 _12871_/A2 sky130_fd_sc_hd__buf_2
Xfanout182 _07086_/Y vssd1 vssd1 vccd1 vccd1 _10246_/A sky130_fd_sc_hd__buf_8
Xfanout160 _06963_/Y vssd1 vssd1 vccd1 vccd1 _11892_/A sky130_fd_sc_hd__buf_4
XFILLER_0_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout193 _09239_/X vssd1 vssd1 vccd1 vccd1 _12416_/C1 sky130_fd_sc_hd__buf_4
XFILLER_0_88_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13048__A2 _06577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12814_ hold92/X _12820_/B vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__or2_1
XFILLER_0_96_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10806__A1 _11990_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12745_ reg1_val[21] _12755_/B vssd1 vssd1 vccd1 vccd1 _12746_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13204__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12676_ _12674_/Y _12676_/B vssd1 vssd1 vccd1 vccd1 _12677_/B sky130_fd_sc_hd__nand2b_2
XANTENNA__07683__B1 _09479_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11627_ _11893_/A _11567_/X _11626_/Y vssd1 vssd1 vccd1 vccd1 _11627_/X sky130_fd_sc_hd__o21a_1
X_11558_ _11646_/B _11645_/B hold180/A vssd1 vssd1 vccd1 vccd1 _11558_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11231__A1 _10283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10034__A2 _12420_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10509_ _10510_/A _10510_/B vssd1 vssd1 vccd1 vccd1 _10511_/A sky130_fd_sc_hd__and2_1
XFILLER_0_80_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07986__A1 _08641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07986__B2 _08627_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11489_ _11929_/A _11489_/B vssd1 vssd1 vccd1 vccd1 _11490_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10563__S _11029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13228_ _13249_/A _13228_/B vssd1 vssd1 vccd1 vccd1 _13387_/D sky130_fd_sc_hd__and2_1
XFILLER_0_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13159_ _13159_/A _13159_/B vssd1 vssd1 vccd1 vccd1 _13159_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08935__B1 _07282_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07720_ _07755_/A _07755_/B _07716_/X vssd1 vssd1 vccd1 vccd1 _07728_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07173__A _10297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07651_ _07652_/A _07652_/B vssd1 vssd1 vccd1 vccd1 _08833_/A sky130_fd_sc_hd__nor2_1
X_06602_ instruction[15] _06590_/X _06601_/X _06675_/B vssd1 vssd1 vccd1 vccd1 reg1_idx[4]
+ sky130_fd_sc_hd__o211a_4
X_07582_ _07198_/Y _08112_/B _10599_/A fanout25/X vssd1 vssd1 vccd1 vccd1 _07583_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09321_ _09321_/A _09321_/B vssd1 vssd1 vccd1 vccd1 _09324_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_48_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09252_ _12445_/A vssd1 vssd1 vccd1 vccd1 _09252_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11470__A1 _10788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09183_ _09175_/X _09182_/X _10295_/S vssd1 vssd1 vccd1 vccd1 _09183_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09415__A1 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08203_ _08454_/A _08203_/B vssd1 vssd1 vccd1 vccd1 _08208_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08134_ _08515_/A2 _10221_/B2 _08501_/B1 _08540_/B vssd1 vssd1 vccd1 vccd1 _08135_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07977__A1 _08538_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07977__B2 _08598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09179__A0 _11134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09547__B _09548_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08065_ _08065_/A _08065_/B _08065_/C vssd1 vssd1 vccd1 vccd1 _08066_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_31_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07016_ _07016_/A _07094_/B vssd1 vssd1 vccd1 vccd1 _07070_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_3_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06952__A2 _09242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12701__B _12702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08967_ _09667_/A _08967_/B vssd1 vssd1 vccd1 vccd1 _08969_/B sky130_fd_sc_hd__xnor2_1
X_07918_ _07918_/A _07918_/B _07915_/Y vssd1 vssd1 vccd1 vccd1 _07970_/A sky130_fd_sc_hd__or3b_1
X_08898_ _08898_/A _08898_/B vssd1 vssd1 vccd1 vccd1 _08899_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_98_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07849_ _08580_/A _07849_/B vssd1 vssd1 vccd1 vccd1 _07850_/B sky130_fd_sc_hd__xnor2_1
X_10860_ _12157_/A _10860_/B vssd1 vssd1 vccd1 vccd1 _10864_/A sky130_fd_sc_hd__xnor2_1
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09519_ _09519_/A _09519_/B vssd1 vssd1 vccd1 vccd1 _09522_/A sky130_fd_sc_hd__nor2_1
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10791_ _11813_/S _10791_/B vssd1 vssd1 vccd1 vccd1 _10791_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_39_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08457__A2 _08457_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _12539_/A _12530_/B vssd1 vssd1 vccd1 vccd1 _12532_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_93_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12461_ _12642_/B _12462_/B vssd1 vssd1 vccd1 vccd1 _12469_/A sky130_fd_sc_hd__nand2_1
X_11412_ _11412_/A _11412_/B vssd1 vssd1 vccd1 vccd1 _11426_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_34_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12392_ _12394_/A vssd1 vssd1 vccd1 vccd1 _12392_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_62_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11343_ _11272_/X _11567_/B _11342_/Y vssd1 vssd1 vccd1 vccd1 _11343_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11274_ _12233_/A fanout47/X fanout45/X _12087_/A vssd1 vssd1 vccd1 vccd1 _11275_/B
+ sky130_fd_sc_hd__o22a_1
X_13013_ _13210_/A hold181/X vssd1 vssd1 vccd1 vccd1 _13316_/D sky130_fd_sc_hd__and2_1
X_10225_ _10225_/A _11946_/C _10225_/C vssd1 vssd1 vccd1 vccd1 _10395_/B sky130_fd_sc_hd__and3_1
X_10156_ _10155_/A _10155_/B _09225_/Y vssd1 vssd1 vccd1 vccd1 _10156_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_89_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10087_ _10088_/A _10088_/B vssd1 vssd1 vccd1 vccd1 _10087_/Y sky130_fd_sc_hd__nand2_1
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08817__A _09834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10989_ _10836_/A _10836_/B _10837_/Y vssd1 vssd1 vccd1 vccd1 _10995_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12728_ reg1_val[17] _12755_/B vssd1 vssd1 vccd1 vccd1 _12739_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12659_ reg1_val[4] _12660_/B vssd1 vssd1 vccd1 vccd1 _12659_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_127_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09648__A _10748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07408__B1 _08649_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12401__B1 _09149_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap102 _07983_/B vssd1 vssd1 vccd1 vccd1 _10944_/B2 sky130_fd_sc_hd__buf_4
Xmax_cap113 _10225_/A vssd1 vssd1 vccd1 vccd1 _12823_/A1 sky130_fd_sc_hd__buf_4
XFILLER_0_52_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09870_ _09766_/X _09909_/B _12356_/B1 vssd1 vssd1 vccd1 vccd1 _09870_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08821_ _08821_/A _08821_/B vssd1 vssd1 vccd1 vccd1 _08822_/B sky130_fd_sc_hd__nor2_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08752_ _08687_/B _08687_/C _08757_/A vssd1 vssd1 vccd1 vccd1 _08753_/B sky130_fd_sc_hd__o21ai_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08136__A1 _08627_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08683_ _08683_/A _08683_/B vssd1 vssd1 vccd1 vccd1 _08741_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08136__B2 _08641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07703_ _07703_/A _07703_/B vssd1 vssd1 vccd1 vccd1 _07804_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout175_A _12816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07634_ _07634_/A _07634_/B vssd1 vssd1 vccd1 vccd1 _07635_/B sky130_fd_sc_hd__or2_1
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07565_ _07565_/A _07565_/B vssd1 vssd1 vccd1 vccd1 _07748_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_118_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09304_ _09306_/B _09306_/C _09672_/A vssd1 vssd1 vccd1 vccd1 _09476_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__07647__B1 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07496_ _07561_/A _07561_/B _07467_/X vssd1 vssd1 vccd1 vccd1 _07503_/A sky130_fd_sc_hd__a21o_1
X_09235_ _12365_/A _11995_/B _08663_/A vssd1 vssd1 vccd1 vccd1 _09235_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_8_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13196__B2 _13223_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09166_ _09164_/X _09165_/X _09383_/S vssd1 vssd1 vccd1 vccd1 _09166_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_114_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09097_ _09097_/A _09097_/B vssd1 vssd1 vccd1 vccd1 _09099_/B sky130_fd_sc_hd__xor2_1
X_08117_ _08121_/A _08121_/B _08111_/X vssd1 vssd1 vccd1 vccd1 _08119_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_16_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07078__A _07078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08048_ _08576_/A2 _08199_/B fanout33/X _09472_/A vssd1 vssd1 vccd1 vccd1 _08049_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10010_ _11630_/A _10010_/B _10010_/C vssd1 vssd1 vccd1 vccd1 _10010_/X sky130_fd_sc_hd__or3_1
XANTENNA_fanout88_A _11284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06710__A _06723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09999_ _09999_/A _09999_/B vssd1 vssd1 vccd1 vccd1 _10542_/A sky130_fd_sc_hd__xnor2_4
X_11961_ _11962_/A _11962_/B _11962_/C vssd1 vssd1 vccd1 vccd1 _11964_/A sky130_fd_sc_hd__a21o_1
X_10912_ _06897_/D _10910_/X _10911_/Y vssd1 vssd1 vccd1 vccd1 _10933_/C sky130_fd_sc_hd__o21a_1
XANTENNA__11682__A1 _12169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11682__B2 _06998_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11892_ _11892_/A _11892_/B _12049_/A vssd1 vssd1 vccd1 vccd1 _11892_/X sky130_fd_sc_hd__or3_1
XANTENNA__07350__A2 _07554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10843_ _10844_/A _10844_/B vssd1 vssd1 vccd1 vccd1 _10845_/A sky130_fd_sc_hd__and2_1
XANTENNA__09627__B2 _07830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09627__A1 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10774_ _10774_/A _10774_/B vssd1 vssd1 vccd1 vccd1 _10777_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_27_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12513_ reg1_val[8] curr_PC[8] _12520_/S vssd1 vssd1 vccd1 vccd1 _12515_/B sky130_fd_sc_hd__mux2_1
XANTENNA__12593__S _12638_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12444_ reg1_val[30] _12444_/B _12444_/C vssd1 vssd1 vccd1 vccd1 _12445_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12375_ _12449_/B1 _12414_/B hold258/A vssd1 vssd1 vccd1 vccd1 _12375_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__08602__A2 _08598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11326_ _11326_/A _11326_/B vssd1 vssd1 vccd1 vccd1 _11329_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11257_ hold275/A _11650_/B _11356_/B _12376_/C1 vssd1 vssd1 vccd1 vccd1 _11258_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_66_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11188_ _11189_/A _11189_/B vssd1 vssd1 vccd1 vccd1 _11190_/A sky130_fd_sc_hd__and2_1
X_10208_ fanout57/X fanout36/X fanout34/X fanout63/X vssd1 vssd1 vccd1 vccd1 _10209_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_66_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09407__S _11138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06977__D _07233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10139_ _09551_/X _09552_/X _10138_/C vssd1 vssd1 vccd1 vccd1 _10139_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09650__B _10476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07350_ _07134_/Y _07554_/B _07175_/A _07166_/Y vssd1 vssd1 vccd1 vccd1 _07351_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07629__B1 _07173_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08841__A2 _10245_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09020_ _08826_/A _08826_/B _08829_/A vssd1 vssd1 vccd1 vccd1 _09025_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_17_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07281_ _11381_/A _07281_/B vssd1 vssd1 vccd1 vccd1 _07287_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold202 hold202/A vssd1 vssd1 vccd1 vccd1 hold202/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold224 hold224/A vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 hold213/A vssd1 vssd1 vccd1 vccd1 hold213/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 hold235/A vssd1 vssd1 vccd1 vccd1 hold235/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold268 hold268/A vssd1 vssd1 vccd1 vccd1 hold268/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold246 hold246/A vssd1 vssd1 vccd1 vccd1 hold246/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 hold257/A vssd1 vssd1 vccd1 vccd1 hold257/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold279 hold279/A vssd1 vssd1 vccd1 vccd1 hold279/X sky130_fd_sc_hd__buf_1
X_09922_ _09922_/A _09922_/B vssd1 vssd1 vccd1 vccd1 _09923_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09853_ _09853_/A _09853_/B vssd1 vssd1 vccd1 vccd1 _09854_/B sky130_fd_sc_hd__xnor2_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11361__B1 _11995_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09784_ _09784_/A _09784_/B vssd1 vssd1 vccd1 vccd1 _09847_/A sky130_fd_sc_hd__xor2_4
X_08804_ _07817_/Y _08702_/B _08704_/Y vssd1 vssd1 vccd1 vccd1 _08807_/B sky130_fd_sc_hd__a21o_1
XANTENNA_fanout292_A _09218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06996_ _06995_/A _06987_/A _06987_/B _07094_/B vssd1 vssd1 vccd1 vccd1 _06998_/B
+ sky130_fd_sc_hd__a31o_2
X_08735_ _10668_/C _10668_/D _10668_/B vssd1 vssd1 vccd1 vccd1 _08735_/Y sky130_fd_sc_hd__a21oi_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08666_ _08666_/A _08666_/B vssd1 vssd1 vccd1 vccd1 _08717_/A sky130_fd_sc_hd__xnor2_1
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07361__A _12224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09609__A1 _09770_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08597_ _08596_/A _08596_/C _08596_/B vssd1 vssd1 vccd1 vccd1 _08603_/B sky130_fd_sc_hd__a21o_1
X_07617_ _10749_/A _07617_/B vssd1 vssd1 vccd1 vccd1 _07620_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07080__B _07080_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09609__B2 _07283_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07548_ _09341_/A _07548_/B vssd1 vssd1 vccd1 vccd1 _07708_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_119_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07479_ _07492_/B _07535_/A _07492_/A vssd1 vssd1 vccd1 vccd1 _07493_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_106_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10490_ _07198_/Y _08877_/B fanout6/X _10599_/A vssd1 vssd1 vccd1 vccd1 _10491_/B
+ sky130_fd_sc_hd__o22a_1
X_09218_ _09218_/A curr_PC[0] vssd1 vssd1 vccd1 vccd1 _09218_/X sky130_fd_sc_hd__or2_1
XFILLER_0_51_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08192__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09288__A _09944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10927__A0 _12420_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09149_ _09234_/C _09239_/B vssd1 vssd1 vccd1 vccd1 _09149_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_44_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12160_ _12161_/B _12160_/B vssd1 vssd1 vccd1 vccd1 _12235_/A sky130_fd_sc_hd__and2b_1
XANTENNA__09793__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11111_ _11111_/A _11111_/B vssd1 vssd1 vccd1 vccd1 _11113_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12091_ _12157_/A _12091_/B vssd1 vssd1 vccd1 vccd1 _12093_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11042_ _11247_/A _09575_/X _09251_/A vssd1 vssd1 vccd1 vccd1 _11042_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_99_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12993_ _13001_/A hold209/X vssd1 vssd1 vccd1 vccd1 hold210/A sky130_fd_sc_hd__and2_1
X_11944_ _12233_/B fanout23/X fanout15/X _12233_/A vssd1 vssd1 vccd1 vccd1 _11945_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10458__A2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11655__B2 _09221_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11655__A1 _12379_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11875_ _11876_/A _11876_/B vssd1 vssd1 vccd1 vccd1 _11962_/A sky130_fd_sc_hd__or2_1
XFILLER_0_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10826_ _10726_/A _10726_/B _10727_/Y vssd1 vssd1 vccd1 vccd1 _10838_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09076__A2 _10245_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10757_ _10758_/A _10758_/B vssd1 vssd1 vccd1 vccd1 _10759_/A sky130_fd_sc_hd__or2_1
XANTENNA__08823__A2 _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10688_ _09228_/X _09234_/X _10688_/S vssd1 vssd1 vccd1 vccd1 _10688_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10091__B1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12427_ _12050_/X _12306_/X _12398_/Y _12399_/X _11892_/A vssd1 vssd1 vccd1 vccd1
+ _12427_/X sky130_fd_sc_hd__a41o_1
XFILLER_0_124_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12358_ _06632_/B _12311_/Y _06630_/X vssd1 vssd1 vccd1 vccd1 _12358_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_50_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11309_ _11309_/A _12017_/A _11309_/C vssd1 vssd1 vccd1 vccd1 _11311_/A sky130_fd_sc_hd__or3_1
X_12289_ _12157_/A _07596_/A _12158_/B _12288_/X vssd1 vssd1 vccd1 vccd1 _12341_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06850_ _11349_/A _06848_/X _06849_/Y vssd1 vssd1 vccd1 vccd1 _06850_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06781_ _06781_/A _06781_/B vssd1 vssd1 vccd1 vccd1 _10155_/A sky130_fd_sc_hd__and2_1
XANTENNA__13096__B1 _13254_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08520_ _08522_/A _08522_/B vssd1 vssd1 vccd1 vccd1 _08521_/C sky130_fd_sc_hd__nand2b_1
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08451_ _08462_/A _08462_/B vssd1 vssd1 vccd1 vccd1 _08464_/A sky130_fd_sc_hd__nand2b_1
X_07402_ _07402_/A _07402_/B vssd1 vssd1 vccd1 vccd1 _07430_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12733__A2_N _07109_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08382_ _10207_/A _08382_/B vssd1 vssd1 vccd1 vccd1 _08408_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_128_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12071__A1 _11829_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07333_ fanout63/X _09943_/B2 _09650_/A fanout61/X vssd1 vssd1 vccd1 vccd1 _07334_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_116_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10082__B1 _10725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout138_A _09794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07264_ _10623_/A _07264_/B vssd1 vssd1 vccd1 vccd1 _07278_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09003_ _10871_/A fanout25/X _10974_/A _08112_/B vssd1 vssd1 vccd1 vccd1 _09004_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_26_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13020__B1 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07195_ _07195_/A _07195_/B vssd1 vssd1 vccd1 vccd1 _07195_/X sky130_fd_sc_hd__xor2_4
XANTENNA__11031__C1 _12446_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09836__A _09836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09905_ _09871_/Y _09873_/Y _09878_/X _09904_/X _06958_/A vssd1 vssd1 vccd1 vccd1
+ _09905_/X sky130_fd_sc_hd__o41a_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09836_ _09836_/A _09836_/B vssd1 vssd1 vccd1 vccd1 _09838_/B sky130_fd_sc_hd__xnor2_2
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06979_ _06983_/A _06983_/B vssd1 vssd1 vccd1 vccd1 _06979_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__06761__B1 _06760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ _09704_/A _09704_/B _09702_/X vssd1 vssd1 vccd1 vccd1 _09862_/A sky130_fd_sc_hd__a21oi_4
X_08718_ _09717_/B _09717_/C vssd1 vssd1 vccd1 vccd1 _08720_/A sky130_fd_sc_hd__nand2_1
X_09698_ _09539_/A _09539_/B _09537_/X vssd1 vssd1 vccd1 vccd1 _09699_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_95_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07091__A _10243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08649_ _09404_/S _08649_/A2 _08649_/B1 _08657_/B vssd1 vssd1 vccd1 vccd1 _08650_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ curr_PC[19] _11749_/C _11659_/Y vssd1 vssd1 vccd1 vccd1 _11660_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_49_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11591_ _11591_/A _11591_/B vssd1 vssd1 vccd1 vccd1 _11593_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_107_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10611_ _10611_/A _10611_/B vssd1 vssd1 vccd1 vccd1 _10612_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13330_ _13360_/CLK _13330_/D vssd1 vssd1 vccd1 vccd1 hold125/A sky130_fd_sc_hd__dfxtp_1
X_10542_ _10542_/A _10661_/A _10661_/B _10661_/C vssd1 vssd1 vccd1 vccd1 _10542_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13261_ hold3/X hold299/X _13260_/X _13259_/A vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__o211a_1
XANTENNA__08018__B1 _10338_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10473_ _10240_/A fanout12/X fanout7/X _10473_/B2 vssd1 vssd1 vccd1 vccd1 _10474_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12212_ _12129_/B _12129_/C _11892_/A vssd1 vssd1 vccd1 vccd1 _12212_/X sky130_fd_sc_hd__a21o_1
X_13192_ _13210_/A hold265/X vssd1 vssd1 vccd1 vccd1 _13379_/D sky130_fd_sc_hd__and2_1
XANTENNA__11995__B _11995_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08650__A _08658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12143_ _09228_/X _09234_/X _12143_/S vssd1 vssd1 vccd1 vccd1 _12143_/X sky130_fd_sc_hd__mux2_1
X_12074_ _12379_/B2 _10299_/X _12073_/X vssd1 vssd1 vccd1 vccd1 _12074_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07266__A _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11025_ _11025_/A _11025_/B vssd1 vssd1 vccd1 vccd1 _11027_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_99_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12976_ hold293/A _13000_/A2 _13257_/A2 hold243/X vssd1 vssd1 vccd1 vccd1 hold244/A
+ sky130_fd_sc_hd__a22o_1
X_11927_ _12096_/A _11927_/B vssd1 vssd1 vccd1 vccd1 _11929_/B sky130_fd_sc_hd__xor2_1
XANTENNA__10851__A2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11858_ _11935_/B _11858_/B vssd1 vssd1 vccd1 vccd1 _11860_/B sky130_fd_sc_hd__and2_1
X_11789_ _11790_/A _11790_/B vssd1 vssd1 vccd1 vccd1 _11881_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_117_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10809_ _12421_/A1 _10808_/X _06754_/B vssd1 vssd1 vccd1 vccd1 _10809_/X sky130_fd_sc_hd__a21o_1
XANTENNA_19 reg1_val[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10603__A2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13002__B1 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07480__B2 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07480__A1 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09757__B1 _12319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08560__A _08664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07951_ _07951_/A _07951_/B vssd1 vssd1 vccd1 vccd1 _07952_/B sky130_fd_sc_hd__and2_1
X_06902_ _06902_/A _06902_/B _06902_/C vssd1 vssd1 vccd1 vccd1 _06902_/X sky130_fd_sc_hd__and3_1
XFILLER_0_128_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07882_ _07842_/A _07841_/B _07841_/C vssd1 vssd1 vccd1 vccd1 _07885_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_128_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06833_ _07215_/A reg1_val[8] vssd1 vssd1 vccd1 vccd1 _06833_/X sky130_fd_sc_hd__and2b_1
X_09621_ _09621_/A _09621_/B _09621_/C vssd1 vssd1 vccd1 vccd1 _09622_/B sky130_fd_sc_hd__and3_1
X_06764_ reg1_val[9] _07237_/A vssd1 vssd1 vccd1 vccd1 _06765_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13117__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09552_ _09552_/A _09552_/B _09863_/A _10004_/A vssd1 vssd1 vccd1 vccd1 _09552_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_78_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08503_ _08641_/B _08561_/A2 _08561_/B1 _08627_/A2 vssd1 vssd1 vccd1 vccd1 _08504_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_93_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06695_ reg2_val[21] _06766_/B _06724_/B1 _06694_/Y vssd1 vssd1 vccd1 vccd1 _06984_/B
+ sky130_fd_sc_hd__o2bb2a_2
XANTENNA_fanout255_A _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09483_ _09484_/A _09484_/B vssd1 vssd1 vccd1 vccd1 _09485_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_92_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08434_ _08434_/A _08434_/B vssd1 vssd1 vccd1 vccd1 _08757_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08365_ _08365_/A _08365_/B vssd1 vssd1 vccd1 vccd1 _08400_/B sky130_fd_sc_hd__xnor2_2
X_07316_ _10476_/B _10476_/C vssd1 vssd1 vccd1 vccd1 _07316_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_34_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08296_ _08297_/A _08297_/B vssd1 vssd1 vccd1 vccd1 _08296_/X sky130_fd_sc_hd__or2_1
XFILLER_0_33_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07247_ _10207_/A vssd1 vssd1 vccd1 vccd1 _10950_/A sky130_fd_sc_hd__inv_6
XFILLER_0_14_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07178_ _07371_/A _07371_/B vssd1 vssd1 vccd1 vccd1 _07372_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_112_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07223__A1 _07959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07223__B2 _12823_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08971__A1 _09298_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08971__B2 _09298_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout70_A _09936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09819_ _09819_/A _09819_/B vssd1 vssd1 vccd1 vccd1 _09820_/B sky130_fd_sc_hd__nor2_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12830_ hold85/X _12862_/B vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__or2_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10240__A _10240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12761_ _12742_/B _12760_/X _12755_/B _07143_/A vssd1 vssd1 vccd1 vccd1 _12763_/B
+ sky130_fd_sc_hd__a2bb2o_2
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _11712_/A _11885_/A vssd1 vssd1 vccd1 vccd1 _11716_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_83_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _12693_/A _12693_/C _12693_/B vssd1 vssd1 vccd1 vccd1 _12699_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_127_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11643_ _12444_/B _11643_/B vssd1 vssd1 vccd1 vccd1 _11643_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_83_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11574_ _11689_/A _11574_/B vssd1 vssd1 vccd1 vccd1 _11578_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_92_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13313_ _13316_/CLK _13313_/D vssd1 vssd1 vccd1 vccd1 hold204/A sky130_fd_sc_hd__dfxtp_1
X_10525_ _10525_/A _10525_/B vssd1 vssd1 vccd1 vccd1 _10527_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_24_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13244_ hold258/A _13243_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13244_/X sky130_fd_sc_hd__mux2_1
X_10456_ _12233_/B _08289_/B fanout74/X _12233_/A vssd1 vssd1 vccd1 vccd1 _10457_/B
+ sky130_fd_sc_hd__o22a_1
X_13175_ hold272/X _13174_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13175_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_110_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12126_ _06672_/A _12125_/X _11637_/A vssd1 vssd1 vccd1 vccd1 _12126_/Y sky130_fd_sc_hd__a21oi_1
X_10387_ _11770_/A _10387_/B vssd1 vssd1 vccd1 vccd1 _10389_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10415__A _10415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08962__A1 _08199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08962__B2 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12057_ _10049_/A _08795_/A _08795_/B vssd1 vssd1 vccd1 vccd1 _12057_/Y sky130_fd_sc_hd__a21oi_1
X_11008_ _11008_/A _11120_/A vssd1 vssd1 vccd1 vccd1 _11229_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07724__A _09341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06725__B1 _06783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12959_ _13216_/A _12958_/B _12882_/X vssd1 vssd1 vccd1 vccd1 _13221_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_90_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06740__A3 _12714_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08150_ _08150_/A _08150_/B vssd1 vssd1 vccd1 vccd1 _08220_/B sky130_fd_sc_hd__xnor2_1
X_07101_ _07442_/A _07442_/B vssd1 vssd1 vccd1 vccd1 _07443_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_15_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08081_ _08081_/A _08081_/B vssd1 vssd1 vccd1 vccd1 _08082_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_113_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07032_ _06995_/A _06994_/X _06995_/Y _06987_/Y vssd1 vssd1 vccd1 vccd1 _07032_/Y
+ sky130_fd_sc_hd__a22oi_4
XANTENNA__12329__A2 _09732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08290__A _08334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10325__A _10581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08983_ _08983_/A _08983_/B vssd1 vssd1 vccd1 vccd1 _08984_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07934_ _07934_/A _07934_/B vssd1 vssd1 vccd1 vccd1 _07941_/B sky130_fd_sc_hd__xor2_4
XANTENNA__07508__A2 _08484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07865_ _07872_/A _07872_/B vssd1 vssd1 vccd1 vccd1 _07946_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_98_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10512__B2 _11476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10512__A1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09604_ _11752_/S _09603_/Y _09444_/X vssd1 vssd1 vccd1 vccd1 dest_val[2] sky130_fd_sc_hd__o21ai_4
XFILLER_0_97_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06816_ reg2_val[0] _06766_/B _06817_/B1 _06815_/X vssd1 vssd1 vccd1 vccd1 _09103_/A
+ sky130_fd_sc_hd__a22oi_4
X_07796_ _09341_/A _07796_/B vssd1 vssd1 vccd1 vccd1 _07823_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__11068__A2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12265__A1 _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06747_ reg1_val[12] _07195_/A vssd1 vssd1 vccd1 vccd1 _06748_/B sky130_fd_sc_hd__nor2_1
X_09535_ _09336_/A _09334_/Y _09333_/X vssd1 vssd1 vccd1 vccd1 _09538_/A sky130_fd_sc_hd__a21bo_1
X_06678_ _07036_/A reg1_val[23] vssd1 vssd1 vccd1 vccd1 _11995_/A sky130_fd_sc_hd__and2b_1
X_09466_ _09347_/A _09347_/B _09344_/A vssd1 vssd1 vccd1 vccd1 _09469_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_109_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08417_ _08649_/A2 _10221_/B2 _08501_/B1 _08657_/B vssd1 vssd1 vccd1 vccd1 _08418_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_108_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09397_ _09193_/X _09195_/X _09419_/B vssd1 vssd1 vccd1 vccd1 _09397_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10579__A1 _12356_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08348_ _08355_/B _08355_/A vssd1 vssd1 vccd1 vccd1 _08357_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__07444__A1 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07444__B2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08279_ _08280_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08279_/Y sky130_fd_sc_hd__nor2_1
X_11290_ _11291_/A _11291_/B vssd1 vssd1 vccd1 vccd1 _11417_/B sky130_fd_sc_hd__nor2_1
X_10310_ reg1_val[7] curr_PC[7] vssd1 vssd1 vccd1 vccd1 _10310_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__06798__A3 _12660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10241_ _10242_/B _10242_/C _08454_/A vssd1 vssd1 vccd1 vccd1 _10243_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_14_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10235__A _12224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ hold260/A _09425_/C _10303_/B _10171_/Y _12416_/C1 vssd1 vssd1 vccd1 vccd1
+ _10172_/Y sky130_fd_sc_hd__a311oi_1
XFILLER_0_30_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout183 _06969_/Y vssd1 vssd1 vccd1 vccd1 _07094_/B sky130_fd_sc_hd__buf_6
Xfanout172 _12826_/B vssd1 vssd1 vccd1 vccd1 _12820_/B sky130_fd_sc_hd__buf_4
Xfanout161 _11538_/A vssd1 vssd1 vccd1 vccd1 _11809_/A sky130_fd_sc_hd__buf_4
Xfanout150 _07037_/X vssd1 vssd1 vccd1 vccd1 _09298_/A1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07544__A _09836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout194 _12205_/B1 vssd1 vssd1 vccd1 vccd1 _11648_/A sky130_fd_sc_hd__buf_4
XANTENNA__07380__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12813_ _07173_/Y _13101_/B2 hold71/X _13147_/A vssd1 vssd1 vccd1 vccd1 _13267_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ reg1_val[21] _12755_/B vssd1 vssd1 vccd1 vccd1 _12744_/Y sky130_fd_sc_hd__nor2_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07132__B1 _07117_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ reg1_val[7] _12675_/B vssd1 vssd1 vccd1 vccd1 _12676_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07683__A1 fanout72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07683__B2 _10595_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11626_ _11841_/A vssd1 vssd1 vccd1 vccd1 _11626_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_37_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11557_ hold177/A _11557_/B vssd1 vssd1 vccd1 vccd1 _11645_/B sky130_fd_sc_hd__or2_1
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10508_ _11770_/A _10508_/B vssd1 vssd1 vccd1 vccd1 _10510_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07986__A2 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07719__A _08334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11488_ _12233_/B fanout45/X fanout17/X fanout47/X vssd1 vssd1 vccd1 vccd1 _11489_/B
+ sky130_fd_sc_hd__o22a_1
X_13227_ hold284/X _13248_/B1 _13226_/X _13248_/A2 vssd1 vssd1 vccd1 vccd1 _13228_/B
+ sky130_fd_sc_hd__a22o_1
X_10439_ _09425_/C _10438_/X hold252/A vssd1 vssd1 vccd1 vccd1 _10439_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13158_ _13158_/A _13158_/B vssd1 vssd1 vccd1 vccd1 _13159_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09934__A _09934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08935__B2 _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08935__A1 _07554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12109_ _12177_/B _12109_/B vssd1 vssd1 vccd1 vccd1 _12111_/C sky130_fd_sc_hd__nand2_1
X_13089_ _09922_/A _13089_/A2 hold76/X vssd1 vssd1 vccd1 vccd1 _13354_/D sky130_fd_sc_hd__o21a_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07650_ _09667_/A _07650_/B vssd1 vssd1 vccd1 vccd1 _07652_/B sky130_fd_sc_hd__xnor2_1
X_06601_ instruction[22] _06944_/B vssd1 vssd1 vccd1 vccd1 _06601_/X sky130_fd_sc_hd__or2_1
XFILLER_0_88_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07581_ _07581_/A _07581_/B vssd1 vssd1 vccd1 vccd1 _07584_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_19_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09320_ _09321_/A _09321_/B vssd1 vssd1 vccd1 vccd1 _09463_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_118_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09251_ _09251_/A _11247_/B _11247_/C vssd1 vssd1 vccd1 vccd1 _12445_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_56_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08202_ _09940_/B2 _08484_/B _09479_/B1 _08561_/A2 vssd1 vssd1 vccd1 vccd1 _08203_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_90_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09182_ _09178_/X _09181_/X _09727_/S vssd1 vssd1 vccd1 vccd1 _09182_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11758__B1 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout120_A _07194_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08133_ _08215_/A _08215_/B _08125_/X vssd1 vssd1 vccd1 vccd1 _08153_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_28_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12535__A _12696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13130__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout218_A _07149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08064_ _08064_/A _08064_/B _08064_/C vssd1 vssd1 vccd1 vccd1 _08068_/A sky130_fd_sc_hd__and3_1
XANTENNA__07977__A2 _10595_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07015_ _07011_/A _07011_/B _09302_/A vssd1 vssd1 vccd1 vccd1 _07015_/X sky130_fd_sc_hd__mux2_2
XANTENNA__11930__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08966_ fanout98/X fanout78/X fanout74/X fanout84/X vssd1 vssd1 vccd1 vccd1 _08967_/B
+ sky130_fd_sc_hd__o22a_1
X_07917_ _07913_/A _07913_/B _07913_/C vssd1 vssd1 vccd1 vccd1 _07917_/X sky130_fd_sc_hd__a21o_1
X_08897_ _08898_/A _08898_/B vssd1 vssd1 vccd1 vccd1 _08899_/A sky130_fd_sc_hd__and2_1
X_07848_ _09943_/B2 fanout80/X fanout76/X _08538_/A1 vssd1 vssd1 vccd1 vccd1 _07849_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09518_ _09518_/A _09518_/B vssd1 vssd1 vccd1 vccd1 _09519_/B sky130_fd_sc_hd__nor2_1
X_07779_ _08575_/A _07779_/B vssd1 vssd1 vccd1 vccd1 _07845_/B sky130_fd_sc_hd__xor2_1
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10790_ _10672_/A _10670_/Y _10688_/S vssd1 vssd1 vccd1 vccd1 _10791_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_66_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout33_A _07201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08195__A _08580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _09936_/A _09449_/B vssd1 vssd1 vccd1 vccd1 _09453_/B sky130_fd_sc_hd__xnor2_1
X_12460_ _09218_/A curr_PC[0] _12520_/S vssd1 vssd1 vccd1 vccd1 _12462_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11411_ _11410_/A _11410_/B _11410_/C vssd1 vssd1 vccd1 vccd1 _11412_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_117_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12391_ _12391_/A _12391_/B _12391_/C vssd1 vssd1 vccd1 vccd1 _12394_/A sky130_fd_sc_hd__and3_1
XFILLER_0_46_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08614__B1 _09672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11342_ _11272_/X _11567_/B _12356_/B1 vssd1 vssd1 vccd1 vccd1 _11342_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11273_ _11193_/A _11193_/B _11190_/A vssd1 vssd1 vccd1 vccd1 _11282_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13012_ hold180/X _13171_/B2 _13209_/A2 hold172/X vssd1 vssd1 vccd1 vccd1 hold181/A
+ sky130_fd_sc_hd__a22o_1
X_10224_ _10224_/A _10224_/B vssd1 vssd1 vccd1 vccd1 _10225_/C sky130_fd_sc_hd__xor2_1
X_10155_ _10155_/A _10155_/B vssd1 vssd1 vccd1 vccd1 _10155_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07274__A _11038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10086_ _10086_/A _10086_/B vssd1 vssd1 vccd1 vccd1 _10088_/B sky130_fd_sc_hd__xor2_2
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10488__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10988_ _10886_/A _10886_/B _10884_/Y vssd1 vssd1 vccd1 vccd1 _10997_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_97_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12727_ reg1_val[16] _12755_/B _12739_/A vssd1 vssd1 vccd1 vccd1 _12729_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_38_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12658_ _12657_/A _12654_/Y _12656_/B vssd1 vssd1 vccd1 vccd1 _12662_/A sky130_fd_sc_hd__o21a_2
X_11609_ _11609_/A _11609_/B vssd1 vssd1 vccd1 vccd1 _11610_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07408__B2 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07408__A1 _09298_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12589_ _12633_/A _12589_/B vssd1 vssd1 vccd1 vccd1 _12590_/B sky130_fd_sc_hd__or2_1
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap103 _06701_/A vssd1 vssd1 vccd1 vccd1 _06902_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11912__B1 _12376_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _08821_/A _08821_/B vssd1 vssd1 vccd1 vccd1 _08822_/A sky130_fd_sc_hd__and2_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06800__B _07165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ _08751_/A _08751_/B _08751_/C vssd1 vssd1 vccd1 vccd1 _08751_/X sky130_fd_sc_hd__or3_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08682_ _08739_/A _08549_/X _08683_/A vssd1 vssd1 vccd1 vccd1 _08682_/Y sky130_fd_sc_hd__a21oi_1
X_07702_ _07784_/A _07784_/B _07698_/X vssd1 vssd1 vccd1 vccd1 _07804_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__08136__A2 _10595_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07912__A _09302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07633_ _07634_/A _07634_/B vssd1 vssd1 vccd1 vccd1 _08893_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07344__B1 _07173_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout168_A _12805_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13125__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07564_ _07565_/A _07565_/B vssd1 vssd1 vccd1 vccd1 _07564_/Y sky130_fd_sc_hd__nand2_1
X_09303_ _09302_/B _09302_/C _09302_/A vssd1 vssd1 vccd1 vccd1 _09306_/C sky130_fd_sc_hd__a21o_1
XANTENNA__11443__A2 _11840_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07647__A1 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07647__B2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07495_ _07495_/A _07495_/B vssd1 vssd1 vccd1 vccd1 _07561_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_118_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09234_ instruction[6] _09234_/B _09234_/C vssd1 vssd1 vccd1 vccd1 _09234_/X sky130_fd_sc_hd__or3_4
XFILLER_0_61_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13196__A2 _13223_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09165_ reg1_val[7] reg1_val[24] _09180_/S vssd1 vssd1 vccd1 vccd1 _09165_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08116_ _08116_/A _08116_/B vssd1 vssd1 vccd1 vccd1 _08121_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_16_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09096_ _09097_/A _09097_/B vssd1 vssd1 vccd1 vccd1 _09330_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08047_ _08099_/A _08099_/B _08043_/X vssd1 vssd1 vccd1 vccd1 _08051_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12156__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10513__A _11929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06710__B _12655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ _09998_/A _09998_/B vssd1 vssd1 vccd1 vccd1 _09999_/B sky130_fd_sc_hd__xnor2_4
X_08949_ fanout61/X _10473_/B2 _10240_/A fanout53/X vssd1 vssd1 vccd1 vccd1 _08950_/B
+ sky130_fd_sc_hd__o22a_1
X_11960_ _12040_/B _11960_/B vssd1 vssd1 vccd1 vccd1 _11962_/C sky130_fd_sc_hd__nand2_1
X_10911_ _06897_/D _10910_/X _11637_/A vssd1 vssd1 vccd1 vccd1 _10911_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11682__A2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11891_ _11892_/A _11892_/B _12049_/A vssd1 vssd1 vccd1 vccd1 _11891_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10842_ _11929_/A _10842_/B vssd1 vssd1 vccd1 vccd1 _10844_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09627__A2 _10871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10773_ _10774_/B _10774_/A vssd1 vssd1 vccd1 vccd1 _10897_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08835__B1 _10240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12512_ _12518_/B _12512_/B vssd1 vssd1 vccd1 vccd1 new_PC[7] sky130_fd_sc_hd__and2_4
XFILLER_0_26_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12443_ _12364_/A _08924_/X _09040_/D _12365_/A vssd1 vssd1 vccd1 vccd1 _12443_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_50_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12374_ hold287/A _12374_/B vssd1 vssd1 vccd1 vccd1 _12414_/B sky130_fd_sc_hd__or2_1
XANTENNA__07269__A _07270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11325_ _11326_/A _11326_/B vssd1 vssd1 vccd1 vccd1 _11431_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_50_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11256_ _11650_/B _11356_/B hold275/A vssd1 vssd1 vccd1 vccd1 _11258_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11187_ _11770_/A _11187_/B vssd1 vssd1 vccd1 vccd1 _11189_/B sky130_fd_sc_hd__xnor2_1
X_10207_ _10207_/A _10207_/B vssd1 vssd1 vccd1 vccd1 _10211_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10173__A2 _12422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11370__A1 _12365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10138_ _10138_/A _10138_/B _10138_/C vssd1 vssd1 vccd1 vccd1 _10138_/X sky130_fd_sc_hd__or3_1
XANTENNA__06782__D1 _06927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10069_ _10069_/A _10069_/B vssd1 vssd1 vccd1 vccd1 _10077_/A sky130_fd_sc_hd__xor2_2
XANTENNA__11658__C1 _11657_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07326__B1 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09650__C _10476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11254__A _11648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07629__B2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07629__A1 _07417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07280_ _07191_/X _10725_/A _07202_/Y _07232_/X vssd1 vssd1 vccd1 vccd1 _07281_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11830__C1 _12421_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold225 hold225/A vssd1 vssd1 vccd1 vccd1 hold225/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold203 hold203/A vssd1 vssd1 vccd1 vccd1 hold203/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 hold214/A vssd1 vssd1 vccd1 vccd1 hold214/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold269 hold269/A vssd1 vssd1 vccd1 vccd1 hold269/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12138__B1 _12416_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold258 hold258/A vssd1 vssd1 vccd1 vccd1 hold258/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold247 hold247/A vssd1 vssd1 vccd1 vccd1 hold247/X sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _07175_/A _10234_/A2 _07274_/Y _07554_/B vssd1 vssd1 vccd1 vccd1 _09922_/B
+ sky130_fd_sc_hd__a22o_1
Xhold236 hold236/A vssd1 vssd1 vccd1 vccd1 hold236/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07907__A _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09003__B1 _10974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11361__A1 _06727_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09852_ _09850_/A _09850_/B _09853_/B vssd1 vssd1 vccd1 vccd1 _09852_/Y sky130_fd_sc_hd__a21oi_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _09783_/A _09783_/B vssd1 vssd1 vccd1 vccd1 _09784_/B sky130_fd_sc_hd__nor2_2
X_08803_ _12258_/B _12258_/C vssd1 vssd1 vccd1 vccd1 _09040_/A sky130_fd_sc_hd__and2_2
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06995_ _06995_/A _07094_/B vssd1 vssd1 vccd1 vccd1 _06995_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout285_A _12404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08734_ _08733_/A _08733_/C _08733_/B vssd1 vssd1 vccd1 vccd1 _10668_/D sky130_fd_sc_hd__a21o_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12861__A1 _12169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08665_ _08665_/A _08665_/B vssd1 vssd1 vccd1 vccd1 _08666_/B sky130_fd_sc_hd__xor2_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09609__A2 _07362_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08596_ _08596_/A _08596_/B _08596_/C vssd1 vssd1 vccd1 vccd1 _08603_/A sky130_fd_sc_hd__nand3_1
X_07616_ fanout51/X _10473_/B2 _10240_/A _09661_/B2 vssd1 vssd1 vccd1 vccd1 _07617_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_119_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07547_ _09934_/A fanout25/X _07283_/X _08112_/B vssd1 vssd1 vccd1 vccd1 _07548_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10624__B1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11821__C1 _09242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12707__B _12708_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07478_ _07534_/A _07534_/B vssd1 vssd1 vccd1 vccd1 _07535_/A sky130_fd_sc_hd__and2_1
XANTENNA__08473__A _08564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10508__A _11770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09217_ _09218_/A curr_PC[0] vssd1 vssd1 vccd1 vccd1 _09413_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_106_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12377__B1 _12421_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09148_ _10049_/A _10321_/A _10321_/B vssd1 vssd1 vccd1 vccd1 _09148_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10927__A1 _09422_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09793__A1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09793__B2 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09079_ _09079_/A _09079_/B vssd1 vssd1 vccd1 vccd1 _09102_/A sky130_fd_sc_hd__xnor2_2
X_11110_ _11111_/B _11111_/A vssd1 vssd1 vccd1 vccd1 _11110_/Y sky130_fd_sc_hd__nand2b_1
X_12090_ fanout17/X fanout15/X _12335_/A fanout23/X vssd1 vssd1 vccd1 vccd1 _12091_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11339__A _11526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11041_ _11036_/Y _11037_/X _11038_/Y _11040_/X vssd1 vssd1 vccd1 vccd1 _11041_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10243__A _10243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11058__B _11058_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12992_ hold217/A _13000_/A2 _13257_/A2 hold208/X vssd1 vssd1 vccd1 vccd1 hold209/A
+ sky130_fd_sc_hd__a22o_1
X_11943_ _12009_/B _11943_/B vssd1 vssd1 vccd1 vccd1 _11950_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11074__A _12096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11874_ _11874_/A _11874_/B vssd1 vssd1 vccd1 vccd1 _11876_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10825_ _10768_/A _10768_/B _10769_/Y vssd1 vssd1 vccd1 vccd1 _10894_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10756_ _10756_/A _10756_/B vssd1 vssd1 vccd1 vccd1 _10758_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09481__B1 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10687_ hold213/A _11990_/A1 _10805_/B _12205_/B1 vssd1 vssd1 vccd1 vccd1 _10687_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_70_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10091__A1 _11868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10091__B2 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12368__B1 _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12426_ _08973_/C _06961_/X _12402_/Y _12425_/X _12631_/S vssd1 vssd1 vccd1 vccd1
+ dest_val[30] sky130_fd_sc_hd__o221a_4
XFILLER_0_35_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12357_ _12399_/B _12355_/X _12356_/Y vssd1 vssd1 vccd1 vccd1 _12357_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07795__B1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11308_ _11308_/A _11308_/B vssd1 vssd1 vccd1 vccd1 _11309_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12288_ fanout15/X fanout7/X _11844_/A vssd1 vssd1 vccd1 vccd1 _12288_/X sky130_fd_sc_hd__o21a_1
X_11239_ _11239_/A _11239_/B vssd1 vssd1 vccd1 vccd1 _11239_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11249__A _11820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07547__B1 _07283_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06780_ reg1_val[6] _07283_/A vssd1 vssd1 vccd1 vccd1 _06781_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12843__A1 _07097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08450_ _08450_/A _08450_/B vssd1 vssd1 vccd1 vccd1 _08462_/B sky130_fd_sc_hd__nand2_1
X_07401_ _07401_/A _07401_/B vssd1 vssd1 vccd1 vccd1 _07402_/B sky130_fd_sc_hd__nor2_2
X_08381_ _08649_/B1 _08411_/B _10476_/A _09404_/S vssd1 vssd1 vccd1 vccd1 _08382_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12808__A _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07332_ _10749_/A _07332_/B vssd1 vssd1 vccd1 vccd1 _07336_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08293__A _08664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10082__A1 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10082__B2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07263_ fanout86/X fanout84/X fanout82/X fanout80/X vssd1 vssd1 vccd1 vccd1 _07264_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_116_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07194_ _07195_/A _07195_/B vssd1 vssd1 vccd1 vccd1 _07194_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_5_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09002_ _08825_/A _08825_/B _08822_/A vssd1 vssd1 vccd1 vccd1 _09014_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_26_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12543__A _12702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout200_A _09149_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07637__A _09922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09904_ _12379_/B2 _09880_/Y _09886_/X _09887_/X _09903_/Y vssd1 vssd1 vccd1 vccd1
+ _09904_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_1_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09835_ _07959_/B _07256_/Y _07262_/X fanout29/X vssd1 vssd1 vccd1 vccd1 _09836_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06978_ _07262_/A _07270_/A _06978_/C _06978_/D vssd1 vssd1 vccd1 vccd1 _06983_/B
+ sky130_fd_sc_hd__nor4_4
X_09766_ _12364_/A _09909_/A vssd1 vssd1 vccd1 vccd1 _09766_/X sky130_fd_sc_hd__or2_1
XFILLER_0_68_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08717_ _08717_/A _08717_/B vssd1 vssd1 vccd1 vccd1 _09717_/C sky130_fd_sc_hd__xor2_1
X_09697_ _09697_/A _09697_/B vssd1 vssd1 vccd1 vccd1 _09699_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ _08656_/A _08648_/B vssd1 vssd1 vccd1 vccd1 _08665_/A sky130_fd_sc_hd__xnor2_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08579_ _12808_/A _09650_/A _09325_/A _09943_/B2 vssd1 vssd1 vccd1 vccd1 _08580_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11590_ _11591_/A _11591_/B vssd1 vssd1 vccd1 vccd1 _11590_/Y sky130_fd_sc_hd__nand2_1
X_10610_ _10611_/A _10611_/B vssd1 vssd1 vccd1 vccd1 _10610_/Y sky130_fd_sc_hd__nand2_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09299__A _09673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06816__A2 _06766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10073__B2 _10243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10541_ _10541_/A _10780_/A vssd1 vssd1 vccd1 vccd1 _10541_/X sky130_fd_sc_hd__and2_1
XFILLER_0_36_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13260_ hold3/X _12803_/B hold68/A _12804_/A vssd1 vssd1 vccd1 vccd1 _13260_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_52_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08018__A1 _08598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12211_ _12211_/A _12211_/B _12211_/C _12211_/D vssd1 vssd1 vccd1 vccd1 _12215_/C
+ sky130_fd_sc_hd__or4_1
X_10472_ _10393_/A _10393_/B _10390_/A vssd1 vssd1 vccd1 vccd1 _10487_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08018__B2 _08538_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08931__A _09779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13191_ hold264/X _13223_/A2 _13190_/X _13223_/B2 vssd1 vssd1 vccd1 vccd1 hold265/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12142_ _13322_/Q _12447_/B1 _12203_/B _12205_/B1 vssd1 vssd1 vccd1 vccd1 _12142_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11069__A _11770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12073_ _06658_/B _12422_/A _09221_/Y _10293_/X _12072_/X vssd1 vssd1 vccd1 vccd1
+ _12073_/X sky130_fd_sc_hd__a221o_1
XANTENNA__07266__B _07267_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11024_ reg1_val[13] curr_PC[13] vssd1 vssd1 vccd1 vccd1 _11025_/B sky130_fd_sc_hd__or2_1
XANTENNA__11089__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12825__A1 _10337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12975_ _13001_/A _12975_/B vssd1 vssd1 vccd1 vccd1 _13297_/D sky130_fd_sc_hd__and2_1
X_11926_ fanout41/X _07316_/Y _07608_/Y fanout43/X vssd1 vssd1 vccd1 vccd1 _11927_/B
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_2_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13304_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11857_ _11857_/A _11857_/B vssd1 vssd1 vccd1 vccd1 _11858_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11788_ _11788_/A _11788_/B vssd1 vssd1 vccd1 vccd1 _11790_/B sky130_fd_sc_hd__xnor2_1
X_10808_ _12420_/A0 _09422_/B _10808_/S vssd1 vssd1 vccd1 vccd1 _10808_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_55_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10739_ _10739_/A _10739_/B vssd1 vssd1 vccd1 vccd1 _10740_/B sky130_fd_sc_hd__or2_1
XFILLER_0_82_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09757__A1 _09221_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07480__A2 _09298_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13389_ _13390_/CLK _13389_/D vssd1 vssd1 vccd1 vccd1 hold287/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09757__B2 _12379_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12409_ _09040_/C _12408_/X _10788_/A vssd1 vssd1 vccd1 vccd1 _12409_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07768__B1 _09325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07457__A _09947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07950_ _07948_/X _07950_/B vssd1 vssd1 vccd1 vccd1 _08711_/A sky130_fd_sc_hd__nand2b_2
X_06901_ _11349_/A _06901_/B _06901_/C _06901_/D vssd1 vssd1 vccd1 vccd1 _06902_/C
+ sky130_fd_sc_hd__and4b_1
XANTENNA__09672__A _09672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12810__B _12820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07881_ _07944_/A _07944_/B vssd1 vssd1 vccd1 vccd1 _07948_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_128_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06832_ _10291_/A _06830_/Y _06831_/X vssd1 vssd1 vccd1 vccd1 _06832_/X sky130_fd_sc_hd__a21o_1
XANTENNA__13069__A1 _09667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09620_ _09621_/A _09621_/B _09621_/C vssd1 vssd1 vccd1 vccd1 _09622_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__08288__A _10207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06763_ reg1_val[9] _07237_/A vssd1 vssd1 vccd1 vccd1 _06763_/Y sky130_fd_sc_hd__nor2_1
X_09551_ _09371_/A _09371_/B _09550_/Y vssd1 vssd1 vccd1 vccd1 _09551_/X sky130_fd_sc_hd__a21bo_1
X_08502_ _08502_/A _08502_/B vssd1 vssd1 vccd1 vccd1 _08506_/A sky130_fd_sc_hd__xnor2_1
X_06694_ _06703_/A _12670_/B vssd1 vssd1 vccd1 vccd1 _06694_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_77_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09482_ _09944_/A _09482_/B vssd1 vssd1 vccd1 vccd1 _09484_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08433_ _08403_/X _08433_/B vssd1 vssd1 vccd1 vccd1 _08759_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_92_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout248_A _12218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09445__B1 _10049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08364_ _08364_/A _08364_/B vssd1 vssd1 vccd1 vccd1 _08400_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_128_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07315_ _07315_/A _07315_/B vssd1 vssd1 vccd1 vccd1 _10476_/C sky130_fd_sc_hd__nor2_8
XFILLER_0_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10058__A _10950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08295_ _09670_/A _08295_/B vssd1 vssd1 vccd1 vccd1 _08297_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07246_ reg1_val[13] _07246_/B vssd1 vssd1 vccd1 vccd1 _09794_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__09748__A1 _12322_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07177_ _09922_/A _07177_/B vssd1 vssd1 vccd1 vccd1 _07371_/B sky130_fd_sc_hd__xor2_1
XANTENNA__07223__A2 _10337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08971__A2 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09818_ _09819_/A _09819_/B vssd1 vssd1 vccd1 vccd1 _09820_/A sky130_fd_sc_hd__and2_1
XANTENNA__12807__A1 _12428_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout63_A _07014_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09749_ hold221/A _12322_/A1 _09747_/X _12205_/B1 vssd1 vssd1 vccd1 vccd1 _09749_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10240__B _10476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12760_ _12760_/A _12760_/B _12760_/C _12760_/D vssd1 vssd1 vccd1 vccd1 _12760_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__08487__A1 _08454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _11711_/A _11799_/A vssd1 vssd1 vccd1 vccd1 _11885_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _12687_/A _12691_/B vssd1 vssd1 vccd1 vccd1 _12693_/C sky130_fd_sc_hd__nand2b_1
XANTENNA__07830__A _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11642_ _11642_/A _11642_/B vssd1 vssd1 vccd1 vccd1 _11642_/Y sky130_fd_sc_hd__xnor2_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11573_ _11572_/B _11573_/B vssd1 vssd1 vccd1 vccd1 _11574_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_107_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13312_ _13316_/CLK hold184/X vssd1 vssd1 vccd1 vccd1 hold182/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10524_ _10468_/B _10344_/B _10368_/B _10367_/B _10367_/A vssd1 vssd1 vccd1 vccd1
+ _10527_/A sky130_fd_sc_hd__a32o_1
X_13243_ _13243_/A _13243_/B vssd1 vssd1 vccd1 vccd1 _13243_/Y sky130_fd_sc_hd__xnor2_1
X_10455_ _10356_/A _10356_/B _10354_/Y vssd1 vssd1 vccd1 vccd1 _10471_/A sky130_fd_sc_hd__a21o_1
XANTENNA__08380__B _08384_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13174_ _13174_/A _13174_/B vssd1 vssd1 vccd1 vccd1 _13174_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10349__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12125_ _06882_/X _12124_/X _12404_/S vssd1 vssd1 vccd1 vccd1 _12125_/X sky130_fd_sc_hd__mux2_1
X_10386_ _11764_/A fanout32/X fanout30/X _11592_/A vssd1 vssd1 vccd1 vccd1 _10387_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10415__B _10415_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08962__A2 _11198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12056_ _06672_/B _12054_/X _12055_/Y vssd1 vssd1 vccd1 vccd1 _12056_/X sky130_fd_sc_hd__o21a_1
XANTENNA__09492__A _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11007_ _11007_/A _11007_/B vssd1 vssd1 vccd1 vccd1 _11227_/A sky130_fd_sc_hd__or2_4
XFILLER_0_74_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07922__B1 _09479_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12958_ _12882_/X _12958_/B vssd1 vssd1 vccd1 vccd1 _13216_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__12274__A2 _09257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08836__A _10749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12889_ hold246/X hold121/X vssd1 vssd1 vccd1 vccd1 _13188_/B sky130_fd_sc_hd__nand2b_1
X_11909_ hold219/A _12447_/B1 _11989_/B _11648_/A vssd1 vssd1 vccd1 vccd1 _11909_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__07150__A1 _11134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13223__B2 _13223_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07989__B1 _07256_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07100_ _10479_/A _07100_/B vssd1 vssd1 vccd1 vccd1 _07442_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12982__B1 _13257_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09667__A _09667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08080_ _08065_/B _08027_/C _08027_/B vssd1 vssd1 vccd1 vccd1 _08083_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12093__A _12093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07031_ _07031_/A _07031_/B vssd1 vssd1 vccd1 vccd1 _07031_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_2_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07187__A _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06803__B _06810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10325__B _10581_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_699 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08982_ _08982_/A _08982_/B vssd1 vssd1 vccd1 vccd1 _08983_/B sky130_fd_sc_hd__xor2_4
XANTENNA__07915__A _09673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07933_ _07956_/A _07956_/B _07901_/Y vssd1 vssd1 vccd1 vccd1 _07941_/A sky130_fd_sc_hd__a21o_2
XANTENNA_fanout198_A _12144_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07864_ _07934_/A _07934_/B _07844_/Y vssd1 vssd1 vccd1 vccd1 _07872_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__10512__A2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06815_ _06815_/A _12645_/B vssd1 vssd1 vccd1 vccd1 _06815_/X sky130_fd_sc_hd__and2_1
X_09603_ _12365_/A _09557_/X _09602_/X vssd1 vssd1 vccd1 vccd1 _09603_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_78_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07795_ _08561_/B1 _08112_/B fanout25/X _08576_/A2 vssd1 vssd1 vccd1 vccd1 _07796_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12265__A2 _09880_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06746_ reg1_val[12] _07195_/A vssd1 vssd1 vccd1 vccd1 _10927_/S sky130_fd_sc_hd__and2_1
XANTENNA__09666__B1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09534_ _09280_/A _09280_/B _09279_/A vssd1 vssd1 vccd1 vccd1 _09539_/A sky130_fd_sc_hd__a21o_1
X_06677_ reg2_val[23] _06766_/B _06677_/B1 _06676_/Y vssd1 vssd1 vccd1 vccd1 _07036_/A
+ sky130_fd_sc_hd__o2bb2a_4
X_09465_ _09319_/A _09319_/B _09316_/A vssd1 vssd1 vccd1 vccd1 _09471_/A sky130_fd_sc_hd__o21a_1
XANTENNA__07650__A _09667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11172__A _12336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08416_ _08664_/A _08416_/B vssd1 vssd1 vccd1 vccd1 _08452_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13214__B2 _13223_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09396_ _09394_/X _09395_/X _09725_/S vssd1 vssd1 vccd1 vccd1 _09396_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08347_ _08347_/A _08347_/B vssd1 vssd1 vccd1 vccd1 _08355_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07444__A2 _10473_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08278_ _08278_/A _08278_/B vssd1 vssd1 vccd1 vccd1 _08779_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_104_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07229_ _11381_/A _07230_/B vssd1 vssd1 vccd1 vccd1 _07231_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_21_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07097__A _07097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10240_ _10240_/A _10476_/B _10476_/C vssd1 vssd1 vccd1 vccd1 _10242_/C sky130_fd_sc_hd__or3_1
XFILLER_0_42_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10171_ _09425_/C _10303_/B hold260/A vssd1 vssd1 vccd1 vccd1 _10171_/Y sky130_fd_sc_hd__a21oi_1
Xfanout140 _07172_/Y vssd1 vssd1 vccd1 vccd1 _09472_/A sky130_fd_sc_hd__buf_6
Xfanout173 _12816_/B vssd1 vssd1 vccd1 vccd1 _12826_/B sky130_fd_sc_hd__clkbuf_4
Xfanout162 _12322_/A1 vssd1 vssd1 vccd1 vccd1 _11538_/A sky130_fd_sc_hd__clkbuf_4
Xfanout151 _07031_/Y vssd1 vssd1 vccd1 vccd1 _08657_/B sky130_fd_sc_hd__buf_6
XFILLER_0_89_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout195 _09237_/X vssd1 vssd1 vccd1 vccd1 _12205_/B1 sky130_fd_sc_hd__buf_4
Xfanout184 _07314_/B vssd1 vssd1 vccd1 vccd1 _07215_/B sky130_fd_sc_hd__buf_8
XANTENNA__07904__B1 _09940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07380__A1 _10871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07380__B2 _07198_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12812_ hold70/X _12820_/B vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__or2_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12743_ _12743_/A _12743_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[20] sky130_fd_sc_hd__nor2_8
XFILLER_0_96_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13205__B2 _13223_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10019__A1 _10297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12674_ reg1_val[7] _12675_/B vssd1 vssd1 vccd1 vccd1 _12674_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07683__A2 _08484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11625_ _11799_/A _11625_/B vssd1 vssd1 vccd1 vccd1 _11841_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__12413__C1 _12446_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11556_ _10159_/A _11030_/B _11042_/Y _09222_/Y _11555_/X vssd1 vssd1 vccd1 vccd1
+ _11556_/X sky130_fd_sc_hd__o221a_1
XANTENNA__09487__A _10479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10507_ _11779_/A fanout32/X fanout30/X _11764_/A vssd1 vssd1 vccd1 vccd1 _10508_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13226_ hold276/X _13225_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13226_/X sky130_fd_sc_hd__mux2_1
X_11487_ _11487_/A _11487_/B vssd1 vssd1 vccd1 vccd1 _11490_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_110_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10438_ hold281/A _10569_/C vssd1 vssd1 vccd1 vccd1 _10438_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13157_ _13246_/A hold289/X vssd1 vssd1 vccd1 vccd1 _13372_/D sky130_fd_sc_hd__and2_1
X_10369_ _10201_/A _10201_/B _10198_/A vssd1 vssd1 vccd1 vccd1 _10379_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09934__B _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12641__A _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08935__A2 _12823_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12108_ _12108_/A _12108_/B _12108_/C vssd1 vssd1 vccd1 vccd1 _12109_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_85_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13088_ hold72/X _13094_/A2 _13250_/B hold13/X _13039_/A vssd1 vssd1 vccd1 vccd1
+ hold76/A sky130_fd_sc_hd__o221a_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12039_ _12041_/A vssd1 vssd1 vccd1 vccd1 _12039_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08148__B1 _10476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06600_ instruction[12] _06590_/X _06599_/X _06716_/B vssd1 vssd1 vccd1 vccd1 reg1_idx[1]
+ sky130_fd_sc_hd__o211a_4
X_07580_ _07580_/A _07580_/B vssd1 vssd1 vccd1 vccd1 _07581_/B sky130_fd_sc_hd__nor2_1
X_09250_ _11138_/A _09250_/B vssd1 vssd1 vccd1 vccd1 _11247_/C sky130_fd_sc_hd__or2_2
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08201_ _08211_/A _08211_/B vssd1 vssd1 vccd1 vccd1 _08201_/X sky130_fd_sc_hd__and2b_1
XANTENNA__11758__A1 _07051_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09181_ _09179_/X _09180_/X _09403_/S vssd1 vssd1 vccd1 vccd1 _09181_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_50_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11758__B2 _12169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06814__A _12644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08132_ _08215_/A _08215_/B vssd1 vssd1 vccd1 vccd1 _08216_/A sky130_fd_sc_hd__and2_1
XFILLER_0_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08063_ _07974_/A _07974_/C _07974_/B vssd1 vssd1 vccd1 vccd1 _08064_/C sky130_fd_sc_hd__o21ai_1
X_07014_ _07014_/A _07014_/B vssd1 vssd1 vccd1 vccd1 _07014_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__10336__A _12087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08387__B1 _09940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10194__B1 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08965_ _08965_/A _08965_/B vssd1 vssd1 vccd1 vccd1 _08969_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11167__A _12096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07916_ _07913_/A _07913_/B _07913_/C vssd1 vssd1 vccd1 vccd1 _07918_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__10071__A _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09887__B1 _09221_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08896_ _08896_/A _08896_/B vssd1 vssd1 vccd1 vccd1 _08898_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07847_ _08454_/A _07847_/B vssd1 vssd1 vccd1 vccd1 _07850_/A sky130_fd_sc_hd__xnor2_1
X_07778_ _09298_/B2 fanout53/X fanout51/X _09298_/A1 vssd1 vssd1 vccd1 vccd1 _07779_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06729_ reg2_val[15] _06810_/B vssd1 vssd1 vccd1 vccd1 _06729_/X sky130_fd_sc_hd__and2_1
X_09517_ _09518_/A _09518_/B vssd1 vssd1 vccd1 vccd1 _09519_/A sky130_fd_sc_hd__and2_1
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11997__A1 _07036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout26_A _07235_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09448_ _07283_/X _07362_/B fanout16/X _09934_/A vssd1 vssd1 vccd1 vccd1 _09449_/B
+ sky130_fd_sc_hd__o22a_1
X_09379_ _09154_/X _09157_/X _09383_/S vssd1 vssd1 vccd1 vccd1 _09379_/X sky130_fd_sc_hd__mux2_1
X_11410_ _11410_/A _11410_/B _11410_/C vssd1 vssd1 vccd1 vccd1 _11412_/A sky130_fd_sc_hd__and3_1
X_12390_ _12390_/A _12390_/B vssd1 vssd1 vccd1 vccd1 _12391_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_62_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11341_ _11840_/A _11840_/B vssd1 vssd1 vccd1 vccd1 _11567_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_105_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10246__A _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11272_ _11893_/A _12050_/A vssd1 vssd1 vccd1 vccd1 _11272_/X sky130_fd_sc_hd__or2_1
XANTENNA__08378__B1 _09479_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13011_ _13210_/A hold192/X vssd1 vssd1 vccd1 vccd1 _13315_/D sky130_fd_sc_hd__and2_1
XANTENNA__12461__A _12642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10223_ _10224_/A _10224_/B vssd1 vssd1 vccd1 vccd1 _10395_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10185__B1 _11752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10154_ _06828_/X _10153_/Y _12054_/S vssd1 vssd1 vccd1 vccd1 _10155_/B sky130_fd_sc_hd__mux2_1
X_10085_ _10085_/A _10085_/B vssd1 vssd1 vccd1 vccd1 _10086_/B sky130_fd_sc_hd__xnor2_2
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10488__B2 _10595_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10488__A1 _10974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06618__B _06675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10987_ _10879_/A _10879_/B _10878_/A vssd1 vssd1 vccd1 vccd1 _10998_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_85_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08302__B1 _09479_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12726_ _12726_/A _12726_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[16] sky130_fd_sc_hd__xor2_4
XFILLER_0_29_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12657_ _12657_/A _12657_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[3] sky130_fd_sc_hd__xnor2_4
X_11608_ _11609_/B _11609_/A vssd1 vssd1 vccd1 vccd1 _11705_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__13231__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07408__A2 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12588_ _12633_/A _12589_/B vssd1 vssd1 vccd1 vccd1 _12598_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_108_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11539_ _06721_/B _11447_/B _06719_/X vssd1 vssd1 vccd1 vccd1 _11539_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13209_ hold266/X _13209_/A2 _13208_/X _13223_/B2 vssd1 vssd1 vccd1 vccd1 hold267/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06919__A1 _06783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09156__S _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12215__D_N _12214_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08750_ _08751_/B _08751_/C vssd1 vssd1 vccd1 vccd1 _11128_/B sky130_fd_sc_hd__nor2_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11676__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09680__A _11946_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08681_ _08681_/A _08681_/B _08681_/C vssd1 vssd1 vccd1 vccd1 _08737_/A sky130_fd_sc_hd__nand3_1
X_07701_ _07701_/A _07701_/B vssd1 vssd1 vccd1 vccd1 _07784_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07344__A1 _07148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07632_ _09834_/A _07632_/B vssd1 vssd1 vccd1 vccd1 _07634_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07344__B2 _07417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09302_ _09302_/A _09302_/B _09302_/C vssd1 vssd1 vccd1 vccd1 _09306_/B sky130_fd_sc_hd__nand3_1
X_07563_ _07563_/A _07563_/B vssd1 vssd1 vccd1 vccd1 _07565_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_118_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07647__A2 fanout86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07494_ _07566_/A _07566_/B _07493_/A vssd1 vssd1 vccd1 vccd1 _07561_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_29_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09233_ _09234_/C _09233_/B instruction[5] vssd1 vssd1 vccd1 vccd1 _11995_/B sky130_fd_sc_hd__and3b_4
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_15_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13354_/CLK sky130_fd_sc_hd__clkbuf_8
X_09164_ reg1_val[6] reg1_val[25] _09180_/S vssd1 vssd1 vccd1 vccd1 _09164_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08115_ _09341_/A _08159_/B _08159_/A vssd1 vssd1 vccd1 vccd1 _08121_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_16_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09095_ _06993_/A _12158_/B _09672_/A vssd1 vssd1 vccd1 vccd1 _09097_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08046_ _08046_/A _08046_/B vssd1 vssd1 vccd1 vccd1 _08099_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_102_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12156__B2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12156__A1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09997_ _09997_/A _09997_/B vssd1 vssd1 vccd1 vccd1 _09998_/B sky130_fd_sc_hd__xor2_4
X_08948_ _08948_/A _08948_/B vssd1 vssd1 vccd1 vccd1 _09001_/A sky130_fd_sc_hd__xnor2_2
X_08879_ _09936_/A _08879_/B vssd1 vssd1 vccd1 vccd1 _08880_/B sky130_fd_sc_hd__xnor2_2
X_10910_ _06840_/X _10909_/Y _11813_/S vssd1 vssd1 vccd1 vccd1 _10910_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_98_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11890_ _12042_/A _11890_/B vssd1 vssd1 vccd1 vccd1 _12049_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_67_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10841_ _11868_/A fanout47/X fanout45/X fanout62/X vssd1 vssd1 vccd1 vccd1 _10842_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_94_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10772_ _10772_/A _10772_/B vssd1 vssd1 vccd1 vccd1 _10774_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07099__B1 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08835__B2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08835__A1 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12511_ _12511_/A _12511_/B _12511_/C vssd1 vssd1 vccd1 vccd1 _12512_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_82_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12442_ _12364_/A _08924_/X _09040_/D vssd1 vssd1 vccd1 vccd1 _12442_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08599__B1 _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12373_ _12373_/A _12373_/B vssd1 vssd1 vccd1 vccd1 _12380_/A sky130_fd_sc_hd__nor2_1
X_11324_ _11324_/A _11324_/B vssd1 vssd1 vccd1 vccd1 _11326_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_120_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11255_ hold272/A _11255_/B vssd1 vssd1 vccd1 vccd1 _11356_/B sky130_fd_sc_hd__or2_1
X_10206_ fanout56/X fanout86/X fanout82/X _12233_/A vssd1 vssd1 vccd1 vccd1 _10207_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07285__A _09836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11186_ _07051_/X fanout32/X fanout30/X _12169_/A vssd1 vssd1 vccd1 vccd1 _11187_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06782__C1 _12670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10137_ _10137_/A _10137_/B _10331_/A _10542_/A vssd1 vssd1 vccd1 vccd1 _10138_/C
+ sky130_fd_sc_hd__or4_4
X_10068_ _10069_/A _10069_/B vssd1 vssd1 vccd1 vccd1 _10068_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13226__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07326__B2 _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07326__A1 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07629__A2 _07166_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12709_ _12717_/A _12709_/B vssd1 vssd1 vccd1 vccd1 _12711_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_127_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12386__A1 _08859_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold226 hold226/A vssd1 vssd1 vccd1 vccd1 hold226/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 hold204/A vssd1 vssd1 vccd1 vccd1 hold204/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 hold215/A vssd1 vssd1 vccd1 vccd1 hold215/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold259 hold259/A vssd1 vssd1 vccd1 vccd1 hold259/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09920_ _09920_/A _09920_/B vssd1 vssd1 vccd1 vccd1 _09923_/A sky130_fd_sc_hd__nor2_1
Xhold248 hold248/A vssd1 vssd1 vccd1 vccd1 hold248/X sky130_fd_sc_hd__buf_1
Xhold237 hold237/A vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09003__A1 _10871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07195__A _07195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07907__B _07907_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09003__B2 _08112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09851_ _09686_/A _09686_/B _09684_/Y vssd1 vssd1 vccd1 vccd1 _09853_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_0_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06994_ _06987_/A _06987_/B _07094_/B vssd1 vssd1 vccd1 vccd1 _06994_/X sky130_fd_sc_hd__a21o_1
XANTENNA__11361__A2 _12422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09782_ _09782_/A _09782_/B _09782_/C vssd1 vssd1 vccd1 vccd1 _09783_/B sky130_fd_sc_hd__and3_1
X_08802_ _08802_/A _08802_/B vssd1 vssd1 vccd1 vccd1 _12258_/C sky130_fd_sc_hd__xnor2_2
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08733_ _08733_/A _08733_/B _08733_/C vssd1 vssd1 vccd1 vccd1 _10668_/C sky130_fd_sc_hd__nand3_2
XANTENNA__07923__A _08454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout180_A _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12861__A2 _12863_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08664_ _08664_/A _08664_/B _09556_/B vssd1 vssd1 vccd1 vccd1 _08714_/A sky130_fd_sc_hd__or3_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08595_ _08583_/A _08582_/C _08582_/B vssd1 vssd1 vccd1 vccd1 _08596_/C sky130_fd_sc_hd__a21o_1
X_07615_ _07615_/A _07615_/B vssd1 vssd1 vccd1 vccd1 _07628_/A sky130_fd_sc_hd__xor2_2
X_07546_ _07546_/A _07546_/B vssd1 vssd1 vccd1 vccd1 _07708_/A sky130_fd_sc_hd__xor2_2
XANTENNA__10624__A1 _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10624__B2 _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09216_ _09184_/X _09215_/X _11247_/A vssd1 vssd1 vccd1 vccd1 _09216_/X sky130_fd_sc_hd__mux2_2
X_07477_ _09341_/A _07477_/B vssd1 vssd1 vccd1 vccd1 _07534_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09147_ _09147_/A _09863_/A vssd1 vssd1 vccd1 vccd1 _10321_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09793__A2 fanout86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09078_ _09079_/B vssd1 vssd1 vccd1 vccd1 _09078_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08029_ _08065_/B _08027_/B _08027_/C _08024_/Y vssd1 vssd1 vccd1 vccd1 _08056_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout93_A _09779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11339__B _11340_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11040_ _12421_/A1 _11039_/X _06743_/B vssd1 vssd1 vccd1 vccd1 _11040_/X sky130_fd_sc_hd__a21o_1
XANTENNA__08929__A _09834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12991_ _13001_/A hold218/X vssd1 vssd1 vccd1 vccd1 _13305_/D sky130_fd_sc_hd__and2_1
X_11942_ _12087_/A fanout10/X fanout5/X _12009_/A vssd1 vssd1 vccd1 vccd1 _11943_/B
+ sky130_fd_sc_hd__o22a_1
X_11873_ _11873_/A _11873_/B vssd1 vssd1 vccd1 vccd1 _11874_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_39_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10824_ _11538_/A _10824_/B vssd1 vssd1 vccd1 vccd1 _10824_/X sky130_fd_sc_hd__and2_1
XANTENNA__10615__A1 _10748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08664__A _08664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11090__A _12017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10755_ _10755_/A _10755_/B vssd1 vssd1 vccd1 vccd1 _10756_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_82_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09481__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09481__B2 _09943_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10686_ _11990_/A1 _10805_/B hold213/A vssd1 vssd1 vccd1 vccd1 _10686_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10091__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12425_ _12425_/A _12425_/B _12425_/C _12424_/X vssd1 vssd1 vccd1 vccd1 _12425_/X
+ sky130_fd_sc_hd__or4b_1
X_12356_ _12399_/B _12355_/X _12356_/B1 vssd1 vssd1 vccd1 vccd1 _12356_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11040__A1 _12421_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11307_ _12017_/A _11307_/B vssd1 vssd1 vccd1 vccd1 _11308_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07795__A1 _08561_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07795__B2 _08576_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12125__S _12404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12287_ _12287_/A _12287_/B vssd1 vssd1 vccd1 vccd1 _12291_/A sky130_fd_sc_hd__xnor2_1
X_11238_ _06846_/X _11237_/X _11813_/S vssd1 vssd1 vccd1 vccd1 _11239_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07547__A1 _09934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11169_ _11168_/B _11169_/B vssd1 vssd1 vccd1 vccd1 _11170_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__11343__A2 _11567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07547__B2 _08112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13096__A2 _06577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12843__A2 _12863_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07400_ _07400_/A _07400_/B _07435_/A vssd1 vssd1 vccd1 vccd1 _07401_/B sky130_fd_sc_hd__nor3_1
X_08380_ _08384_/A _08384_/B vssd1 vssd1 vccd1 vccd1 _08380_/X sky130_fd_sc_hd__and2_1
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12808__B _12820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07331_ _09661_/B2 _10473_/B2 _10240_/A fanout98/X vssd1 vssd1 vccd1 vccd1 _07332_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12096__A _12096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06806__B _07172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07262_ _07262_/A _07262_/B vssd1 vssd1 vccd1 vccd1 _07262_/X sky130_fd_sc_hd__xor2_4
XANTENNA__10082__A2 _10234_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07193_ _07133_/A _06974_/B _06978_/C _06976_/X _07215_/B vssd1 vssd1 vccd1 vccd1
+ _07195_/B sky130_fd_sc_hd__o41a_4
XFILLER_0_5_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09001_ _09001_/A _09001_/B vssd1 vssd1 vccd1 vccd1 _09016_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_14_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13020__A2 _13171_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11031__A1 _12412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09903_ _09889_/Y _09890_/X _09902_/X vssd1 vssd1 vccd1 vccd1 _09903_/Y sky130_fd_sc_hd__o21ai_1
X_09834_ _09834_/A _09834_/B vssd1 vssd1 vccd1 vccd1 _09838_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06977_ _11038_/A _07195_/A _10813_/A _07233_/A vssd1 vssd1 vccd1 vccd1 _06978_/D
+ sky130_fd_sc_hd__or4_4
XANTENNA__12819__C1 _13147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09765_ _09765_/A _09765_/B _10321_/C _09715_/B vssd1 vssd1 vccd1 vccd1 _09909_/A
+ sky130_fd_sc_hd__nor4b_1
X_08716_ _08575_/A _08666_/A _08660_/X _08714_/A vssd1 vssd1 vccd1 vccd1 _08717_/B
+ sky130_fd_sc_hd__o31ai_1
X_09696_ _09696_/A _09696_/B vssd1 vssd1 vccd1 vccd1 _09697_/B sky130_fd_sc_hd__xnor2_4
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08647_ _12642_/A _07166_/Y _07173_/Y _07983_/A vssd1 vssd1 vccd1 vccd1 _08648_/B
+ sky130_fd_sc_hd__a22o_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08578_ _08608_/A _08608_/B _08578_/C vssd1 vssd1 vccd1 vccd1 _08583_/A sky130_fd_sc_hd__nand3_2
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08484__A _09404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07529_ _07529_/A _07735_/A vssd1 vssd1 vccd1 vccd1 _07559_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10073__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10540_ _10661_/B _10661_/C vssd1 vssd1 vccd1 vccd1 _10780_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11270__A1 _12471_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10471_ _10471_/A _10471_/B vssd1 vssd1 vccd1 vccd1 _10519_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08018__A2 _10595_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12210_ _09221_/Y _10016_/Y _10026_/X _12379_/B2 _12209_/Y vssd1 vssd1 vccd1 vccd1
+ _12211_/D sky130_fd_sc_hd__a221o_1
XFILLER_0_44_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13190_ hold246/X _13189_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13190_/X sky130_fd_sc_hd__mux2_1
XANTENNA__06732__A _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12141_ _12447_/B1 _12203_/B _13322_/Q vssd1 vssd1 vccd1 vccd1 _12141_/Y sky130_fd_sc_hd__a21oi_1
X_12072_ _11554_/A _12071_/X _06659_/B vssd1 vssd1 vccd1 vccd1 _12072_/X sky130_fd_sc_hd__o21a_1
X_11023_ reg1_val[13] curr_PC[13] vssd1 vssd1 vccd1 vccd1 _11025_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11089__B2 _11198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11089__A1 _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12974_ hold293/X _13257_/A2 fanout2/X _13000_/A2 vssd1 vssd1 vccd1 vccd1 _12975_/B
+ sky130_fd_sc_hd__a22o_1
X_11925_ _11874_/A _11874_/B _11873_/A vssd1 vssd1 vccd1 vccd1 _11959_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_86_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09151__B1 _09150_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_0_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11856_ _11857_/A _11857_/B vssd1 vssd1 vccd1 vccd1 _11935_/B sky130_fd_sc_hd__or2_1
XFILLER_0_67_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06626__B _06675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11787_ _11788_/A _11788_/B vssd1 vssd1 vccd1 vccd1 _11878_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_95_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10807_ hold185/A _11990_/A1 _10921_/B _12205_/B1 vssd1 vssd1 vccd1 vccd1 _10807_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_103_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10738_ _10739_/A _10739_/B vssd1 vssd1 vccd1 vccd1 _10740_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11261__A1 _07262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13002__A2 _13171_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11013__A1 _10006_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12408_ _09040_/A _09040_/B _12364_/A vssd1 vssd1 vccd1 vccd1 _12408_/X sky130_fd_sc_hd__a21o_1
X_10669_ _10669_/A _10669_/B vssd1 vssd1 vccd1 vccd1 _10669_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12644__A _12644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13388_ _13390_/CLK _13388_/D vssd1 vssd1 vccd1 vccd1 hold282/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12210__B1 _10026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09757__A2 _09732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07768__A1 _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12339_ _12339_/A _12339_/B vssd1 vssd1 vccd1 vccd1 _12341_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_50_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12761__B2 _07143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07768__B2 _07830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06900_ _06900_/A _06900_/B _06900_/C vssd1 vssd1 vccd1 vccd1 _06901_/D sky130_fd_sc_hd__and3_1
XFILLER_0_37_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07880_ _07880_/A _07880_/B vssd1 vssd1 vccd1 vccd1 _07944_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07473__A _09836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06831_ _07222_/A reg1_val[7] vssd1 vssd1 vccd1 vccd1 _06831_/X sky130_fd_sc_hd__and2b_1
XANTENNA__13069__A2 _12826_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06762_ _07237_/A vssd1 vssd1 vccd1 vccd1 _07238_/A sky130_fd_sc_hd__inv_2
X_09550_ _09146_/A _09146_/B _09371_/A _09371_/B vssd1 vssd1 vccd1 vccd1 _09550_/Y
+ sky130_fd_sc_hd__o22ai_1
X_09481_ fanout56/X _09650_/A fanout17/X _09943_/B2 vssd1 vssd1 vccd1 vccd1 _09482_/B
+ sky130_fd_sc_hd__o22a_1
X_08501_ _08613_/A _10221_/B2 _08501_/B1 _06992_/A vssd1 vssd1 vccd1 vccd1 _08502_/B
+ sky130_fd_sc_hd__o22a_1
X_06693_ instruction[0] instruction[1] instruction[2] instruction[31] pred_val vssd1
+ vssd1 vccd1 vccd1 _12670_/B sky130_fd_sc_hd__o311a_4
XFILLER_0_77_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08432_ _08434_/A _08434_/B vssd1 vssd1 vccd1 vccd1 _08432_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_93_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10339__A _12157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout143_A _09325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08363_ _08326_/Y _08362_/Y _08325_/Y vssd1 vssd1 vccd1 vccd1 _08363_/X sky130_fd_sc_hd__a21o_1
X_07314_ _08973_/B _07314_/B vssd1 vssd1 vccd1 vccd1 _07315_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_46_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07456__B1 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08294_ _08641_/B _08457_/A2 _08501_/B1 _08627_/A2 vssd1 vssd1 vccd1 vccd1 _08295_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_128_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07245_ reg1_val[11] reg1_val[12] _07248_/B _07248_/A vssd1 vssd1 vccd1 vccd1 _07246_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12201__B1 _12376_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07648__A _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07176_ _07166_/Y _07554_/B _07173_/Y _07175_/A vssd1 vssd1 vccd1 vccd1 _07177_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11555__A2 _09257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09817_ _09817_/A _09817_/B vssd1 vssd1 vccd1 vccd1 _09819_/B sky130_fd_sc_hd__xor2_1
XANTENNA__07383__A _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12268__B1 _11648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09748_ _12322_/A1 _09747_/X hold221/A vssd1 vssd1 vccd1 vccd1 _09748_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10240__C _10476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _11710_/A _11710_/B vssd1 vssd1 vccd1 vccd1 _11884_/A sky130_fd_sc_hd__nand2_4
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _09934_/A _08877_/B fanout6/X _09822_/A vssd1 vssd1 vccd1 vccd1 _09680_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12690_ _12699_/A _12690_/B vssd1 vssd1 vccd1 vccd1 _12693_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07830__B _07830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11641_ _11545_/B _11547_/B _11545_/A vssd1 vssd1 vccd1 vccd1 _11642_/B sky130_fd_sc_hd__a21boi_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09103__A _09103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11572_ _11573_/B _11572_/B vssd1 vssd1 vccd1 vccd1 _11689_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_37_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13311_ _13316_/CLK hold195/X vssd1 vssd1 vccd1 vccd1 hold193/A sky130_fd_sc_hd__dfxtp_1
X_10523_ _10397_/A _10396_/B _10394_/X vssd1 vssd1 vccd1 vccd1 _10528_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_37_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13242_ _13246_/A hold259/X vssd1 vssd1 vccd1 vccd1 _13390_/D sky130_fd_sc_hd__and2_1
XFILLER_0_107_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10454_ _10409_/A _10409_/B _10407_/Y vssd1 vssd1 vccd1 vccd1 _10536_/A sky130_fd_sc_hd__a21o_1
X_13173_ _13173_/A _13173_/B vssd1 vssd1 vccd1 vccd1 _13174_/B sky130_fd_sc_hd__nand2_1
X_10385_ _11182_/A _10385_/B vssd1 vssd1 vccd1 vccd1 _10389_/A sky130_fd_sc_hd__xnor2_1
X_12124_ _06672_/B _12053_/Y _12071_/S vssd1 vssd1 vccd1 vccd1 _12124_/X sky130_fd_sc_hd__o21a_1
XANTENNA__09773__A _09922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10712__A _11929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12055_ _06672_/B _12054_/X _11637_/A vssd1 vssd1 vccd1 vccd1 _12055_/Y sky130_fd_sc_hd__a21oi_1
X_11006_ _11006_/A _11006_/B _11006_/C vssd1 vssd1 vccd1 vccd1 _11007_/B sky130_fd_sc_hd__and3_1
XANTENNA__07922__A1 _08457_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07922__B2 _08501_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10809__A1 _12421_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12957_ hold254/X hold77/X vssd1 vssd1 vccd1 vccd1 _12958_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12888_ hold121/X hold246/X vssd1 vssd1 vccd1 vccd1 _12888_/X sky130_fd_sc_hd__and2b_1
X_11908_ _12447_/B1 _11989_/B hold219/A vssd1 vssd1 vccd1 vccd1 _11908_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10285__A2 _10581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07150__A2 _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10159__A _10159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11839_ _11752_/S _11835_/X _11838_/X vssd1 vssd1 vccd1 vccd1 dest_val[21] sky130_fd_sc_hd__o21ai_4
XFILLER_0_28_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13223__A2 _13223_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09427__B2 _11820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08852__A _09667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07030_ _07030_/A _07030_/B vssd1 vssd1 vccd1 vccd1 _07030_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_3_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08981_ _08981_/A _08981_/B vssd1 vssd1 vccd1 vccd1 _08982_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__11718__A _11884_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08299__A _08575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07932_ _07932_/A _07932_/B vssd1 vssd1 vccd1 vccd1 _07956_/B sky130_fd_sc_hd__xor2_2
XANTENNA__09902__A2 _12420_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07863_ _07863_/A _07863_/B vssd1 vssd1 vccd1 vccd1 _07934_/B sky130_fd_sc_hd__xnor2_4
X_09602_ _09602_/A _09602_/B _09600_/X vssd1 vssd1 vccd1 vccd1 _09602_/X sky130_fd_sc_hd__or3b_1
X_06814_ _12644_/A _09725_/S vssd1 vssd1 vccd1 vccd1 _09418_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_3_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07794_ _07800_/B _07800_/A vssd1 vssd1 vccd1 vccd1 _07794_/X sky130_fd_sc_hd__and2b_1
X_09533_ _09362_/A _09362_/B _09360_/Y vssd1 vssd1 vccd1 vccd1 _09540_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12549__A _12708_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout260_A hold191/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06745_ _06927_/A _06723_/A _12708_/B _06744_/X vssd1 vssd1 vccd1 vccd1 _07195_/A
+ sky130_fd_sc_hd__a31o_4
XANTENNA__09666__A1 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09666__B2 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06676_ _06723_/A _12680_/B vssd1 vssd1 vccd1 vccd1 _06676_/Y sky130_fd_sc_hd__nor2_1
X_09464_ _09464_/A _09464_/B vssd1 vssd1 vccd1 vccd1 _09531_/A sky130_fd_sc_hd__and2_2
XFILLER_0_93_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09395_ _09189_/X _09192_/X _09419_/B vssd1 vssd1 vccd1 vccd1 _09395_/X sky130_fd_sc_hd__mux2_1
X_08415_ _06992_/A _10338_/B2 _08457_/A2 _08613_/A vssd1 vssd1 vccd1 vccd1 _08416_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13214__A2 _13223_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08346_ _08367_/A _08367_/B _08345_/A vssd1 vssd1 vccd1 vccd1 _08355_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_117_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08277_ _08229_/X _08276_/Y _08228_/X vssd1 vssd1 vccd1 vccd1 _08277_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_116_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07228_ reg1_val[18] _07228_/B vssd1 vssd1 vccd1 vccd1 _07230_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07159_ _07158_/B _12158_/A _12224_/A vssd1 vssd1 vccd1 vccd1 _07159_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06955__A2 _12359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10170_ hold248/A hold290/A _10170_/C vssd1 vssd1 vccd1 vccd1 _10303_/B sky130_fd_sc_hd__or3_1
XFILLER_0_100_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout130 _07120_/X vssd1 vssd1 vccd1 vccd1 _09934_/A sky130_fd_sc_hd__clkbuf_4
Xfanout174 _12870_/B vssd1 vssd1 vccd1 vccd1 _12862_/B sky130_fd_sc_hd__buf_4
Xfanout163 _12322_/A1 vssd1 vssd1 vccd1 vccd1 _10049_/A sky130_fd_sc_hd__buf_4
Xfanout141 _07165_/Y vssd1 vssd1 vccd1 vccd1 _08576_/A2 sky130_fd_sc_hd__buf_6
Xfanout152 _07031_/Y vssd1 vssd1 vccd1 vccd1 _09298_/B2 sky130_fd_sc_hd__buf_4
Xfanout185 _06921_/Y vssd1 vssd1 vccd1 vccd1 _13101_/A2 sky130_fd_sc_hd__buf_4
Xfanout196 _09234_/X vssd1 vssd1 vccd1 vccd1 _09422_/B sky130_fd_sc_hd__buf_4
XANTENNA__07904__B2 _08289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07904__A1 _08561_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07380__A2 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12811_ _07148_/Y _13101_/B2 hold155/X _13039_/A vssd1 vssd1 vccd1 vccd1 _13266_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _12760_/A _12742_/B _12742_/C vssd1 vssd1 vccd1 vccd1 _12743_/B sky130_fd_sc_hd__and3_2
XFILLER_0_96_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _12672_/A _12671_/A _12671_/B vssd1 vssd1 vccd1 vccd1 _12677_/A sky130_fd_sc_hd__o21ba_2
XANTENNA__13205__A2 _13223_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11624_ _10784_/B _11229_/X _11620_/Y _11622_/X _11623_/X vssd1 vssd1 vccd1 vccd1
+ _11625_/B sky130_fd_sc_hd__a311o_2
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10707__A _10707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11555_ _07087_/A _09257_/S _11554_/Y _06715_/B vssd1 vssd1 vccd1 vccd1 _11555_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10424__C1 _11637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11486_ _11486_/A _11486_/B vssd1 vssd1 vccd1 vccd1 _11487_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_107_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10506_ _11398_/A _10506_/B vssd1 vssd1 vccd1 vccd1 _10510_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_80_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13225_ _13225_/A _13225_/B vssd1 vssd1 vccd1 vccd1 _13225_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10437_ _06770_/B _11829_/B _11554_/A vssd1 vssd1 vccd1 vccd1 _10437_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13156_ hold288/X _13248_/B1 _13155_/X _13248_/A2 vssd1 vssd1 vccd1 vccd1 hold289/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10368_ _10368_/A _10368_/B vssd1 vssd1 vccd1 vccd1 _10381_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__06920__A _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12641__B _12642_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12107_ _12108_/A _12108_/B _12108_/C vssd1 vssd1 vccd1 vccd1 _12177_/B sky130_fd_sc_hd__a21o_1
XANTENNA__06650__A_N _06998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13087_ _07168_/C _13089_/A2 hold73/X vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__o21a_1
X_10299_ _10296_/X _10298_/X _11247_/A vssd1 vssd1 vccd1 vccd1 _10299_/X sky130_fd_sc_hd__mux2_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12038_ _12040_/A _12040_/B _12040_/C vssd1 vssd1 vccd1 vccd1 _12041_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__13141__B2 _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08148__A1 _08561_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08148__B2 _08561_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09345__B1 _07274_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08200_ _10092_/A _08265_/A _08265_/B vssd1 vssd1 vccd1 vccd1 _08211_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_90_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09180_ _11242_/A reg1_val[16] _09180_/S vssd1 vssd1 vccd1 vccd1 _09180_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12816__B _12816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11758__A2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11720__B _11720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08131_ _08131_/A _08131_/B vssd1 vssd1 vccd1 vccd1 _08215_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_126_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07831__B1 _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08062_ _08062_/A _08062_/B vssd1 vssd1 vccd1 vccd1 _08064_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_113_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07013_ _07014_/A _07014_/B vssd1 vssd1 vccd1 vccd1 _07013_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout106_A _08484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08387__A1 _08538_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10194__A1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10194__B2 _11671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09584__B1 _12205_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07926__A _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08387__B2 _08598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11930__A2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08964_ _08965_/A _08965_/B vssd1 vssd1 vccd1 vccd1 _08964_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_11_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07137__S _11929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07915_ _09673_/A _07915_/B vssd1 vssd1 vccd1 vccd1 _07915_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__09887__A1 _11820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08895_ _08896_/A _08896_/B vssd1 vssd1 vccd1 vccd1 _09022_/B sky130_fd_sc_hd__and2b_1
X_07846_ _10338_/B2 _08484_/B _09479_/B1 _08457_/A2 vssd1 vssd1 vccd1 vccd1 _07847_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07898__B1 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07777_ _07777_/A _07777_/B vssd1 vssd1 vccd1 vccd1 _07845_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06728_ _06726_/X _06728_/B vssd1 vssd1 vccd1 vccd1 _11349_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_78_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09516_ _09834_/A _09516_/B vssd1 vssd1 vccd1 vccd1 _09518_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11997__A2 _09257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09447_ _09364_/A _09364_/B _09365_/Y vssd1 vssd1 vccd1 vccd1 _09545_/A sky130_fd_sc_hd__o21ai_4
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06659_ _12071_/S _06659_/B vssd1 vssd1 vccd1 vccd1 _06672_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_93_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09378_ _10049_/A _09765_/A _09765_/B _09150_/X vssd1 vssd1 vccd1 vccd1 _09378_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout19_A _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08329_ _08358_/A _08358_/B vssd1 vssd1 vccd1 vccd1 _08690_/A sky130_fd_sc_hd__or2_1
XANTENNA__10957__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11340_ _11526_/A _11340_/B vssd1 vssd1 vccd1 vccd1 _11840_/B sky130_fd_sc_hd__and2_1
XFILLER_0_62_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13010_ hold177/X _13171_/B2 _13209_/A2 hold180/X vssd1 vssd1 vccd1 vccd1 hold192/A
+ sky130_fd_sc_hd__a22o_1
X_11271_ _11271_/A _11271_/B _11271_/C _11124_/Y vssd1 vssd1 vccd1 vccd1 _12050_/A
+ sky130_fd_sc_hd__nor4b_4
XANTENNA__08378__A1 _08576_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10222_ _11497_/A _10222_/B vssd1 vssd1 vccd1 vccd1 _10224_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08378__B2 _07172_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07836__A _09947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11382__B1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10153_ _06790_/A _10012_/B _06788_/Y vssd1 vssd1 vccd1 vccd1 _10153_/Y sky130_fd_sc_hd__o21ai_1
X_10084_ _10085_/A _10085_/B vssd1 vssd1 vccd1 vccd1 _10084_/Y sky130_fd_sc_hd__nand2_1
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10488__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11093__A _11093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10986_ _10986_/A _10986_/B vssd1 vssd1 vccd1 vccd1 _11000_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_97_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08302__A1 _08561_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08302__B2 _08576_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12085__A_N _12084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12725_ _12726_/A _12726_/B vssd1 vssd1 vccd1 vccd1 _12739_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_84_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12656_ _12654_/Y _12656_/B vssd1 vssd1 vccd1 vccd1 _12657_/B sky130_fd_sc_hd__and2b_1
X_11607_ _11705_/A _11607_/B vssd1 vssd1 vccd1 vccd1 _11609_/B sky130_fd_sc_hd__nand2_1
X_12587_ reg1_val[19] curr_PC[19] _12638_/S vssd1 vssd1 vccd1 vccd1 _12589_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_53_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06634__B _12719_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10948__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09010__B _11946_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap116 _07199_/X vssd1 vssd1 vccd1 vccd1 _10725_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11538_ _11538_/A _11538_/B _11538_/C vssd1 vssd1 vccd1 vccd1 _11538_/X sky130_fd_sc_hd__and3_1
XFILLER_0_123_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11469_ _11637_/A _11449_/X _11456_/X _11468_/X vssd1 vssd1 vccd1 vccd1 _11469_/X
+ sky130_fd_sc_hd__o211a_1
X_13208_ hold268/A _13207_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13208_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13139_ _13139_/A _13139_/B vssd1 vssd1 vccd1 vccd1 _13139_/Y sky130_fd_sc_hd__xnor2_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11125__B1 _09150_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07700_ _08575_/A _07700_/B vssd1 vssd1 vccd1 vccd1 _07784_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11676__A1 _12009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11676__B2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10900__A _10900_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08577__A _09302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08680_ _08681_/B _08739_/B vssd1 vssd1 vccd1 vccd1 _08733_/B sky130_fd_sc_hd__and2_1
XANTENNA__07481__A _07604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07631_ _07830_/B _07221_/X _09940_/B2 fanout46/X vssd1 vssd1 vccd1 vccd1 _07632_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07344__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07562_ _07562_/A _07562_/B vssd1 vssd1 vccd1 vccd1 _07565_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09301_ _09301_/A _10476_/B _10476_/C vssd1 vssd1 vccd1 vccd1 _09302_/C sky130_fd_sc_hd__or3_1
XFILLER_0_118_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07493_ _07493_/A _07493_/B vssd1 vssd1 vccd1 vccd1 _07566_/B sky130_fd_sc_hd__nor2_1
X_09232_ _09232_/A _09239_/B vssd1 vssd1 vccd1 vccd1 _10788_/A sky130_fd_sc_hd__or2_4
XFILLER_0_29_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09163_ _09161_/X _09162_/X _09383_/S vssd1 vssd1 vccd1 vccd1 _09163_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout223_A _07165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08114_ _10092_/A _08114_/B vssd1 vssd1 vccd1 vccd1 _08159_/B sky130_fd_sc_hd__xnor2_1
X_09094_ _09302_/A _09094_/B vssd1 vssd1 vccd1 vccd1 _09097_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08045_ _08575_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08099_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07280__B2 _07232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12156__A2 _12335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11178__A _11179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09996_ _09997_/A _09997_/B vssd1 vssd1 vccd1 vccd1 _09996_/X sky130_fd_sc_hd__and2_1
X_08947_ _08948_/A _08948_/B vssd1 vssd1 vccd1 vccd1 _09060_/B sky130_fd_sc_hd__nand2b_1
X_08878_ _07172_/Y _07362_/B fanout16/X _09325_/A vssd1 vssd1 vccd1 vccd1 _08879_/B
+ sky130_fd_sc_hd__o22a_1
X_07829_ _07935_/A _07827_/Y _07825_/Y vssd1 vssd1 vccd1 vccd1 _07863_/A sky130_fd_sc_hd__o21a_2
X_10840_ _12096_/A _10840_/B vssd1 vssd1 vccd1 vccd1 _10844_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_79_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10771_ _10772_/A _10772_/B vssd1 vssd1 vccd1 vccd1 _10897_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07099__B2 _10245_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07099__A1 _09661_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08835__A2 _10473_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_5_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12510_ _12511_/A _12511_/B _12511_/C vssd1 vssd1 vccd1 vccd1 _12518_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_81_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12441_ _06962_/B _12439_/X _12440_/Y vssd1 vssd1 vccd1 vccd1 _12441_/X sky130_fd_sc_hd__o21a_1
XANTENNA__08048__B1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08599__B2 _08641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08599__A1 _08627_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12372_ hold241/A _12447_/B1 _12417_/B _11648_/A vssd1 vssd1 vccd1 vccd1 _12373_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_34_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08950__A _10749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11323_ _11324_/B _11324_/A vssd1 vssd1 vccd1 vccd1 _11323_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_120_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12472__A _12650_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11254_ _11648_/A _11254_/B _11254_/C vssd1 vssd1 vccd1 vccd1 _11254_/X sky130_fd_sc_hd__or3_1
XANTENNA__09257__S _09257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10205_ _10116_/A _10116_/B _10113_/A vssd1 vssd1 vccd1 vccd1 _10220_/A sky130_fd_sc_hd__a21oi_1
X_11185_ _12093_/A _11185_/B vssd1 vssd1 vccd1 vccd1 _11189_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_100_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10136_ _10136_/A _10136_/B vssd1 vssd1 vccd1 vccd1 _10661_/A sky130_fd_sc_hd__xnor2_4
X_10067_ _09976_/A _09976_/B _09972_/X vssd1 vssd1 vccd1 vccd1 _10069_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11658__B2 _10788_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07326__A2 _09943_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10969_ _11198_/A fanout10/X fanout5/X _11093_/A vssd1 vssd1 vccd1 vccd1 _10970_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08287__B1 _10476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12708_ reg1_val[13] _12708_/B vssd1 vssd1 vccd1 vccd1 _12709_/B sky130_fd_sc_hd__or2_1
XFILLER_0_73_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10581__D_N _10453_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08039__B1 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12639_ _12639_/A _12639_/B vssd1 vssd1 vccd1 vccd1 _12640_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold205 hold205/A vssd1 vssd1 vccd1 vccd1 hold205/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold216 hold216/A vssd1 vssd1 vccd1 vccd1 hold216/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 hold227/A vssd1 vssd1 vccd1 vccd1 hold227/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 hold249/A vssd1 vssd1 vccd1 vccd1 hold249/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 hold238/A vssd1 vssd1 vccd1 vccd1 hold238/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07907__C _07907_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09003__A2 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09850_ _09850_/A _09850_/B vssd1 vssd1 vccd1 vccd1 _09853_/A sky130_fd_sc_hd__nand2_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _09782_/A _09782_/B _09782_/C vssd1 vssd1 vccd1 vccd1 _09783_/A sky130_fd_sc_hd__a21oi_1
X_06993_ _06993_/A _12644_/A vssd1 vssd1 vccd1 vccd1 _06993_/Y sky130_fd_sc_hd__nand2_8
X_08801_ _08800_/A _08800_/B _08712_/Y _08795_/A _08795_/B vssd1 vssd1 vccd1 vccd1
+ _12258_/B sky130_fd_sc_hd__a2111oi_2
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ _08727_/A _08727_/B _08588_/X _08607_/X vssd1 vssd1 vccd1 vccd1 _08733_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08663_ _08663_/A _09432_/A vssd1 vssd1 vccd1 vccd1 _09556_/B sky130_fd_sc_hd__or2_1
XANTENNA_fanout173_A _12816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07614_ _07614_/A _07614_/B vssd1 vssd1 vccd1 vccd1 _07615_/B sky130_fd_sc_hd__xnor2_2
X_08594_ _08594_/A _08594_/B vssd1 vssd1 vccd1 vccd1 _08596_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_119_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12557__A _12714_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12074__A1 _12379_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07545_ _07546_/A _07546_/B vssd1 vssd1 vccd1 vccd1 _07556_/B sky130_fd_sc_hd__and2_1
XANTENNA__11821__A1 _11820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10624__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07476_ _07221_/X _08112_/B fanout25/X _07283_/X vssd1 vssd1 vccd1 vccd1 _07477_/B
+ sky130_fd_sc_hd__o22a_1
X_09215_ _09199_/X _09214_/X _11138_/A vssd1 vssd1 vccd1 vccd1 _09215_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_64_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12377__A2 _12420_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09778__B1 _07238_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09146_ _09146_/A _09146_/B vssd1 vssd1 vccd1 vccd1 _09863_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_17_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09077_ _10479_/A _09077_/B vssd1 vssd1 vccd1 vccd1 _09079_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08028_ _08024_/Y _08083_/A vssd1 vssd1 vccd1 vccd1 _08028_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout86_A _08411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08202__B1 _09479_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09950__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ _09979_/A _09979_/B vssd1 vssd1 vccd1 vccd1 _09980_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_99_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12990_ hold215/X _13000_/A2 _13257_/A2 hold217/X vssd1 vssd1 vccd1 vccd1 hold218/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09106__A _11946_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11941_ _11851_/A _11851_/B _11861_/A vssd1 vssd1 vccd1 vccd1 _11955_/A sky130_fd_sc_hd__o21a_1
X_11872_ _11872_/A _11872_/B _11872_/C vssd1 vssd1 vccd1 vccd1 _11873_/B sky130_fd_sc_hd__nor3_1
XANTENNA__13262__B1 _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10823_ _11271_/A _11050_/A _11050_/B vssd1 vssd1 vccd1 vccd1 _10824_/B sky130_fd_sc_hd__or3_1
XFILLER_0_39_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10754_ _10755_/A _10755_/B vssd1 vssd1 vccd1 vccd1 _10754_/X sky130_fd_sc_hd__and2_1
XFILLER_0_94_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09481__A2 _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13014__B1 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10685_ hold208/A _10685_/B vssd1 vssd1 vccd1 vccd1 _10805_/B sky130_fd_sc_hd__or2_1
X_12424_ _12418_/Y _12419_/X _12423_/X _12416_/X vssd1 vssd1 vccd1 vccd1 _12424_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12355_ _12050_/X _12399_/A _12306_/X _11892_/A vssd1 vssd1 vccd1 vccd1 _12355_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11306_ _11476_/A fanout10/X fanout5/X _11406_/A vssd1 vssd1 vccd1 vccd1 _11307_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07296__A _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07795__A2 _08112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12286_ _12286_/A _12335_/B vssd1 vssd1 vccd1 vccd1 _12287_/B sky130_fd_sc_hd__nor2_1
X_11237_ _11131_/A _11129_/Y _11150_/S vssd1 vssd1 vccd1 vccd1 _11237_/X sky130_fd_sc_hd__a21o_1
X_11168_ _11169_/B _11168_/B vssd1 vssd1 vccd1 vccd1 _11318_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__10000__B1 _09862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07547__A2 fanout25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10119_ _10120_/A _10120_/B vssd1 vssd1 vccd1 vccd1 _10119_/Y sky130_fd_sc_hd__nand2b_1
X_11099_ _11097_/Y _11099_/B vssd1 vssd1 vccd1 vccd1 _11100_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_117_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07330_ _07387_/A _07387_/B vssd1 vssd1 vccd1 vccd1 _07388_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_18_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07261_ _07262_/A _07262_/B vssd1 vssd1 vccd1 vccd1 _07261_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_5_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09000_ _09000_/A _09000_/B vssd1 vssd1 vccd1 vccd1 _09001_/B sky130_fd_sc_hd__xor2_2
X_07192_ _07189_/Y _07192_/B vssd1 vssd1 vccd1 vccd1 _07192_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_0_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07235__A1 _11582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12824__B _12826_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10625__A _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13001__A _13001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09902_ _06898_/C _12420_/A0 _09901_/X vssd1 vssd1 vccd1 vccd1 _09902_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_6_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09833_ _07830_/B _11093_/A fanout72/X fanout46/X vssd1 vssd1 vccd1 vccd1 _09834_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10360__A _12224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06761__A3 _12689_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06976_ _10813_/A _07233_/A vssd1 vssd1 vccd1 vccd1 _06976_/X sky130_fd_sc_hd__or2_1
X_09764_ _10821_/A _09760_/X _09761_/X _09763_/Y vssd1 vssd1 vccd1 vccd1 dest_val[3]
+ sky130_fd_sc_hd__a22o_4
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08715_ _09556_/B _08715_/B vssd1 vssd1 vccd1 vccd1 _09717_/B sky130_fd_sc_hd__nor2_1
X_09695_ _09694_/A _09694_/B _09696_/A vssd1 vssd1 vccd1 vccd1 _09695_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08646_ _08646_/A _08646_/B _08646_/C vssd1 vssd1 vccd1 vccd1 _08671_/B sky130_fd_sc_hd__and3_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12047__A1 _11340_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08577_ _09302_/A _08577_/B vssd1 vssd1 vccd1 vccd1 _08578_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__08484__B _08484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07528_ _07734_/B _07734_/C _07734_/A vssd1 vssd1 vccd1 vccd1 _07735_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_91_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07459_ _09943_/B2 fanout51/X _09661_/B2 _09650_/A vssd1 vssd1 vccd1 vccd1 _07460_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10470_ _10471_/B _10471_/A vssd1 vssd1 vccd1 vccd1 _10645_/B sky130_fd_sc_hd__and2b_1
XANTENNA__09596__A _12064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09129_ _09127_/Y _09129_/B vssd1 vssd1 vccd1 vccd1 _09130_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_121_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12140_ hold206/A _12140_/B vssd1 vssd1 vccd1 vccd1 _12203_/B sky130_fd_sc_hd__or2_1
XANTENNA__08974__A1 _12359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06732__B _07262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10230__B1 _07269_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11130__S _11813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10781__A1 _10539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12071_ _11995_/B _11829_/B _12071_/S vssd1 vssd1 vccd1 vccd1 _12071_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11022_ _11022_/A _11022_/B vssd1 vssd1 vccd1 vccd1 _11022_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_99_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11089__A2 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12973_ _12973_/A _13247_/B vssd1 vssd1 vccd1 vccd1 fanout2/A sky130_fd_sc_hd__or2_2
X_11924_ _12050_/A _12050_/B _12049_/A _11892_/A vssd1 vssd1 vccd1 vccd1 _11973_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09151__A1 _10049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11855_ _07136_/Y _12158_/B _11854_/X _11929_/A vssd1 vssd1 vccd1 vccd1 _11857_/B
+ sky130_fd_sc_hd__a22o_1
X_11786_ _11878_/A _11786_/B vssd1 vssd1 vccd1 vccd1 _11788_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_103_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10806_ _11990_/A1 _10921_/B hold185/A vssd1 vssd1 vccd1 vccd1 _10806_/Y sky130_fd_sc_hd__a21oi_1
X_10737_ _10737_/A _10737_/B vssd1 vssd1 vccd1 vccd1 _10739_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_94_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11261__A2 _12422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08662__B1 _07148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12407_ _12406_/A _12404_/X _12405_/Y vssd1 vssd1 vccd1 vccd1 _12425_/A sky130_fd_sc_hd__o21a_1
X_10668_ _11809_/A _10668_/B _10668_/C _10668_/D vssd1 vssd1 vccd1 vccd1 _10669_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12644__B _12645_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13387_ _13390_/CLK _13387_/D vssd1 vssd1 vccd1 vccd1 hold284/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12210__A1 _09221_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11013__A2 _10542_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12210__B2 _12379_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10599_ _10599_/A _12087_/B _10600_/A vssd1 vssd1 vccd1 vccd1 _10599_/X sky130_fd_sc_hd__or3_1
XANTENNA__10221__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07768__A2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12338_ _12338_/A _12338_/B vssd1 vssd1 vccd1 vccd1 _12339_/B sky130_fd_sc_hd__and2_1
XFILLER_0_11_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12269_ _12269_/A _12269_/B vssd1 vssd1 vccd1 vccd1 _12277_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09914__B1 _07232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11721__B1 _12356_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06830_ _10155_/A _06828_/X _06829_/Y vssd1 vssd1 vccd1 vccd1 _06830_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06761_ _06815_/A _06817_/B1 _12689_/B _06760_/X vssd1 vssd1 vccd1 vccd1 _07237_/A
+ sky130_fd_sc_hd__a31o_4
X_06692_ reg1_val[20] _07016_/A vssd1 vssd1 vccd1 vccd1 _11726_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09480_ _10749_/A _09480_/B vssd1 vssd1 vccd1 vccd1 _09484_/A sky130_fd_sc_hd__xnor2_1
X_08500_ _08500_/A _08500_/B vssd1 vssd1 vccd1 vccd1 _08522_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08431_ _08431_/A _08431_/B vssd1 vssd1 vccd1 vccd1 _08434_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08362_ _08691_/A vssd1 vssd1 vccd1 vccd1 _08362_/Y sky130_fd_sc_hd__inv_2
X_07313_ _07314_/B _08973_/D _08973_/B vssd1 vssd1 vccd1 vccd1 _10476_/B sky130_fd_sc_hd__a21oi_4
X_08293_ _08664_/A _08293_/B vssd1 vssd1 vccd1 vccd1 _08297_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__07456__B2 _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07456__A1 _09669_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07244_ _07244_/A _07244_/B vssd1 vssd1 vccd1 vccd1 _07370_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_116_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07175_ _07175_/A vssd1 vssd1 vccd1 vccd1 _07175_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_14_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09905__B1 _06958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09816_ _09817_/B _09817_/A vssd1 vssd1 vccd1 vccd1 _09816_/X sky130_fd_sc_hd__and2b_1
X_06959_ _09233_/B instruction[5] vssd1 vssd1 vccd1 vccd1 _09228_/B sky130_fd_sc_hd__nand2_2
X_09747_ hold237/A hold301/A hold293/A vssd1 vssd1 vccd1 vccd1 _09747_/X sky130_fd_sc_hd__or3_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10279__B1 _10136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout49_A _11770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09678_ _09505_/A _09505_/B _09501_/Y vssd1 vssd1 vccd1 vccd1 _09682_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__06727__B _06727_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _08630_/A _08630_/B _08628_/Y vssd1 vssd1 vccd1 vccd1 _08637_/A sky130_fd_sc_hd__nor3b_1
X_11640_ _11640_/A _11640_/B vssd1 vssd1 vccd1 vccd1 _11642_/A sky130_fd_sc_hd__nand2_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09103__B _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11571_ _12093_/A _11571_/B vssd1 vssd1 vccd1 vccd1 _11572_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_119_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13310_ _13316_/CLK hold171/X vssd1 vssd1 vccd1 vccd1 _13310_/Q sky130_fd_sc_hd__dfxtp_1
X_10522_ _10382_/B _10398_/B _10380_/Y vssd1 vssd1 vccd1 vccd1 _10532_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13241_ hold258/X _13248_/B1 _13240_/X _13248_/A2 vssd1 vssd1 vccd1 vccd1 hold259/A
+ sky130_fd_sc_hd__a22o_1
X_10453_ _10453_/A _10453_/B vssd1 vssd1 vccd1 vccd1 _10549_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13172_ _13249_/A hold273/X vssd1 vssd1 vccd1 vccd1 _13375_/D sky130_fd_sc_hd__and2_1
X_10384_ fanout59/X fanout36/X fanout34/X fanout57/X vssd1 vssd1 vccd1 vccd1 _10385_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_58_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12123_ _12184_/B _12123_/B vssd1 vssd1 vccd1 vccd1 _12123_/X sky130_fd_sc_hd__or2_1
X_12054_ _06864_/Y _12053_/Y _12054_/S vssd1 vssd1 vccd1 vccd1 _12054_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12480__A _12655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11005_ _11006_/A _11006_/B _11006_/C vssd1 vssd1 vccd1 vccd1 _11007_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07922__A2 _08484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12956_ _13211_/A _13212_/A _13211_/B vssd1 vssd1 vccd1 vccd1 _13216_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_59_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12887_ hold264/X hold96/X vssd1 vssd1 vccd1 vccd1 _13193_/A sky130_fd_sc_hd__nand2b_1
X_11907_ hold188/A _11907_/B vssd1 vssd1 vccd1 vccd1 _11989_/B sky130_fd_sc_hd__or2_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ _12471_/S _11838_/B _12003_/C vssd1 vssd1 vccd1 vccd1 _11838_/X sky130_fd_sc_hd__or3_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10159__B _10159_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11769_ _12093_/A _11769_/B vssd1 vssd1 vccd1 vccd1 _11770_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07989__A2 _07097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12982__A2 _13000_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11942__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07205__A4 _07109_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08980_ _08981_/A _08981_/B vssd1 vssd1 vccd1 vccd1 _08980_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07931_ _07968_/A _07968_/B _07929_/B _07930_/Y vssd1 vssd1 vccd1 vccd1 _07956_/A
+ sky130_fd_sc_hd__o31ai_4
X_07862_ _07937_/A _07937_/B _07855_/X vssd1 vssd1 vccd1 vccd1 _07934_/A sky130_fd_sc_hd__a21o_2
X_09601_ _07172_/A _12422_/A _12356_/B1 _09555_/Y vssd1 vssd1 vccd1 vccd1 _09602_/A
+ sky130_fd_sc_hd__a22o_1
X_06813_ _12644_/A _07149_/A vssd1 vssd1 vccd1 vccd1 _09586_/A sky130_fd_sc_hd__or2_1
XFILLER_0_3_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07793_ _07826_/A _07826_/B _07789_/Y vssd1 vssd1 vccd1 vccd1 _07800_/B sky130_fd_sc_hd__o21ba_1
X_09532_ _09352_/A _09352_/B _09355_/A vssd1 vssd1 vccd1 vccd1 _09542_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_78_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06744_ reg2_val[12] _06810_/B vssd1 vssd1 vccd1 vccd1 _06744_/X sky130_fd_sc_hd__and2_1
X_06675_ instruction[33] _06675_/B vssd1 vssd1 vccd1 vccd1 _12680_/B sky130_fd_sc_hd__and2_4
X_09463_ _09463_/A _09463_/B _09463_/C vssd1 vssd1 vccd1 vccd1 _09464_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_93_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09394_ _09186_/X _09188_/X _09403_/S vssd1 vssd1 vccd1 vccd1 _09394_/X sky130_fd_sc_hd__mux2_1
X_08414_ _08427_/A _08427_/B vssd1 vssd1 vccd1 vccd1 _08414_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_86_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08345_ _08345_/A _08345_/B vssd1 vssd1 vccd1 vccd1 _08367_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_19_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13160__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08276_ _08280_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08276_/Y sky130_fd_sc_hd__nand2_1
X_07227_ _07227_/A _07227_/B vssd1 vssd1 vccd1 vccd1 _07241_/A sky130_fd_sc_hd__nor2_2
XANTENNA__12186__B1 _09150_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07158_ _12224_/A _07158_/B vssd1 vssd1 vccd1 vccd1 _07158_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_14_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09051__B1 _12823_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07089_ reg1_val[8] _07089_/B vssd1 vssd1 vccd1 vccd1 _07091_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_100_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout120 _07194_/Y vssd1 vssd1 vccd1 vccd1 _10871_/A sky130_fd_sc_hd__buf_4
Xfanout131 _07098_/X vssd1 vssd1 vccd1 vccd1 _08515_/A2 sky130_fd_sc_hd__buf_6
Xfanout164 _11990_/A1 vssd1 vssd1 vccd1 vccd1 _11646_/B sky130_fd_sc_hd__buf_4
Xfanout142 _07165_/Y vssd1 vssd1 vccd1 vccd1 _09677_/A sky130_fd_sc_hd__buf_4
Xfanout153 _07015_/X vssd1 vssd1 vccd1 vccd1 _08627_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout175 _12816_/B vssd1 vssd1 vccd1 vccd1 _12870_/B sky130_fd_sc_hd__buf_2
Xfanout197 _09228_/X vssd1 vssd1 vccd1 vccd1 _12420_/A0 sky130_fd_sc_hd__buf_4
Xfanout186 _06921_/Y vssd1 vssd1 vccd1 vccd1 _13250_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__07904__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12810_ hold154/X _12820_/B vssd1 vssd1 vccd1 vccd1 hold155/A sky130_fd_sc_hd__or2_1
XFILLER_0_97_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ _12742_/B _12742_/C _12760_/A vssd1 vssd1 vccd1 vccd1 _12743_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_96_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ _12672_/A _12672_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[6] sky130_fd_sc_hd__xor2_4
X_11623_ _11623_/A _11623_/B _11800_/A vssd1 vssd1 vccd1 vccd1 _11623_/X sky130_fd_sc_hd__and3_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12413__A1 _12412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11554_ _11554_/A _11554_/B vssd1 vssd1 vccd1 vccd1 _11554_/Y sky130_fd_sc_hd__nor2_1
X_11485_ _11486_/A _11486_/B vssd1 vssd1 vccd1 vccd1 _11487_/A sky130_fd_sc_hd__and2_1
X_10505_ _07097_/X _07171_/A _07175_/A _07256_/Y vssd1 vssd1 vccd1 vccd1 _10506_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13224_ _13249_/A hold277/X vssd1 vssd1 vccd1 vccd1 _13386_/D sky130_fd_sc_hd__and2_1
XFILLER_0_100_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10436_ hold217/A _11990_/A1 _10565_/B _12205_/B1 vssd1 vssd1 vccd1 vccd1 _10436_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_110_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11924__B1 _11892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13155_ hold279/X _13154_/Y fanout2/A vssd1 vssd1 vccd1 vccd1 _13155_/X sky130_fd_sc_hd__mux2_1
X_10367_ _10367_/A _10367_/B vssd1 vssd1 vccd1 vccd1 _10368_/B sky130_fd_sc_hd__xor2_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12106_ _12177_/A _12106_/B vssd1 vssd1 vccd1 vccd1 _12108_/C sky130_fd_sc_hd__nand2_1
X_10298_ _11247_/B _10297_/X _11138_/A vssd1 vssd1 vccd1 vccd1 _10298_/X sky130_fd_sc_hd__mux2_1
X_13086_ hold108/A _13094_/A2 _13250_/B hold72/X _13259_/A vssd1 vssd1 vccd1 vccd1
+ hold73/A sky130_fd_sc_hd__o221a_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12037_ _12111_/B _12037_/B vssd1 vssd1 vccd1 vccd1 _12040_/C sky130_fd_sc_hd__nand2_1
XANTENNA__13141__A2 _13254_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09345__A1 _10234_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08148__A2 _08411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09345__B2 _07959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11152__A1 _07270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11554__A _11554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06648__A _06723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12939_ _13173_/A _13174_/A _13173_/B vssd1 vssd1 vccd1 vccd1 _13179_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_88_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08856__B1 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12385__A fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08130_ _08198_/A _08198_/B vssd1 vssd1 vccd1 vccd1 _08215_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_126_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07831__A1 _07020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08061_ _07965_/B _08061_/B vssd1 vssd1 vccd1 vccd1 _08062_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_114_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07012_ _06987_/A _06986_/C _07094_/B vssd1 vssd1 vccd1 vccd1 _07014_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_3_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12832__B _12862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08387__A2 _08561_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07595__B1 _11844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10194__A2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08963_ _10092_/A _08963_/B vssd1 vssd1 vccd1 vccd1 _08965_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07914_ _07030_/Y _07983_/B _07097_/X _07038_/X vssd1 vssd1 vccd1 vccd1 _07915_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09887__A2 _12446_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08894_ _09022_/A _08894_/B vssd1 vssd1 vccd1 vccd1 _08896_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_75_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07845_ _07845_/A _07845_/B vssd1 vssd1 vccd1 vccd1 _07861_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07898__A1 _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07898__B2 _07172_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07776_ _07777_/A _07777_/B vssd1 vssd1 vccd1 vccd1 _07776_/Y sky130_fd_sc_hd__nand2_1
X_06727_ reg1_val[16] _06727_/B vssd1 vssd1 vccd1 vccd1 _06728_/B sky130_fd_sc_hd__or2_1
XFILLER_0_79_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09515_ _07830_/B _10595_/A1 _10338_/B2 fanout46/X vssd1 vssd1 vccd1 vccd1 _09516_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08847__B1 _10974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09446_ _09369_/A _09369_/B _09367_/X vssd1 vssd1 vccd1 vccd1 _09548_/A sky130_fd_sc_hd__a21oi_4
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06658_ reg1_val[24] _06658_/B vssd1 vssd1 vccd1 vccd1 _06659_/B sky130_fd_sc_hd__or2_1
XFILLER_0_38_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06589_ instruction[1] instruction[2] instruction[0] pred_val vssd1 vssd1 vccd1 vccd1
+ _06944_/B sky130_fd_sc_hd__and4b_4
X_09377_ _10049_/A _09765_/A _09765_/B vssd1 vssd1 vccd1 vccd1 _09377_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10957__A1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08328_ _08328_/A _08328_/B vssd1 vssd1 vccd1 vccd1 _08358_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_19_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09272__B1 _07282_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10957__B2 _11868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08259_ _08255_/A _08255_/B _08258_/Y vssd1 vssd1 vccd1 vccd1 _08286_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_104_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11270_ _12471_/S _11266_/X _11267_/X _11269_/Y vssd1 vssd1 vccd1 vccd1 dest_val[15]
+ sky130_fd_sc_hd__a22o_4
XANTENNA__08378__A2 _10473_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11382__A1 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10221_ _10500_/A _08877_/B fanout6/X _10221_/B2 vssd1 vssd1 vccd1 vccd1 _10222_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11382__B2 _07231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10152_ _10788_/A _10152_/B _10151_/X vssd1 vssd1 vccd1 vccd1 _10152_/X sky130_fd_sc_hd__or3b_1
X_10083_ _12224_/A _10083_/B vssd1 vssd1 vccd1 vccd1 _10085_/B sky130_fd_sc_hd__xor2_2
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07852__A _10246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11093__B _12087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10985_ _10984_/A _10984_/B _10984_/C vssd1 vssd1 vccd1 vccd1 _10986_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09779__A _09779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12724_ reg1_val[15] _12719_/B _12722_/A vssd1 vssd1 vccd1 vccd1 _12726_/B sky130_fd_sc_hd__a21o_2
XANTENNA__08302__A2 _08484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07510__B1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12655_ reg1_val[3] _12655_/B vssd1 vssd1 vccd1 vccd1 _12656_/B sky130_fd_sc_hd__nand2_1
X_11606_ _11606_/A _11606_/B vssd1 vssd1 vccd1 vccd1 _11607_/B sky130_fd_sc_hd__nand2_1
X_12586_ _12591_/B _12586_/B vssd1 vssd1 vccd1 vccd1 new_PC[18] sky130_fd_sc_hd__and2_4
XFILLER_0_108_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06616__A2 _12796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10948__A1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10948__B2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11537_ _11538_/A _11538_/B _11538_/C vssd1 vssd1 vccd1 vccd1 _11537_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11468_ _10159_/A _11141_/B _11460_/Y _11467_/X vssd1 vssd1 vccd1 vccd1 _11468_/X
+ sky130_fd_sc_hd__o211a_1
Xmax_cap139 _07221_/B vssd1 vssd1 vccd1 vccd1 _07222_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13207_ _13207_/A _13207_/B vssd1 vssd1 vccd1 vccd1 _13207_/Y sky130_fd_sc_hd__xnor2_1
X_11399_ _11399_/A _11399_/B vssd1 vssd1 vccd1 vccd1 _11401_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11373__A1 _12471_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10419_ _11630_/A _10420_/B _10420_/C vssd1 vssd1 vccd1 vccd1 _10419_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_0_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07577__B1 _07238_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13138_ _13138_/A _13138_/B vssd1 vssd1 vccd1 vccd1 _13139_/B sky130_fd_sc_hd__nand2_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _09667_/A _12826_/B hold136/X vssd1 vssd1 vccd1 vccd1 _13344_/D sky130_fd_sc_hd__a21boi_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11676__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10900__B _11008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11284__A _11284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07630_ _09779_/A _07630_/B vssd1 vssd1 vccd1 vccd1 _07634_/A sky130_fd_sc_hd__xor2_1
X_07561_ _07561_/A _07561_/B vssd1 vssd1 vccd1 vccd1 _07568_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_88_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09300_ _07608_/A _07608_/B _09669_/B2 vssd1 vssd1 vccd1 vccd1 _09302_/B sky130_fd_sc_hd__a21o_1
X_07492_ _07492_/A _07492_/B _07535_/A vssd1 vssd1 vccd1 vccd1 _07493_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_29_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09231_ _09232_/A _09239_/B vssd1 vssd1 vccd1 vccd1 _12365_/A sky130_fd_sc_hd__nor2_8
XANTENNA__06825__B _11029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09162_ reg1_val[5] reg1_val[26] _09180_/S vssd1 vssd1 vccd1 vccd1 _09162_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11061__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08113_ _09472_/A _08199_/B fanout33/X _08649_/B1 vssd1 vssd1 vccd1 vccd1 _08114_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout216_A _09103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09093_ _09669_/B2 _10476_/B _10476_/C _09301_/A fanout56/X vssd1 vssd1 vccd1 vccd1
+ _09094_/B sky130_fd_sc_hd__o32a_1
XFILLER_0_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08044_ _08657_/B fanout84/X fanout80/X _08649_/A2 vssd1 vssd1 vccd1 vccd1 _08045_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07280__A2 _10725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12054__S _12054_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10572__C1 _06958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09995_ _09995_/A _09995_/B vssd1 vssd1 vccd1 vccd1 _09997_/B sky130_fd_sc_hd__xnor2_2
X_08946_ _08946_/A _08946_/B vssd1 vssd1 vccd1 vccd1 _08948_/B sky130_fd_sc_hd__xnor2_2
X_08877_ _12808_/A _08877_/B vssd1 vssd1 vccd1 vccd1 _09010_/A sky130_fd_sc_hd__nor2_2
X_07828_ _07828_/A _07828_/B vssd1 vssd1 vccd1 vccd1 _07935_/B sky130_fd_sc_hd__xor2_1
X_07759_ _08580_/A _07759_/B vssd1 vssd1 vccd1 vccd1 _07763_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10770_ _10770_/A _10770_/B vssd1 vssd1 vccd1 vccd1 _10772_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout31_A fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07099__A2 _10245_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09429_ _09415_/Y _09429_/B _09429_/C _09429_/D vssd1 vssd1 vccd1 vccd1 _09429_/X
+ sky130_fd_sc_hd__and4b_1
X_12440_ _06962_/B _12439_/X _09226_/X vssd1 vssd1 vccd1 vccd1 _12440_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08048__A1 _08576_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08048__B2 _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08599__A2 _08649_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12371_ _12447_/B1 _12417_/B hold241/A vssd1 vssd1 vccd1 vccd1 _12373_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11322_ _11322_/A _11322_/B vssd1 vssd1 vccd1 vccd1 _11324_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07847__A _08454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11253_ _11646_/B _11363_/B hold182/A vssd1 vssd1 vccd1 vccd1 _11254_/C sky130_fd_sc_hd__a21oi_1
X_10204_ _10204_/A _10204_/B vssd1 vssd1 vccd1 vccd1 _10260_/A sky130_fd_sc_hd__xnor2_4
X_11184_ _11946_/B _07171_/A fanout38/X _07013_/X vssd1 vssd1 vccd1 vccd1 _11185_/B
+ sky130_fd_sc_hd__a22o_1
X_10135_ _10135_/A _10135_/B vssd1 vssd1 vccd1 vccd1 _10136_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__12855__A1 _11946_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10066_ _10066_/A _10066_/B vssd1 vssd1 vccd1 vccd1 _10069_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_max_cap9_A _08974_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10968_ _10967_/A _10967_/B _10967_/C vssd1 vssd1 vccd1 vccd1 _10976_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08287__A1 _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08287__B2 _08649_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11830__A2 _09422_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09302__A _09302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12707_ reg1_val[13] _12708_/B vssd1 vssd1 vccd1 vccd1 _12717_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_128_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10899_ _10656_/A _10776_/X _10778_/B vssd1 vssd1 vccd1 vccd1 _10899_/Y sky130_fd_sc_hd__a21oi_2
X_12638_ reg1_val[27] curr_PC[27] _12638_/S vssd1 vssd1 vccd1 vccd1 _12639_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_38_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08039__B2 _08613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08039__A1 _06992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12569_ reg1_val[16] curr_PC[16] _12638_/S vssd1 vssd1 vccd1 vccd1 _12570_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_41_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold206 hold206/A vssd1 vssd1 vccd1 vccd1 hold206/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold217 hold217/A vssd1 vssd1 vccd1 vccd1 hold217/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold228 hold228/A vssd1 vssd1 vccd1 vccd1 hold228/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 hold300/A vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08800_ _08800_/A _08800_/B vssd1 vssd1 vccd1 vccd1 _08800_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_0_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12602__S _12631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09780_ _09780_/A _09780_/B vssd1 vssd1 vccd1 vccd1 _09782_/C sky130_fd_sc_hd__xor2_1
X_06992_ _06992_/A _12644_/A vssd1 vssd1 vccd1 vccd1 _07983_/A sky130_fd_sc_hd__and2_2
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ _08730_/A _08730_/B _10420_/C _10420_/B vssd1 vssd1 vccd1 vccd1 _10668_/B
+ sky130_fd_sc_hd__o211ai_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08662_ _07959_/A _07983_/A _07148_/Y _12642_/A vssd1 vssd1 vccd1 vccd1 _09432_/A
+ sky130_fd_sc_hd__a22o_1
X_07613_ _07614_/A _07614_/B vssd1 vssd1 vccd1 vccd1 _07613_/X sky130_fd_sc_hd__or2_1
XANTENNA_fanout166_A _12322_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08593_ _08593_/A _08593_/B vssd1 vssd1 vccd1 vccd1 _08594_/B sky130_fd_sc_hd__and2_1
XFILLER_0_119_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07544_ _09836_/A _07544_/B vssd1 vssd1 vccd1 vccd1 _07546_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07475_ _07475_/A _07475_/B vssd1 vssd1 vccd1 vccd1 _07534_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_119_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10358__A _11393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09214_ _09206_/X _09213_/X _10295_/S vssd1 vssd1 vccd1 vccd1 _09214_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11034__B1 _11648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09778__A1 _07417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09778__B2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09145_ _09146_/A _09146_/B vssd1 vssd1 vccd1 vccd1 _09711_/A sky130_fd_sc_hd__and2_1
XFILLER_0_16_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09076_ fanout59/X _10245_/B2 _10245_/A1 fanout57/X vssd1 vssd1 vccd1 vccd1 _09077_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08027_ _08065_/B _08027_/B _08027_/C vssd1 vssd1 vccd1 vccd1 _08083_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_102_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08202__A1 _09940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08202__B2 _08561_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09950__A1 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09950__B2 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09978_ _09979_/A _09979_/B vssd1 vssd1 vccd1 vccd1 _09978_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12837__A1 _07269_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08929_ _09834_/A _08929_/B vssd1 vssd1 vccd1 vccd1 _08933_/A sky130_fd_sc_hd__xnor2_1
X_11940_ _12030_/B _11940_/B vssd1 vssd1 vccd1 vccd1 _11957_/A sky130_fd_sc_hd__and2_1
XFILLER_0_98_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11871_ _11872_/A _11872_/B _11872_/C vssd1 vssd1 vccd1 vccd1 _11873_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_79_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10822_ _10821_/A _10818_/X _10819_/X _10821_/Y vssd1 vssd1 vccd1 vccd1 dest_val[11]
+ sky130_fd_sc_hd__a22o_4
X_10753_ _10588_/A _10588_/B _10593_/A vssd1 vssd1 vccd1 vccd1 _10755_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10615__A3 fanout8/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10684_ _11820_/A _10682_/X _10683_/X _09242_/B vssd1 vssd1 vccd1 vccd1 _10684_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_70_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08961__A _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12423_ _10159_/A _09409_/Y _12412_/B _09222_/Y _12422_/Y vssd1 vssd1 vccd1 vccd1
+ _12423_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_63_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12354_ _12429_/A _12354_/B vssd1 vssd1 vccd1 vccd1 _12399_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_62_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11305_ _11183_/A _11183_/B _11180_/A vssd1 vssd1 vccd1 vccd1 _11308_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_77_18 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12285_ _12285_/A _12285_/B vssd1 vssd1 vccd1 vccd1 _12287_/A sky130_fd_sc_hd__nor2_1
XANTENNA__09792__A _10749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11236_ _11809_/A _08751_/X _08753_/X _10788_/A _11235_/Y vssd1 vssd1 vccd1 vccd1
+ _11236_/Y sky130_fd_sc_hd__a311oi_1
XANTENNA__10000__A1 _09707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11167_ _12096_/A _11167_/B vssd1 vssd1 vccd1 vccd1 _11168_/B sky130_fd_sc_hd__xor2_1
X_10118_ _10118_/A _10118_/B vssd1 vssd1 vccd1 vccd1 _10120_/B sky130_fd_sc_hd__xor2_4
X_11098_ _11098_/A _11098_/B vssd1 vssd1 vccd1 vccd1 _11099_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10839__B1 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10049_ _10049_/A _10049_/B vssd1 vssd1 vccd1 vccd1 _10049_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_98_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07260_ _07270_/A _06974_/X _06978_/C _06978_/D _07215_/B vssd1 vssd1 vccd1 vccd1
+ _07262_/B sky130_fd_sc_hd__o41a_4
XFILLER_0_73_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07191_ _07189_/Y _07192_/B vssd1 vssd1 vccd1 vccd1 _07191_/X sky130_fd_sc_hd__and2b_2
XFILLER_0_26_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09901_ reg1_val[4] _07117_/C _11995_/B _09894_/X _09900_/X vssd1 vssd1 vccd1 vccd1
+ _09901_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_1_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12840__B _12862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09832_ _09611_/Y _09614_/B _09619_/A vssd1 vssd1 vccd1 vccd1 _09843_/A sky130_fd_sc_hd__a21o_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12819__A1 _07121_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09763_ _10821_/A _10045_/C vssd1 vssd1 vccd1 vccd1 _09763_/Y sky130_fd_sc_hd__nor2_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06975_ _07237_/A _07215_/A vssd1 vssd1 vccd1 vccd1 _06978_/C sky130_fd_sc_hd__or2_4
X_08714_ _08714_/A _08714_/B vssd1 vssd1 vccd1 vccd1 _08715_/B sky130_fd_sc_hd__and2_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09694_ _09694_/A _09694_/B vssd1 vssd1 vccd1 vccd1 _09696_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08645_ _08646_/A _08646_/C _08646_/B vssd1 vssd1 vccd1 vccd1 _08645_/X sky130_fd_sc_hd__a21o_1
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11472__A _12050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09448__B1 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08576_ _08641_/B _08576_/A2 _09472_/A _08627_/A2 vssd1 vssd1 vccd1 vccd1 _08577_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07527_ _07721_/A _07721_/B vssd1 vssd1 vccd1 vccd1 _07734_/C sky130_fd_sc_hd__or2_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07458_ _07461_/A _07461_/B vssd1 vssd1 vccd1 vccd1 _07458_/X sky130_fd_sc_hd__or2_1
XFILLER_0_9_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09596__B _09596_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07389_ _08199_/B _10599_/A _10500_/A fanout33/X vssd1 vssd1 vccd1 vccd1 _07390_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_115_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07397__A _09341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09128_ _09128_/A _09128_/B vssd1 vssd1 vccd1 vccd1 _09129_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10230__A1 _07171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10230__B2 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09059_ _09060_/A _09060_/B _09060_/C vssd1 vssd1 vccd1 vccd1 _09357_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_20_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12070_ hold278/A _12449_/B1 _12136_/B _12069_/Y _12376_/C1 vssd1 vssd1 vccd1 vccd1
+ _12070_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11021_ _11022_/A _11022_/B vssd1 vssd1 vccd1 vccd1 _11021_/X sky130_fd_sc_hd__or2_1
XANTENNA__09117__A _09834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08021__A _08564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12972_ hold48/X _12971_/B hold250/X vssd1 vssd1 vccd1 vccd1 _13247_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_99_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08956__A _10479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11494__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11923_ _12631_/S _11920_/X _11921_/X _11922_/Y vssd1 vssd1 vccd1 vccd1 dest_val[22]
+ sky130_fd_sc_hd__a22o_4
X_11854_ _11854_/A fanout7/X vssd1 vssd1 vccd1 vccd1 _11854_/X sky130_fd_sc_hd__or2_1
X_10805_ hold213/A _10805_/B vssd1 vssd1 vccd1 vccd1 _10921_/B sky130_fd_sc_hd__or2_1
X_11785_ _11785_/A _11785_/B _11785_/C vssd1 vssd1 vccd1 vccd1 _11786_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_82_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10736_ _11582_/A _10736_/B vssd1 vssd1 vccd1 vccd1 _10737_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12994__B1 _13257_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08662__B2 _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08662__A1 _07959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10667_ _11809_/A _10668_/B _10668_/C _10668_/D vssd1 vssd1 vccd1 vccd1 _10669_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12406_ _12406_/A _12406_/B vssd1 vssd1 vccd1 vccd1 _12406_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13386_ _13390_/CLK _13386_/D vssd1 vssd1 vccd1 vccd1 hold276/A sky130_fd_sc_hd__dfxtp_1
X_10598_ _10599_/A _12087_/B vssd1 vssd1 vccd1 vccd1 _10600_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10221__A1 _10500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07100__A _10479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12337_ _12338_/A _12338_/B vssd1 vssd1 vccd1 vccd1 _12339_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10221__B2 _10221_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12268_ hold224/A _12447_/B1 _12321_/B _11648_/A vssd1 vssd1 vccd1 vccd1 _12269_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09726__S _10297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11219_ _11219_/A _11219_/B vssd1 vssd1 vccd1 vccd1 _11222_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09914__A1 _07417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09914__B2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12660__B _12660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12199_ hold276/A _12199_/B vssd1 vssd1 vccd1 vccd1 _12270_/B sky130_fd_sc_hd__or2_1
XANTENNA__07925__B1 _10338_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06760_ reg2_val[9] _06810_/B vssd1 vssd1 vccd1 vccd1 _06760_/X sky130_fd_sc_hd__and2_2
XFILLER_0_37_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06691_ reg1_val[20] _07016_/A vssd1 vssd1 vccd1 vccd1 _06691_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_78_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08430_ _08407_/A _08407_/B _08429_/X vssd1 vssd1 vccd1 vccd1 _08434_/A sky130_fd_sc_hd__o21bai_4
XFILLER_0_93_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08361_ _08690_/A _08690_/B _08690_/C vssd1 vssd1 vccd1 vccd1 _08691_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_116_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08292_ _06992_/A fanout76/X fanout72/X _08613_/A vssd1 vssd1 vccd1 vccd1 _08293_/B
+ sky130_fd_sc_hd__o22a_2
XANTENNA__07456__A2 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07312_ _07604_/A _07312_/B vssd1 vssd1 vccd1 vccd1 _07325_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_5_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07243_ _07104_/A _07104_/B _07244_/B vssd1 vssd1 vccd1 vccd1 _07243_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_5_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07174_ _07170_/A _07170_/B _12093_/A vssd1 vssd1 vccd1 vccd1 _07174_/X sky130_fd_sc_hd__mux2_2
XANTENNA__07010__A _09673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10763__A2 _10707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10371__A _10950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ _09302_/A _07011_/A fanout8/X _09814_/Y vssd1 vssd1 vccd1 vccd1 _09817_/B
+ sky130_fd_sc_hd__o31ai_4
X_06958_ _06958_/A _06958_/B vssd1 vssd1 vccd1 vccd1 dest_mask[1] sky130_fd_sc_hd__nand2_8
XANTENNA__12268__A2 _12447_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09746_ _09745_/B _09746_/B vssd1 vssd1 vccd1 vccd1 _09746_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__09669__B1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _09677_/A _11497_/A vssd1 vssd1 vccd1 vccd1 _09683_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10279__B2 _10136_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06889_ _06963_/B _06888_/X _06879_/X vssd1 vssd1 vccd1 vccd1 _06889_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07144__A1 _11134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08628_ _09302_/A _08628_/B vssd1 vssd1 vccd1 vccd1 _08628_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08559_ _06992_/A _09770_/B2 _09940_/B2 _08613_/A vssd1 vssd1 vccd1 vccd1 _08560_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_119_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11570_ _07051_/X _07171_/A fanout38/X _12169_/A vssd1 vssd1 vccd1 vccd1 _11571_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12976__B1 _13257_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout8_A fanout8/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10521_ _10521_/A _10521_/B vssd1 vssd1 vccd1 vccd1 _10534_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10451__A1 _11752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13240_ hold287/A _13239_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13240_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_92_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10452_ curr_PC[9] _10699_/C vssd1 vssd1 vccd1 vccd1 _10452_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_33_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13171_ hold272/X _13223_/A2 _13170_/X _13171_/B2 vssd1 vssd1 vccd1 vccd1 hold273/A
+ sky130_fd_sc_hd__a22o_1
X_10383_ _10383_/A _10383_/B vssd1 vssd1 vccd1 vccd1 _10397_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_20_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12122_ _12184_/B _12123_/B vssd1 vssd1 vccd1 vccd1 _12122_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_32_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12053_ _06700_/A _11979_/X _11995_/A vssd1 vssd1 vccd1 vccd1 _12053_/Y sky130_fd_sc_hd__a21oi_1
X_11004_ _11004_/A _11004_/B vssd1 vssd1 vccd1 vccd1 _11006_/C sky130_fd_sc_hd__xnor2_1
X_12955_ hold24/X hold266/X vssd1 vssd1 vccd1 vccd1 _13211_/B sky130_fd_sc_hd__nand2b_1
X_11906_ _10575_/X _11905_/X _12444_/B vssd1 vssd1 vccd1 vccd1 _11906_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08332__B1 _08561_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12886_ hold52/X hold262/X vssd1 vssd1 vccd1 vccd1 _12886_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12416__C1 _12416_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07150__A4 _07143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11837_ curr_PC[21] _11837_/B vssd1 vssd1 vccd1 vccd1 _12003_/C sky130_fd_sc_hd__and2_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _07175_/Y fanout17/X _12335_/A _07171_/Y vssd1 vssd1 vccd1 vccd1 _11769_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10719_ _10719_/A _10719_/B vssd1 vssd1 vccd1 vccd1 _10720_/B sky130_fd_sc_hd__nor2_1
XANTENNA__12655__B _12655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06653__B _06675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11699_ _11793_/A _11699_/B vssd1 vssd1 vccd1 vccd1 _11701_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_113_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13369_ _13369_/CLK _13369_/D vssd1 vssd1 vccd1 vccd1 hold252/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11942__B2 _12009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11942__A1 _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07765__A _08564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07930_ _08003_/A _08003_/B vssd1 vssd1 vccd1 vccd1 _07930_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_48_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07861_ _07861_/A _07861_/B vssd1 vssd1 vccd1 vccd1 _07937_/B sky130_fd_sc_hd__xnor2_1
X_06812_ _06815_/A _06817_/B1 _12650_/B _06810_/X vssd1 vssd1 vccd1 vccd1 _07149_/A
+ sky130_fd_sc_hd__a31o_4
X_09600_ _09583_/Y _09584_/X _09597_/X _09599_/X vssd1 vssd1 vccd1 vccd1 _09600_/X
+ sky130_fd_sc_hd__o211a_1
X_07792_ _09667_/A _07792_/B vssd1 vssd1 vccd1 vccd1 _07826_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11458__B1 _12638_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06743_ _11039_/S _06743_/B vssd1 vssd1 vccd1 vccd1 _11022_/A sky130_fd_sc_hd__or2_2
X_09531_ _09531_/A _09531_/B vssd1 vssd1 vccd1 vccd1 _09544_/A sky130_fd_sc_hd__xor2_4
XANTENNA__13007__A _13019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06674_ _06674_/A vssd1 vssd1 vccd1 vccd1 _06902_/A sky130_fd_sc_hd__inv_2
X_09462_ _09463_/A _09463_/B _09463_/C vssd1 vssd1 vccd1 vccd1 _09464_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_80_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09393_ _09385_/X _09392_/X _11028_/S vssd1 vssd1 vccd1 vccd1 _09393_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07005__A _09947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08413_ _10950_/A _08449_/B _08450_/A vssd1 vssd1 vccd1 vccd1 _08427_/B sky130_fd_sc_hd__o21a_1
XANTENNA_fanout246_A _06958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08344_ _08392_/A _08392_/B _08334_/A vssd1 vssd1 vccd1 vccd1 _08345_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_117_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08275_ _08275_/A _08275_/B vssd1 vssd1 vccd1 vccd1 _08280_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_104_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07226_ _07226_/A _07226_/B vssd1 vssd1 vccd1 vccd1 _07227_/B sky130_fd_sc_hd__nor2_1
Xclkbuf_4_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13373_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07157_ _07158_/B _12158_/A vssd1 vssd1 vccd1 vccd1 _07157_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_42_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09051__A1 _07554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09051__B2 _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07088_ _07088_/A _07088_/B vssd1 vssd1 vccd1 vccd1 _07088_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__10813__B _12422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout110 _07237_/Y vssd1 vssd1 vccd1 vccd1 _10500_/A sky130_fd_sc_hd__buf_4
Xfanout121 _08334_/A vssd1 vssd1 vccd1 vccd1 _09667_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout165 _12447_/B1 vssd1 vssd1 vccd1 vccd1 _11990_/A1 sky130_fd_sc_hd__buf_4
Xfanout132 _07098_/X vssd1 vssd1 vccd1 vccd1 _10245_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout154 _07015_/X vssd1 vssd1 vccd1 vccd1 _09301_/A sky130_fd_sc_hd__clkbuf_8
Xfanout143 _09325_/A vssd1 vssd1 vccd1 vccd1 _08649_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout198 _12144_/A1 vssd1 vssd1 vccd1 vccd1 _12421_/A1 sky130_fd_sc_hd__buf_4
XANTENNA__12520__S _12520_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout187 _13257_/A2 vssd1 vssd1 vccd1 vccd1 _13254_/A2 sky130_fd_sc_hd__buf_4
Xfanout176 _10159_/A vssd1 vssd1 vccd1 vccd1 _09211_/S sky130_fd_sc_hd__clkbuf_8
X_09729_ _09727_/X _09728_/X _10295_/S vssd1 vssd1 vccd1 vccd1 _09729_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout61_A _07019_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12740_ _12755_/B _12740_/B vssd1 vssd1 vccd1 vccd1 _12742_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_96_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _12671_/A _12671_/B vssd1 vssd1 vccd1 vccd1 _12672_/B sky130_fd_sc_hd__or2_2
X_11622_ _11436_/X _11800_/A _11621_/X vssd1 vssd1 vccd1 vccd1 _11622_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_65_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09814__B1 _09302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11553_ _11829_/B _11995_/B _11553_/S vssd1 vssd1 vccd1 vccd1 _11554_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10276__A _10276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11484_ _11484_/A _11484_/B vssd1 vssd1 vccd1 vccd1 _11486_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10504_ _10504_/A _10504_/B vssd1 vssd1 vccd1 vccd1 _10515_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_122_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13223_ hold276/X _13223_/A2 _13222_/X _13223_/B2 vssd1 vssd1 vccd1 vccd1 hold277/A
+ sky130_fd_sc_hd__a22o_1
X_10435_ _11990_/A1 _10565_/B hold217/A vssd1 vssd1 vccd1 vccd1 _10435_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13154_ _13154_/A _13154_/B vssd1 vssd1 vccd1 vccd1 _13154_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__11924__A1 _12050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12105_ _12105_/A _12105_/B vssd1 vssd1 vccd1 vccd1 _12106_/B sky130_fd_sc_hd__or2_1
X_10366_ _10366_/A _10366_/B vssd1 vssd1 vccd1 vccd1 _10367_/B sky130_fd_sc_hd__xor2_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ _11929_/A _13089_/A2 hold109/X vssd1 vssd1 vccd1 vccd1 hold110/A sky130_fd_sc_hd__o21a_1
X_10297_ _09725_/X _09728_/X _10297_/S vssd1 vssd1 vccd1 vccd1 _10297_/X sky130_fd_sc_hd__mux2_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12036_ _12036_/A _12036_/B _12036_/C vssd1 vssd1 vccd1 vccd1 _12037_/B sky130_fd_sc_hd__nand3_1
XANTENNA__09345__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11152__A2 _12422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06648__B _12689_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12938_ hold20/X hold272/X vssd1 vssd1 vccd1 vccd1 _13173_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_34_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08856__B2 _09298_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08856__A1 _09298_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12869_ _08859_/Y _12871_/A2 hold27/X _13246_/A vssd1 vssd1 vccd1 vccd1 _13295_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08871__A4 _12779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09975__A _11582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07831__A2 _07020_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08060_ _08070_/B _08070_/A vssd1 vssd1 vccd1 vccd1 _08072_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_114_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12168__B2 _07051_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12168__A1 _07316_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07011_ _07011_/A _07011_/B vssd1 vssd1 vccd1 vccd1 _07011_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11915__A1 _07014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07595__A1 _12224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09584__A2 _12322_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08962_ _08199_/B _11198_/A _11093_/A fanout33/X vssd1 vssd1 vccd1 vccd1 _08963_/B
+ sky130_fd_sc_hd__o22a_1
X_07913_ _07913_/A _07913_/B _07913_/C vssd1 vssd1 vccd1 vccd1 _07918_/A sky130_fd_sc_hd__and3_1
X_08893_ _08893_/A _08893_/B _08893_/C vssd1 vssd1 vccd1 vccd1 _08894_/B sky130_fd_sc_hd__and3_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07844_ _07863_/A _07863_/B vssd1 vssd1 vccd1 vccd1 _07844_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_98_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07898__A2 _08112_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06783__C_N _12670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07775_ _07777_/A _07777_/B vssd1 vssd1 vccd1 vccd1 _07775_/Y sky130_fd_sc_hd__nor2_1
X_06726_ reg1_val[16] _06727_/B vssd1 vssd1 vccd1 vccd1 _06726_/X sky130_fd_sc_hd__and2_1
XFILLER_0_79_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09514_ _11284_/A _09514_/B vssd1 vssd1 vccd1 vccd1 _09518_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08847__A1 _08199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08847__B2 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06657_ reg1_val[24] _06658_/B vssd1 vssd1 vccd1 vccd1 _12071_/S sky130_fd_sc_hd__nand2_1
X_09445_ _09765_/A _09765_/B _10049_/A vssd1 vssd1 vccd1 vccd1 _09555_/A sky130_fd_sc_hd__o21ai_1
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06588_ instruction[0] instruction[1] instruction[2] pred_val vssd1 vssd1 vccd1 vccd1
+ _06588_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_46_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09376_ _10004_/A _09376_/B vssd1 vssd1 vccd1 vccd1 _09765_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_105_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08327_ _08327_/A _08327_/B vssd1 vssd1 vccd1 vccd1 _08358_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09272__B2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09272__A1 _07417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10957__A2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08258_ _08317_/B _08317_/A vssd1 vssd1 vccd1 vccd1 _08258_/Y sky130_fd_sc_hd__nand2b_1
X_07209_ _07212_/A _07212_/B vssd1 vssd1 vccd1 vccd1 _11284_/A sky130_fd_sc_hd__and2_4
XANTENNA__12159__B2 _12224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10220_ _10220_/A _10220_/B vssd1 vssd1 vccd1 vccd1 _10257_/A sky130_fd_sc_hd__xnor2_1
X_08189_ _08540_/B _10221_/B2 _09770_/B2 _08515_/A2 vssd1 vssd1 vccd1 vccd1 _08190_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11382__A2 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10151_ _11630_/A _10151_/B _10151_/C vssd1 vssd1 vccd1 vccd1 _10151_/X sky130_fd_sc_hd__or3_1
XFILLER_0_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10082_ fanout43/X _10234_/A2 _10725_/A fanout41/X vssd1 vssd1 vccd1 vccd1 _10083_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10984_ _10984_/A _10984_/B _10984_/C vssd1 vssd1 vccd1 vccd1 _10986_/A sky130_fd_sc_hd__and3_1
XANTENNA__12095__B1 _08974_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12723_ reg1_val[16] _12755_/B vssd1 vssd1 vccd1 vccd1 _12726_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_127_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12486__A _12660_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07510__B2 _10500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07510__A1 _08457_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12654_ reg1_val[3] _12655_/B vssd1 vssd1 vccd1 vccd1 _12654_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_127_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11605_ _11606_/A _11606_/B vssd1 vssd1 vccd1 vccd1 _11705_/A sky130_fd_sc_hd__or2_1
X_12585_ _12597_/A _12597_/B _12598_/B vssd1 vssd1 vccd1 vccd1 _12586_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_108_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10948__A2 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11536_ _11536_/A _11536_/B vssd1 vssd1 vccd1 vccd1 _11536_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_108_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13206_ _13210_/A hold269/X vssd1 vssd1 vccd1 vccd1 _13382_/D sky130_fd_sc_hd__and2_1
X_11467_ _11648_/A _11462_/X _11463_/Y _11466_/X vssd1 vssd1 vccd1 vccd1 _11467_/X
+ sky130_fd_sc_hd__o31a_1
Xmax_cap118 _07195_/X vssd1 vssd1 vccd1 vccd1 _10234_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_33_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11398_ _11398_/A _11398_/B vssd1 vssd1 vccd1 vccd1 _11399_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_110_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10418_ _10326_/X _10453_/B _10417_/Y vssd1 vssd1 vccd1 vccd1 _10418_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10453__B _10453_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07577__A1 _10337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13137_ _13147_/A _13137_/B vssd1 vssd1 vccd1 vccd1 _13368_/D sky130_fd_sc_hd__and2_1
X_10349_ _07092_/B fanout8/X _10479_/A vssd1 vssd1 vccd1 vccd1 _10349_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__07577__B2 _07959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ hold135/X _12805_/A _13101_/A2 hold79/X _13039_/A vssd1 vssd1 vccd1 vccd1
+ hold136/A sky130_fd_sc_hd__o221a_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12019_ _12096_/A _12019_/B vssd1 vssd1 vccd1 vccd1 _12021_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12322__A1 _12322_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11125__A2 _11124_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07560_ _07681_/A _07681_/B _07539_/X vssd1 vssd1 vccd1 vccd1 _07568_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_88_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08874__A _12336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09230_ _12144_/A1 _09229_/X _06894_/Y vssd1 vssd1 vccd1 vccd1 _09241_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07491_ _07490_/A _07533_/A vssd1 vssd1 vccd1 vccd1 _07566_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_0_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09161_ reg1_val[4] reg1_val[27] _09180_/S vssd1 vssd1 vccd1 vccd1 _09161_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11061__B2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11061__A1 _12009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09092_ _09673_/A _09092_/B vssd1 vssd1 vccd1 vccd1 _09099_/A sky130_fd_sc_hd__xor2_1
X_08112_ _09404_/S _08112_/B vssd1 vssd1 vccd1 vccd1 _08159_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_16_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08043_ _08046_/A _08046_/B vssd1 vssd1 vccd1 vccd1 _08043_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout111_A _07233_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08114__A _10092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10021__C1 _11029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09994_ _09995_/B _09995_/A vssd1 vssd1 vccd1 vccd1 _09994_/Y sky130_fd_sc_hd__nand2b_1
X_08945_ _08946_/B _08946_/A vssd1 vssd1 vccd1 vccd1 _09060_/A sky130_fd_sc_hd__nand2b_1
X_08876_ _08876_/A _08876_/B vssd1 vssd1 vccd1 vccd1 _08876_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_98_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07827_ _07828_/A _07828_/B vssd1 vssd1 vccd1 vccd1 _07827_/Y sky130_fd_sc_hd__nor2_1
X_07758_ _08598_/B fanout84/X fanout80/X _08538_/A1 vssd1 vssd1 vccd1 vccd1 _07759_/B
+ sky130_fd_sc_hd__o22a_1
X_06709_ instruction[28] _06716_/B vssd1 vssd1 vccd1 vccd1 _12655_/B sky130_fd_sc_hd__and2_4
XFILLER_0_94_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11824__B1 _12376_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07689_ _08540_/B fanout80/X fanout76/X _08515_/A2 vssd1 vssd1 vccd1 vccd1 _07690_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_109_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09428_ _09418_/A _12420_/A0 _09422_/X _09426_/X _09427_/X vssd1 vssd1 vccd1 vccd1
+ _09429_/D sky130_fd_sc_hd__o2111a_1
XFILLER_0_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09245__A1 _09728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08048__A2 _08199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09359_ _09126_/A _09126_/B _09124_/X vssd1 vssd1 vccd1 vccd1 _09361_/B sky130_fd_sc_hd__a21oi_2
X_12370_ hold227/A _12370_/B vssd1 vssd1 vccd1 vccd1 _12417_/B sky130_fd_sc_hd__or2_1
XANTENNA__13041__A2 _13101_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11321_ _11214_/A _11213_/Y _11211_/X vssd1 vssd1 vccd1 vccd1 _11322_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_105_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12001__B1 _11977_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11252_ hold182/A _11646_/B _11363_/B vssd1 vssd1 vccd1 vccd1 _11254_/B sky130_fd_sc_hd__and3_1
XFILLER_0_120_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11183_ _11183_/A _11183_/B vssd1 vssd1 vccd1 vccd1 _11195_/A sky130_fd_sc_hd__xor2_2
X_10203_ _10203_/A _10203_/B vssd1 vssd1 vccd1 vccd1 _10204_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_30_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10134_ _10134_/A _10134_/B vssd1 vssd1 vccd1 vccd1 _10135_/B sky130_fd_sc_hd__xor2_4
XANTENNA__12855__A2 _12863_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10065_ _10065_/A _10065_/B vssd1 vssd1 vccd1 vccd1 _10066_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10967_ _10967_/A _10967_/B _10967_/C vssd1 vssd1 vccd1 vccd1 _10976_/A sky130_fd_sc_hd__and3_1
XFILLER_0_97_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06926__B _06926_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08287__A2 _08411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10898_ _10898_/A _10898_/B vssd1 vssd1 vccd1 vccd1 _11120_/A sky130_fd_sc_hd__or2_4
XFILLER_0_85_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13105__A _13147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12706_ _12711_/B _12706_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[12] sky130_fd_sc_hd__and2_4
XFILLER_0_128_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12637_ _12634_/B _12636_/B _12634_/A vssd1 vssd1 vccd1 vccd1 _12640_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_66_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08039__A2 _09661_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12568_ _12572_/B _12568_/B vssd1 vssd1 vccd1 vccd1 new_PC[15] sky130_fd_sc_hd__and2_4
XANTENNA__11043__B2 _10159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11519_ _11616_/A _11519_/B vssd1 vssd1 vccd1 vccd1 _11522_/A sky130_fd_sc_hd__nand2_1
Xhold207 hold207/A vssd1 vssd1 vccd1 vccd1 hold207/X sky130_fd_sc_hd__dlygate4sd3_1
X_12499_ reg1_val[6] curr_PC[6] _12520_/S vssd1 vssd1 vccd1 vccd1 _12501_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_40_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold229 hold229/A vssd1 vssd1 vccd1 vccd1 hold229/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 hold218/A vssd1 vssd1 vccd1 vccd1 hold218/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06991_ _07046_/B _06991_/B vssd1 vssd1 vccd1 vccd1 _06991_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__13099__A2 _12820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ _08730_/A _08730_/B vssd1 vssd1 vccd1 vccd1 _10552_/C sky130_fd_sc_hd__or2_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08661_ _08661_/A _08667_/S vssd1 vssd1 vccd1 vccd1 _08664_/B sky130_fd_sc_hd__xor2_1
X_07612_ _09947_/A _07612_/B vssd1 vssd1 vccd1 vccd1 _07614_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12838__B _12862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08592_ _08592_/A _08592_/B vssd1 vssd1 vccd1 vccd1 _08678_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11742__B _11829_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07543_ _07134_/Y _07959_/B fanout29/X _07166_/Y vssd1 vssd1 vccd1 vccd1 _07544_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13015__A _13019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout159_A _11892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07474_ _07475_/A _07475_/B vssd1 vssd1 vccd1 vccd1 _07492_/B sky130_fd_sc_hd__and2_1
XANTENNA__07013__A _07014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09213_ _09209_/X _09212_/X _09727_/S vssd1 vssd1 vccd1 vccd1 _09213_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09144_ _09144_/A _09144_/B vssd1 vssd1 vccd1 vccd1 _09146_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__09778__A2 _07232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10793__B1 _09225_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09075_ _09075_/A _09075_/B vssd1 vssd1 vccd1 vccd1 _09079_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_114_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1 fanout2/X vssd1 vssd1 vccd1 vccd1 fanout1/X sky130_fd_sc_hd__buf_6
XANTENNA__07159__S _12224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08026_ _08065_/A _07992_/C _07992_/B vssd1 vssd1 vccd1 vccd1 _08027_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08202__A2 _08484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09950__A2 fanout86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ _09828_/A _09828_/B _09826_/Y vssd1 vssd1 vccd1 vccd1 _09979_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__12837__A2 _12863_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ fanout46/X _07217_/Y _10500_/A _07830_/B vssd1 vssd1 vccd1 vccd1 _08929_/B
+ sky130_fd_sc_hd__o22a_1
X_08859_ _08973_/C _08860_/B vssd1 vssd1 vccd1 vccd1 _08859_/Y sky130_fd_sc_hd__xnor2_4
X_11870_ _11870_/A _11870_/B vssd1 vssd1 vccd1 vccd1 _11872_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10821_ _10821_/A _10821_/B vssd1 vssd1 vccd1 vccd1 _10821_/Y sky130_fd_sc_hd__nor2_1
X_10752_ _10874_/B _10752_/B vssd1 vssd1 vccd1 vccd1 _10755_/A sky130_fd_sc_hd__nor2_1
XANTENNA__06746__B _07195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08019__A _08580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13014__A2 _13171_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12422_ _12422_/A _12422_/B vssd1 vssd1 vccd1 vccd1 _12422_/Y sky130_fd_sc_hd__nor2_1
X_10683_ _10678_/Y _10679_/X _12064_/S vssd1 vssd1 vccd1 vccd1 _10683_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12353_ _11806_/B _12115_/A _12350_/Y _12351_/X _12352_/X vssd1 vssd1 vccd1 vccd1
+ _12354_/B sky130_fd_sc_hd__o311a_1
XFILLER_0_62_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11304_ _11304_/A _11304_/B vssd1 vssd1 vccd1 vccd1 _11313_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_105_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12284_ _12284_/A _12284_/B _12284_/C vssd1 vssd1 vccd1 vccd1 _12285_/B sky130_fd_sc_hd__and3_1
X_11235_ _11809_/A _08751_/X _08753_/X vssd1 vssd1 vccd1 vccd1 _11235_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11166_ _11779_/A fanout43/X fanout41/X _11764_/A vssd1 vssd1 vccd1 vccd1 _11167_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10000__A2 _09707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11097_ _11098_/A _11098_/B vssd1 vssd1 vccd1 vccd1 _11097_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_93_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12004__A _12631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_14_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13396_/CLK sky130_fd_sc_hd__clkbuf_8
X_10117_ _09933_/A _09932_/B _09930_/X vssd1 vssd1 vccd1 vccd1 _10118_/B sky130_fd_sc_hd__a21o_1
XANTENNA__10839__A1 _10944_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09154__A0 _12644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10048_ _09910_/B _10324_/A vssd1 vssd1 vccd1 vccd1 _10049_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_117_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10839__B2 _07097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10459__A _11284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09313__A _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11999_ _11990_/Y _11991_/X _11994_/X _11998_/X vssd1 vssd1 vccd1 vccd1 _11999_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07190_ _09667_/A _07200_/C vssd1 vssd1 vccd1 vccd1 _07192_/B sky130_fd_sc_hd__nand2_2
XANTENNA__12213__B1 _12365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09900_ _12444_/B _12446_/C1 _09899_/X _11554_/A _06796_/A vssd1 vssd1 vccd1 vccd1
+ _09900_/X sky130_fd_sc_hd__a32o_1
XFILLER_0_22_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09831_ _09831_/A _09831_/B vssd1 vssd1 vccd1 vccd1 _09845_/A sky130_fd_sc_hd__xnor2_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06974_ _07133_/A _06974_/B vssd1 vssd1 vccd1 vccd1 _06974_/X sky130_fd_sc_hd__or2_2
X_09762_ curr_PC[3] _09762_/B vssd1 vssd1 vccd1 vccd1 _10045_/C sky130_fd_sc_hd__and2_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12819__A2 _13101_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08713_ _08664_/A _09556_/B _08664_/B vssd1 vssd1 vccd1 vccd1 _08714_/B sky130_fd_sc_hd__o21ai_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout276_A _13162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09693_ _09511_/A _09511_/B _09509_/Y vssd1 vssd1 vccd1 vccd1 _09696_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08644_ _08646_/A _08646_/C _08646_/B vssd1 vssd1 vccd1 vccd1 _08671_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11472__B _11567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09448__A1 _07283_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08575_ _08575_/A _08575_/B vssd1 vssd1 vccd1 vccd1 _08608_/B sky130_fd_sc_hd__xnor2_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12452__B1 _11554_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09448__B2 _09934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07459__B1 _09661_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07526_ _07526_/A _07526_/B vssd1 vssd1 vccd1 vccd1 _07721_/B sky130_fd_sc_hd__xnor2_1
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07457_ _09947_/A _07457_/B vssd1 vssd1 vccd1 vccd1 _07461_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07388_ _07388_/A _07388_/B vssd1 vssd1 vccd1 vccd1 _07400_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_17_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09127_ _09128_/A _09128_/B vssd1 vssd1 vccd1 vccd1 _09127_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10230__A2 _07262_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07631__B1 _09940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09058_ _09058_/A _09058_/B vssd1 vssd1 vccd1 vccd1 _09060_/C sky130_fd_sc_hd__or2_1
XFILLER_0_13_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08009_ _08009_/A _08009_/B vssd1 vssd1 vccd1 vccd1 _08075_/B sky130_fd_sc_hd__nand2_2
XANTENNA_fanout91_A _11398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11020_ _06842_/X _11019_/X _11813_/S vssd1 vssd1 vccd1 vccd1 _11022_/B sky130_fd_sc_hd__mux2_1
XANTENNA__11191__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12971_ hold48/X _12971_/B vssd1 vssd1 vccd1 vccd1 _12973_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11494__B2 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11494__A1 _11868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11922_ curr_PC[22] _12003_/C _06958_/A vssd1 vssd1 vccd1 vccd1 _11922_/Y sky130_fd_sc_hd__a21oi_1
X_11853_ _12093_/A _11853_/B vssd1 vssd1 vccd1 vccd1 _11857_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_86_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09439__A1 _10159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10804_ _12064_/S _10803_/X _10800_/X vssd1 vssd1 vccd1 vccd1 _10804_/X sky130_fd_sc_hd__o21a_1
X_11784_ _11785_/A _11785_/B _11785_/C vssd1 vssd1 vccd1 vccd1 _11878_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12443__B1 _12365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08972__A _09673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10735_ _12087_/A fanout28/X fanout26/X _12009_/A vssd1 vssd1 vccd1 vccd1 _10736_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12494__A _12665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10666_ _11538_/A _11271_/A _11050_/A _09150_/X vssd1 vssd1 vccd1 vccd1 _10666_/X
+ sky130_fd_sc_hd__a31o_1
X_13385_ _13385_/CLK _13385_/D vssd1 vssd1 vccd1 vccd1 hold278/A sky130_fd_sc_hd__dfxtp_1
X_12405_ _12406_/A _12404_/X _11637_/A vssd1 vssd1 vccd1 vccd1 _12405_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10597_ _10597_/A _10597_/B vssd1 vssd1 vccd1 vccd1 _10600_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__10221__A2 _08877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12336_ _12336_/A _12336_/B vssd1 vssd1 vccd1 vccd1 _12338_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12267_ _12447_/B1 _12321_/B hold224/A vssd1 vssd1 vccd1 vccd1 _12269_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__11838__A _12471_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11218_ _11219_/A _11219_/B vssd1 vssd1 vccd1 vccd1 _11331_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13171__B2 _13171_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12198_ _12444_/B _10016_/Y _12197_/X _12446_/C1 vssd1 vssd1 vccd1 vccd1 _12211_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09914__A2 _10725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11149_ hold193/A _11646_/B _11251_/B _11648_/A vssd1 vssd1 vccd1 vccd1 _11149_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11721__A2 _11720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07925__B2 _08515_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07925__A1 _08540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06690_ _07016_/A reg1_val[20] vssd1 vssd1 vccd1 vccd1 _11742_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__07689__B1 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08360_ _08360_/A _08360_/B vssd1 vssd1 vccd1 vccd1 _08690_/C sky130_fd_sc_hd__xnor2_1
X_07311_ fanout68/X _08657_/B _08649_/A2 fanout65/X vssd1 vssd1 vccd1 vccd1 _07312_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08291_ _08350_/A _08350_/B vssd1 vssd1 vccd1 vccd1 _08311_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_116_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07242_ _07242_/A _07242_/B vssd1 vssd1 vccd1 vccd1 _07244_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_27_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12198__C1 _12446_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07173_ _10297_/S _07173_/B vssd1 vssd1 vccd1 vccd1 _07173_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_42_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09218__A _09218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09814_ _07011_/B fanout8/X _09302_/A vssd1 vssd1 vccd1 vccd1 _09814_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_94_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10920__B1 _11820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06957_ _12359_/A is_load _06723_/A _06954_/X vssd1 vssd1 vccd1 vccd1 _06958_/B sky130_fd_sc_hd__a22o_2
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09745_ _09746_/B _09745_/B vssd1 vssd1 vccd1 vccd1 _09745_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__09669__B2 _09669_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09669__A1 _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06888_ _12406_/A _06887_/X _06865_/X vssd1 vssd1 vccd1 vccd1 _06888_/X sky130_fd_sc_hd__a21o_1
X_09676_ _09676_/A _09676_/B vssd1 vssd1 vccd1 vccd1 _09685_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__06577__A _06577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10684__C1 _09242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07144__A2 _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08627_ _09404_/S _08627_/A2 _08649_/B1 _08641_/B vssd1 vssd1 vccd1 vccd1 _08628_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_96_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08558_ _08564_/A _08564_/B vssd1 vssd1 vccd1 vccd1 _08558_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08489_ _08496_/A _08496_/B vssd1 vssd1 vccd1 vccd1 _08489_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_37_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07509_ _08454_/A _07509_/B vssd1 vssd1 vccd1 vccd1 _07515_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10520_ _10519_/B _10519_/C _10519_/A vssd1 vssd1 vccd1 vccd1 _10521_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10451_ _11752_/S _10447_/X _10450_/X vssd1 vssd1 vccd1 vccd1 dest_val[8] sky130_fd_sc_hd__o21ai_4
XFILLER_0_122_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13170_ hold270/X _13169_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13170_/X sky130_fd_sc_hd__mux2_1
X_10382_ _10380_/Y _10382_/B vssd1 vssd1 vccd1 vccd1 _10398_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_32_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12121_ _12184_/A _12050_/X _11892_/A vssd1 vssd1 vccd1 vccd1 _12123_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12052_ _11892_/A _12184_/A _12050_/X _09149_/Y vssd1 vssd1 vccd1 vccd1 _12052_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA__11164__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11003_ _11004_/A _11004_/B vssd1 vssd1 vccd1 vccd1 _11117_/B sky130_fd_sc_hd__or2_1
XANTENNA__10911__B1 _11637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08967__A _09667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12954_ _13207_/A _12953_/B _12884_/X vssd1 vssd1 vccd1 vccd1 _13212_/A sky130_fd_sc_hd__a21o_1
XANTENNA__11393__A _11393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11467__A1 _11648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11905_ _11905_/A _11905_/B vssd1 vssd1 vccd1 vccd1 _11905_/X sky130_fd_sc_hd__xor2_1
XANTENNA__08332__B2 _08515_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08332__A1 _08540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12885_ hold274/A hold34/X vssd1 vssd1 vccd1 vccd1 _13202_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_59_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11836_ curr_PC[21] _11837_/B vssd1 vssd1 vccd1 vccd1 _11838_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _11767_/A _11767_/B vssd1 vssd1 vccd1 vccd1 _11776_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_55_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06934__B _06944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10718_ _10719_/A _10719_/B vssd1 vssd1 vccd1 vccd1 _10720_/A sky130_fd_sc_hd__and2_1
XANTENNA__10442__A2 _09422_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07843__A0 _09834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11698_ _11698_/A _11698_/B _11698_/C vssd1 vssd1 vccd1 vccd1 _11699_/B sky130_fd_sc_hd__and3_1
XFILLER_0_83_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08207__A _10207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10649_ _10649_/A _10649_/B vssd1 vssd1 vccd1 vccd1 _10651_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13368_ _13369_/CLK _13368_/D vssd1 vssd1 vccd1 vccd1 hold281/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11942__A2 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12319_ _12444_/B _12319_/B vssd1 vssd1 vccd1 vccd1 _12319_/X sky130_fd_sc_hd__or2_1
XANTENNA__11287__B _11288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13299_ _13304_/CLK _13299_/D vssd1 vssd1 vccd1 vccd1 hold237/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08877__A _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08020__B1 _08501_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07860_ _07883_/A _07883_/B vssd1 vssd1 vccd1 vccd1 _07937_/A sky130_fd_sc_hd__nor2_1
X_06811_ _06815_/A _06817_/B1 _12650_/B _06810_/X vssd1 vssd1 vccd1 vccd1 _09728_/S
+ sky130_fd_sc_hd__a31oi_4
X_07791_ _07217_/Y _08289_/B fanout75/X _07221_/X vssd1 vssd1 vccd1 vccd1 _07792_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11458__A1 _07097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06742_ reg1_val[13] _11038_/A vssd1 vssd1 vccd1 vccd1 _06743_/B sky130_fd_sc_hd__nor2_1
X_09530_ _09530_/A _09530_/B vssd1 vssd1 vccd1 vccd1 _09531_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_78_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07126__A2 _12740_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09520__B1 _07274_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09461_ _09461_/A _09461_/B vssd1 vssd1 vccd1 vccd1 _09463_/C sky130_fd_sc_hd__xnor2_1
X_06673_ _06673_/A _12313_/A _06673_/C _06672_/X vssd1 vssd1 vccd1 vccd1 _06674_/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_93_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09392_ _09388_/X _10018_/B _10294_/S vssd1 vssd1 vccd1 vccd1 _09392_/X sky130_fd_sc_hd__mux2_1
X_08412_ _08449_/A _08449_/B vssd1 vssd1 vccd1 vccd1 _08450_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_117_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12846__B _12862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09823__A1 _09673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09501__A _09672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08343_ _08393_/A _08393_/B _08339_/X vssd1 vssd1 vccd1 vccd1 _08367_/A sky130_fd_sc_hd__o21a_1
XANTENNA__10969__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout239_A _08502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08274_ _08282_/A _08282_/B _08233_/Y vssd1 vssd1 vccd1 vccd1 _08280_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_116_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07225_ _07226_/A _07226_/B vssd1 vssd1 vccd1 vccd1 _07227_/A sky130_fd_sc_hd__and2_1
XFILLER_0_104_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07156_ _07155_/A _07155_/B _07155_/C vssd1 vssd1 vccd1 vccd1 _12158_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09051__A2 _10337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07087_ _07087_/A _07088_/B vssd1 vssd1 vccd1 vccd1 _07983_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_42_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout122 _08334_/A vssd1 vssd1 vccd1 vccd1 _11179_/A sky130_fd_sc_hd__clkbuf_16
Xfanout100 _07088_/Y vssd1 vssd1 vccd1 vccd1 _09661_/B2 sky130_fd_sc_hd__buf_8
Xfanout111 _07233_/Y vssd1 vssd1 vccd1 vccd1 _08457_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout144 _07149_/Y vssd1 vssd1 vccd1 vccd1 _09325_/A sky130_fd_sc_hd__buf_4
Xfanout155 _09669_/B2 vssd1 vssd1 vccd1 vccd1 _08641_/B sky130_fd_sc_hd__buf_6
Xfanout133 _10245_/B2 vssd1 vssd1 vccd1 vccd1 _08540_/B sky130_fd_sc_hd__clkbuf_8
Xfanout166 _12322_/A1 vssd1 vssd1 vccd1 vccd1 _12447_/B1 sky130_fd_sc_hd__buf_4
Xfanout199 _09224_/X vssd1 vssd1 vccd1 vccd1 _12144_/A1 sky130_fd_sc_hd__clkbuf_4
Xfanout177 _09153_/Y vssd1 vssd1 vccd1 vccd1 _10159_/A sky130_fd_sc_hd__clkbuf_8
Xfanout188 _12803_/B vssd1 vssd1 vccd1 vccd1 _13257_/A2 sky130_fd_sc_hd__clkbuf_8
X_09728_ _09394_/X _09404_/X _09728_/S vssd1 vssd1 vccd1 vccd1 _09728_/X sky130_fd_sc_hd__mux2_1
X_07989_ _07030_/Y _07097_/X _07256_/Y _07038_/X vssd1 vssd1 vccd1 vccd1 _07990_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout54_A _07072_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09659_ fanout57/X fanout86/X fanout82/X fanout63/X vssd1 vssd1 vccd1 vccd1 _09660_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12670_ reg1_val[6] _12670_/B vssd1 vssd1 vccd1 vccd1 _12671_/B sky130_fd_sc_hd__and2_1
X_11621_ _11430_/Y _11523_/Y _11525_/B vssd1 vssd1 vccd1 vccd1 _11621_/X sky130_fd_sc_hd__o21a_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09411__A _12644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11552_ _11552_/A _11552_/B vssd1 vssd1 vccd1 vccd1 _11552_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10276__B _10276_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11483_ fanout30/X _07608_/Y _08859_/Y fanout32/X vssd1 vssd1 vccd1 vccd1 _11484_/B
+ sky130_fd_sc_hd__a22o_1
X_10503_ _10503_/A _10503_/B vssd1 vssd1 vccd1 vccd1 _10504_/B sky130_fd_sc_hd__or2_1
X_13222_ hold278/A _13221_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13222_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_107_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10434_ hold215/A _10434_/B vssd1 vssd1 vccd1 vccd1 _10565_/B sky130_fd_sc_hd__or2_1
XFILLER_0_33_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13153_ _13153_/A _13153_/B vssd1 vssd1 vccd1 vccd1 _13154_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_100_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10365_ _11398_/A _10365_/B vssd1 vssd1 vccd1 vccd1 _10366_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_33_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12104_ _12105_/A _12105_/B vssd1 vssd1 vccd1 vccd1 _12177_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13126__B2 _06577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13084_ hold123/A _13094_/A2 _13250_/B hold108/X _13259_/A vssd1 vssd1 vccd1 vccd1
+ hold109/A sky130_fd_sc_hd__o221a_1
X_10296_ _10294_/X _10295_/X _11246_/S vssd1 vssd1 vccd1 vccd1 _10296_/X sky130_fd_sc_hd__mux2_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12035_ _12036_/A _12036_/B _12036_/C vssd1 vssd1 vccd1 vccd1 _12111_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_88_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12937_ _13168_/A _13169_/A _13168_/B vssd1 vssd1 vccd1 vccd1 _13174_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08856__A2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12868_ hold26/X _12870_/B vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__or2_1
XANTENNA__06841__A_N _07195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11819_ _11819_/A _11819_/B vssd1 vssd1 vccd1 vccd1 _11820_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_56_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06664__B _07147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12799_ hold66/X hold200/X hold298/X hold305/A vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__and4_1
XFILLER_0_7_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07010_ _09673_/A _07010_/B vssd1 vssd1 vccd1 vccd1 _07011_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11915__A2 _09257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11376__B1 _11752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08241__B1 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_14_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08961_ _10623_/A _08961_/B vssd1 vssd1 vccd1 vccd1 _08965_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07912_ _09302_/A _07912_/B vssd1 vssd1 vccd1 vccd1 _07913_/C sky130_fd_sc_hd__xnor2_1
X_08892_ _08893_/A _08893_/B _08893_/C vssd1 vssd1 vccd1 vccd1 _09022_/A sky130_fd_sc_hd__a21oi_1
X_07843_ _09834_/A _07936_/B _07936_/A vssd1 vssd1 vccd1 vccd1 _07863_/B sky130_fd_sc_hd__mux2_2
XANTENNA__10351__A1 _10479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07774_ _09670_/A _07774_/B vssd1 vssd1 vccd1 vccd1 _07777_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07016__A _07016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06725_ _06723_/Y _06724_/B1 _06783_/A reg2_val[16] vssd1 vssd1 vccd1 vccd1 _06727_/B
+ sky130_fd_sc_hd__a2bb2o_2
X_09513_ fanout28/X _11309_/A _11198_/A fanout25/X vssd1 vssd1 vccd1 vccd1 _09514_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08847__A2 _11093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06656_ _06654_/Y _06677_/B1 _06783_/A reg2_val[24] vssd1 vssd1 vccd1 vccd1 _06658_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_09444_ _10821_/A _09762_/B _09444_/C vssd1 vssd1 vccd1 vccd1 _09444_/X sky130_fd_sc_hd__or3_1
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06587_ pred_val instruction[1] vssd1 vssd1 vccd1 vccd1 _06911_/C sky130_fd_sc_hd__and2_1
XFILLER_0_93_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09375_ _09375_/A _09375_/B vssd1 vssd1 vccd1 vccd1 _09376_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_61_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08326_ _08689_/A _08689_/B vssd1 vssd1 vccd1 vccd1 _08326_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09272__A2 _12823_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08257_ _08564_/A _08257_/B vssd1 vssd1 vccd1 vccd1 _08317_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_104_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07208_ reg1_val[19] _07228_/B _07208_/C vssd1 vssd1 vccd1 vccd1 _07212_/B sky130_fd_sc_hd__or3_2
XANTENNA__12159__A2 _12158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07686__A _08580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08188_ _08188_/A _08188_/B vssd1 vssd1 vccd1 vccd1 _08275_/A sky130_fd_sc_hd__xor2_2
X_07139_ _09834_/A _07139_/B vssd1 vssd1 vccd1 vccd1 _07162_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13108__B2 _06577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10150_ _11630_/A _10151_/B _10151_/C vssd1 vssd1 vccd1 vccd1 _10152_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_30_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10840__A _12096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10081_ _11497_/A _10081_/B vssd1 vssd1 vccd1 vccd1 _10085_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__06749__B _06810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10983_ _10983_/A _10983_/B vssd1 vssd1 vccd1 vccd1 _10984_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__12095__A1 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12095__B2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11671__A _11671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12722_ _12722_/A _12722_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[15] sky130_fd_sc_hd__nor2_8
XFILLER_0_85_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07510__A2 _08289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13044__B1 _13254_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12653_ _12652_/A _12649_/Y _12651_/B vssd1 vssd1 vccd1 vccd1 _12657_/A sky130_fd_sc_hd__o21a_2
X_11604_ _11511_/A _11510_/B _11510_/A vssd1 vssd1 vccd1 vccd1 _11606_/B sky130_fd_sc_hd__o21ba_1
X_12584_ _12597_/B _12598_/B _12597_/A vssd1 vssd1 vccd1 vccd1 _12591_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_108_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11535_ _11893_/A _11472_/X _11567_/D _12356_/B1 vssd1 vssd1 vccd1 vccd1 _11536_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_25_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13205_ hold268/X _13223_/A2 _13204_/X _13223_/B2 vssd1 vssd1 vccd1 vccd1 hold269/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11358__B1 _12376_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11466_ hold246/A _11464_/X _11465_/Y vssd1 vssd1 vccd1 vccd1 _11466_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_80_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11397_ _06998_/X _07171_/A fanout38/X _07032_/Y vssd1 vssd1 vccd1 vccd1 _11398_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12007__A _12093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10417_ _10326_/X _10453_/B _12356_/B1 vssd1 vssd1 vccd1 vccd1 _10417_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07577__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10348_ _10748_/A _10348_/B vssd1 vssd1 vccd1 vccd1 _10353_/A sky130_fd_sc_hd__xnor2_2
X_13136_ hold281/X _13254_/A2 _13135_/X _06577_/A vssd1 vssd1 vccd1 vccd1 _13137_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06785__B1 _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11846__A _12096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13067_ _07267_/B _12826_/B hold153/X vssd1 vssd1 vccd1 vccd1 _13343_/D sky130_fd_sc_hd__a21boi_1
X_10279_ _09999_/A _09999_/B _10136_/A _10136_/B vssd1 vssd1 vccd1 vccd1 _10279_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12018_ fanout41/X _07608_/Y _08859_/Y fanout43/X vssd1 vssd1 vccd1 vccd1 _12019_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11581__A _11582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07490_ _07490_/A _07490_/B _07489_/X vssd1 vssd1 vccd1 vccd1 _07533_/A sky130_fd_sc_hd__or3b_1
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09160_ _09156_/X _09159_/X _09725_/S vssd1 vssd1 vccd1 vccd1 _09160_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11061__A2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09091_ _09298_/A1 fanout14/X fanout13/X _09298_/B2 vssd1 vssd1 vccd1 vccd1 _09092_/B
+ sky130_fd_sc_hd__o22a_1
X_08111_ _08110_/A _08157_/A _08116_/A vssd1 vssd1 vccd1 vccd1 _08111_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_126_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08042_ _09670_/A _08042_/B vssd1 vssd1 vccd1 vccd1 _08046_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07017__A1 _07016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout104_A _09479_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09993_ _09993_/A _09993_/B vssd1 vssd1 vccd1 vccd1 _09995_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08944_ _08844_/A _08843_/Y _08839_/Y vssd1 vssd1 vccd1 vccd1 _08946_/B sky130_fd_sc_hd__a21oi_2
X_08875_ _08876_/A _08876_/B vssd1 vssd1 vccd1 vccd1 _08875_/X sky130_fd_sc_hd__and2_1
X_07826_ _07826_/A _07826_/B vssd1 vssd1 vccd1 vccd1 _07935_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07757_ _07866_/A _07866_/B _07753_/Y vssd1 vssd1 vccd1 vccd1 _07802_/A sky130_fd_sc_hd__o21ai_1
X_06708_ _06708_/A vssd1 vssd1 vccd1 vccd1 _11636_/A sky130_fd_sc_hd__inv_2
XFILLER_0_94_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07688_ _07688_/A _07688_/B vssd1 vssd1 vccd1 vccd1 _07752_/A sky130_fd_sc_hd__xor2_2
XANTENNA__13026__B1 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06639_ _12438_/B _06639_/B vssd1 vssd1 vccd1 vccd1 _12406_/A sky130_fd_sc_hd__or2_2
X_09427_ _09586_/A _11554_/A _09414_/X _11820_/A vssd1 vssd1 vccd1 vccd1 _09427_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_47_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09358_ _09112_/A _09112_/B _09110_/Y vssd1 vssd1 vccd1 vccd1 _09361_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11588__B1 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout17_A _12286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08309_ _08352_/B _08352_/A vssd1 vssd1 vccd1 vccd1 _08309_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__08453__B1 _09479_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11320_ _11320_/A _11320_/B vssd1 vssd1 vccd1 vccd1 _11322_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_105_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09289_ fanout57/X _10473_/B2 _10240_/A fanout63/X vssd1 vssd1 vccd1 vccd1 _09290_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_105_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08305__A _08580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11251_ hold193/A _11251_/B vssd1 vssd1 vccd1 vccd1 _11363_/B sky130_fd_sc_hd__or2_1
X_11182_ _11182_/A _11182_/B vssd1 vssd1 vccd1 vccd1 _11183_/B sky130_fd_sc_hd__xnor2_2
X_10202_ _10203_/B _10203_/A vssd1 vssd1 vccd1 vccd1 _10202_/X sky130_fd_sc_hd__and2b_1
X_10133_ _10134_/A _10134_/B vssd1 vssd1 vccd1 vccd1 _10133_/X sky130_fd_sc_hd__and2_1
X_10064_ _10065_/A _10065_/B vssd1 vssd1 vccd1 vccd1 _10064_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10315__A1 _12379_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08040__A _08664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10966_ _10966_/A _10966_/B vssd1 vssd1 vccd1 vccd1 _10967_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_85_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10897_ _10897_/A _10897_/B _10897_/C vssd1 vssd1 vccd1 vccd1 _10898_/B sky130_fd_sc_hd__and3_1
XFILLER_0_85_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12705_ _12705_/A _12705_/B _12705_/C vssd1 vssd1 vccd1 vccd1 _12706_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_122_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12636_ _12636_/A _12636_/B vssd1 vssd1 vccd1 vccd1 new_PC[26] sky130_fd_sc_hd__xnor2_4
XFILLER_0_72_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11579__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06942__B _06944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12567_ _12567_/A _12567_/B _12567_/C vssd1 vssd1 vccd1 vccd1 _12568_/B sky130_fd_sc_hd__nand3_1
XANTENNA__10745__A _10950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11518_ _11518_/A _11518_/B vssd1 vssd1 vccd1 vccd1 _11519_/B sky130_fd_sc_hd__or2_1
X_12498_ _12504_/B _12498_/B vssd1 vssd1 vccd1 vccd1 new_PC[5] sky130_fd_sc_hd__and2_4
XFILLER_0_80_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold208 hold208/A vssd1 vssd1 vccd1 vccd1 hold208/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold219 hold219/A vssd1 vssd1 vccd1 vccd1 hold219/X sky130_fd_sc_hd__dlygate4sd3_1
X_11449_ _11449_/A _11449_/B vssd1 vssd1 vccd1 vccd1 _11449_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11576__A _12096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13119_ _13147_/A hold257/X vssd1 vssd1 vccd1 vccd1 _13364_/D sky130_fd_sc_hd__and2_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06990_ _07046_/B _06991_/B vssd1 vssd1 vccd1 vccd1 _12169_/A sky130_fd_sc_hd__xor2_4
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08660_ _08659_/B _08661_/A vssd1 vssd1 vccd1 vccd1 _08660_/X sky130_fd_sc_hd__and2b_1
X_07611_ fanout65/X _09669_/B2 _09301_/A fanout59/X vssd1 vssd1 vccd1 vccd1 _07612_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08591_ _08592_/A _08592_/B vssd1 vssd1 vccd1 vccd1 _08733_/A sky130_fd_sc_hd__or2_1
XFILLER_0_48_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07542_ _11381_/A _07542_/B vssd1 vssd1 vccd1 vccd1 _07546_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__13008__B1 _13209_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07473_ _09836_/A _07473_/B vssd1 vssd1 vccd1 vccd1 _07475_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10490__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09212_ _09210_/X _09211_/X _09403_/S vssd1 vssd1 vccd1 vccd1 _09212_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_127_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12854__B _12862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09143_ _09143_/A _09143_/B vssd1 vssd1 vccd1 vccd1 _09144_/B sky130_fd_sc_hd__xor2_4
XANTENNA__13031__A _13162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08986__A1 _12404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_551 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09074_ _09075_/A _09075_/B vssd1 vssd1 vccd1 vccd1 _09074_/Y sky130_fd_sc_hd__nor2_1
Xfanout2 fanout2/A vssd1 vssd1 vccd1 vccd1 fanout2/X sky130_fd_sc_hd__buf_6
X_08025_ _08095_/A _08025_/B vssd1 vssd1 vccd1 vccd1 _08027_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_114_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09935__B1 _07238_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07964__A _09341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10545__A1 _10415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09976_ _09976_/A _09976_/B vssd1 vssd1 vccd1 vccd1 _09979_/A sky130_fd_sc_hd__xnor2_2
X_08927_ _08943_/B _08855_/B _08868_/B _08869_/B _08869_/A vssd1 vssd1 vccd1 vccd1
+ _08940_/B sky130_fd_sc_hd__a32o_1
X_08858_ _06866_/B _06867_/B _07315_/A _07094_/B vssd1 vssd1 vccd1 vccd1 _08860_/B
+ sky130_fd_sc_hd__a31o_2
X_07809_ _07807_/A _07807_/B _07879_/A vssd1 vssd1 vccd1 vccd1 _07820_/A sky130_fd_sc_hd__o21ba_1
X_08789_ _08076_/A _08076_/B _08788_/X vssd1 vssd1 vccd1 vccd1 _08793_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10820_ curr_PC[11] _10934_/C vssd1 vssd1 vccd1 vccd1 _10821_/B sky130_fd_sc_hd__and2_1
XFILLER_0_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10751_ _10751_/A _10751_/B vssd1 vssd1 vccd1 vccd1 _10752_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_67_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07204__A _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12421_ _12421_/A1 _12420_/X _06639_/B vssd1 vssd1 vccd1 vccd1 _12422_/B sky130_fd_sc_hd__a21oi_1
X_10682_ _10015_/Y _10681_/Y _11029_/S vssd1 vssd1 vccd1 vccd1 _10682_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12352_ _12246_/X _12350_/B _12350_/Y _12117_/Y vssd1 vssd1 vccd1 vccd1 _12352_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_90_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08035__A _10207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11303_ _11303_/A _11303_/B vssd1 vssd1 vccd1 vccd1 _11304_/B sky130_fd_sc_hd__or2_1
XANTENNA__11981__B1 _09225_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12283_ _12284_/A _12284_/B _12284_/C vssd1 vssd1 vccd1 vccd1 _12285_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11234_ _11234_/A _11271_/B vssd1 vssd1 vccd1 vccd1 _11234_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11165_ _12087_/B _11165_/B vssd1 vssd1 vccd1 vccd1 _11169_/B sky130_fd_sc_hd__xnor2_1
X_11096_ _11096_/A _11096_/B vssd1 vssd1 vccd1 vccd1 _11098_/B sky130_fd_sc_hd__xor2_1
XANTENNA__12289__A1 _12157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10116_ _10116_/A _10116_/B vssd1 vssd1 vccd1 vccd1 _10118_/A sky130_fd_sc_hd__xor2_4
XANTENNA__10839__A2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10047_ _10821_/A _10043_/X _10044_/X _10046_/Y vssd1 vssd1 vccd1 vccd1 dest_val[5]
+ sky130_fd_sc_hd__a22o_4
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06912__B1 _12218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11998_ _10159_/A _10432_/Y _10444_/Y _09222_/Y _11997_/X vssd1 vssd1 vccd1 vccd1
+ _11998_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_128_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10949_ _11182_/A _10949_/B vssd1 vssd1 vccd1 vccd1 _10950_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12674__B _12675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12619_ reg1_val[24] curr_PC[24] _12638_/S vssd1 vssd1 vccd1 vccd1 _12620_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_54_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11016__A2 _11050_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08417__B1 _08501_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09830_ _09830_/A _09830_/B vssd1 vssd1 vccd1 vccd1 _09831_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_6_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06973_ _07133_/A _06974_/B vssd1 vssd1 vccd1 vccd1 _06983_/A sky130_fd_sc_hd__nor2_4
X_09761_ curr_PC[3] _09762_/B vssd1 vssd1 vccd1 vccd1 _09761_/X sky130_fd_sc_hd__or2_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08712_ _12129_/B vssd1 vssd1 vccd1 vccd1 _08712_/Y sky130_fd_sc_hd__inv_2
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09692_ _09461_/A _09461_/B _09464_/A vssd1 vssd1 vccd1 vccd1 _09697_/A sky130_fd_sc_hd__o21ai_4
XANTENNA_fanout171_A _12805_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06847__B _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08643_ _08637_/A _08637_/C _08637_/B vssd1 vssd1 vccd1 vccd1 _08646_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08574_ _07030_/Y _07134_/Y _07166_/Y _07038_/X vssd1 vssd1 vccd1 vccd1 _08575_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09448__A2 _07362_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07459__A1 _09943_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07459__B2 _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07525_ _09944_/A _07525_/B vssd1 vssd1 vccd1 vccd1 _07721_/A sky130_fd_sc_hd__xnor2_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07959__A _07959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07456_ _09669_/B2 fanout61/X fanout53/X _09301_/A vssd1 vssd1 vccd1 vccd1 _07457_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12204__A1 _12447_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10385__A _11182_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07387_ _07387_/A _07387_/B vssd1 vssd1 vccd1 vccd1 _07388_/B sky130_fd_sc_hd__and2_1
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09126_ _09126_/A _09126_/B vssd1 vssd1 vccd1 vccd1 _09128_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07631__A1 _07830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09057_ _09056_/B _09057_/B vssd1 vssd1 vccd1 vccd1 _09058_/B sky130_fd_sc_hd__and2b_1
XANTENNA__07631__B2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08008_ _08009_/A _08009_/B vssd1 vssd1 vccd1 vccd1 _08008_/X sky130_fd_sc_hd__and2_1
XANTENNA__11191__A1 _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11191__B2 _12009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ _09959_/A _09959_/B vssd1 vssd1 vccd1 vccd1 _09960_/B sky130_fd_sc_hd__xor2_4
XANTENNA_fanout84_A _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12970_ _12874_/B _13243_/B _12874_/A vssd1 vssd1 vccd1 vccd1 _12971_/B sky130_fd_sc_hd__o21ba_1
XANTENNA__11494__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11921_ curr_PC[22] _12003_/C vssd1 vssd1 vccd1 vccd1 _11921_/X sky130_fd_sc_hd__or2_1
XANTENNA__06757__B _07233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11852_ fanout38/X _07608_/Y _08859_/Y _07171_/A vssd1 vssd1 vccd1 vccd1 _11853_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09439__A2 _12412_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10803_ _09879_/Y _10802_/Y _11029_/S vssd1 vssd1 vccd1 vccd1 _10803_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08647__B1 _07173_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11783_ _11783_/A _11783_/B vssd1 vssd1 vccd1 vccd1 _11785_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_95_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10734_ _10734_/A _10734_/B vssd1 vssd1 vccd1 vccd1 _10737_/A sky130_fd_sc_hd__xor2_1
XANTENNA__12994__A2 _13000_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10665_ _11809_/A _11271_/A _11050_/A vssd1 vssd1 vccd1 vccd1 _10665_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07588__B _11844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13384_ _13385_/CLK _13384_/D vssd1 vssd1 vccd1 vccd1 hold254/A sky130_fd_sc_hd__dfxtp_1
X_12404_ _06887_/X _12406_/B _12404_/S vssd1 vssd1 vccd1 vccd1 _12404_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10206__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13102__C fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09072__B1 _10240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10596_ _12087_/B _10596_/B vssd1 vssd1 vccd1 vccd1 _10597_/B sky130_fd_sc_hd__xnor2_2
X_12335_ _12335_/A _12335_/B vssd1 vssd1 vccd1 vccd1 _12336_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_51_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12266_ hold229/A _12266_/B vssd1 vssd1 vccd1 vccd1 _12321_/B sky130_fd_sc_hd__or2_1
X_11217_ _11217_/A _11217_/B vssd1 vssd1 vccd1 vccd1 _11219_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13171__A2 _13223_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12015__A _12336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12197_ _12192_/X _12195_/X _12196_/Y vssd1 vssd1 vccd1 vccd1 _12197_/X sky130_fd_sc_hd__a21o_1
X_11148_ _11646_/B _11251_/B hold193/A vssd1 vssd1 vccd1 vccd1 _11148_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07925__A2 _10595_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11079_ _11182_/A _11079_/B vssd1 vssd1 vccd1 vccd1 _11084_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12669__B _12670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07138__B1 _09822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07689__A1 _08540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07689__B2 _08515_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07310_ _07310_/A _07310_/B vssd1 vssd1 vccd1 vccd1 _07368_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08290_ _08334_/A _08290_/B vssd1 vssd1 vccd1 vccd1 _08350_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__07779__A _08575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07241_ _07241_/A _07241_/B vssd1 vssd1 vccd1 vccd1 _07242_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_27_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07172_ _07172_/A _07173_/B vssd1 vssd1 vccd1 vccd1 _07172_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09813_ _09944_/A _09813_/B vssd1 vssd1 vccd1 vccd1 _09817_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07019__A _07020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11764__A _11764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06956_ _06958_/A _06956_/B vssd1 vssd1 vccd1 vccd1 dest_mask[0] sky130_fd_sc_hd__nand2_8
X_09744_ _12054_/S _06822_/X _09743_/X vssd1 vssd1 vccd1 vccd1 _09746_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__09669__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06887_ _06625_/Y _12359_/B _06877_/A vssd1 vssd1 vccd1 vccd1 _06887_/X sky130_fd_sc_hd__a21bo_1
X_09675_ _09675_/A _09675_/B vssd1 vssd1 vccd1 vccd1 _09676_/B sky130_fd_sc_hd__xor2_2
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08626_ _08618_/A _08618_/B _08618_/C vssd1 vssd1 vccd1 vccd1 _08630_/B sky130_fd_sc_hd__a21oi_2
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13190__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08557_ _08557_/A _08557_/B vssd1 vssd1 vccd1 vccd1 _08564_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_119_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10436__B1 _12205_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12976__A2 _13000_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08488_ _08498_/A _08498_/B _08482_/Y vssd1 vssd1 vccd1 vccd1 _08496_/B sky130_fd_sc_hd__a21bo_1
X_07508_ fanout76/X _08484_/B _09479_/B1 fanout72/X vssd1 vssd1 vccd1 vccd1 _07509_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_91_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07439_ _07562_/A vssd1 vssd1 vccd1 vccd1 _07439_/Y sky130_fd_sc_hd__inv_2
X_10450_ _10821_/A _10699_/C _10450_/C vssd1 vssd1 vccd1 vccd1 _10450_/X sky130_fd_sc_hd__or3_1
XANTENNA__09054__B1 _07282_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09109_ _09109_/A _09109_/B vssd1 vssd1 vccd1 vccd1 _09111_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12534__S _12638_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10381_ _10381_/A _10381_/B vssd1 vssd1 vccd1 vccd1 _10382_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_32_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12120_ _12300_/B _12120_/B vssd1 vssd1 vccd1 vccd1 _12184_/B sky130_fd_sc_hd__xor2_2
X_12051_ _11892_/A _12050_/X _12184_/A vssd1 vssd1 vccd1 vccd1 _12051_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11164__B2 _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11164__A1 _11406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11002_ _10888_/A _10888_/B _10889_/Y vssd1 vssd1 vccd1 vccd1 _11004_/B sky130_fd_sc_hd__o21a_1
XANTENNA__12361__B1 _09225_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12953_ _12884_/X _12953_/B vssd1 vssd1 vccd1 vccd1 _13207_/B sky130_fd_sc_hd__nand2b_1
X_11904_ _11819_/A _11819_/B _11817_/A vssd1 vssd1 vccd1 vccd1 _11905_/B sky130_fd_sc_hd__o21a_1
XANTENNA__08332__A2 _08561_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12884_ hold62/X hold268/A vssd1 vssd1 vccd1 vccd1 _12884_/X sky130_fd_sc_hd__and2b_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ _11807_/Y _11808_/X _11810_/X _10788_/A _11834_/X vssd1 vssd1 vccd1 vccd1
+ _11835_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_23_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _11766_/A _11766_/B vssd1 vssd1 vccd1 vccd1 _11767_/B sky130_fd_sc_hd__or2_1
XFILLER_0_95_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11840__C _11840_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09293__B1 _10245_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10717_ _12093_/A _10717_/B vssd1 vssd1 vccd1 vccd1 _10719_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_83_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11697_ _11698_/A _11698_/B _11698_/C vssd1 vssd1 vccd1 vccd1 _11793_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10648_ _10649_/B _10649_/A vssd1 vssd1 vccd1 vccd1 _10648_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_23_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13367_ _13369_/CLK _13367_/D vssd1 vssd1 vccd1 vccd1 hold260/A sky130_fd_sc_hd__dfxtp_1
X_10579_ _12356_/B1 _10549_/Y _10550_/X _10578_/X vssd1 vssd1 vccd1 vccd1 _10579_/X
+ sky130_fd_sc_hd__a31o_1
X_12318_ reg1_val[28] _12366_/C vssd1 vssd1 vccd1 vccd1 _12318_/X sky130_fd_sc_hd__xor2_1
X_13298_ _13304_/CLK _13298_/D vssd1 vssd1 vccd1 vccd1 hold301/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12249_ _12430_/A _12249_/B vssd1 vssd1 vccd1 vccd1 _12306_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08020__A1 _08540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08020__B2 _08515_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08877__B _08877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11584__A _11584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06810_ reg2_val[1] _06810_/B vssd1 vssd1 vccd1 vccd1 _06810_/X sky130_fd_sc_hd__and2_2
X_07790_ _07790_/A _07790_/B vssd1 vssd1 vccd1 vccd1 _07826_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11458__A2 _09257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06741_ reg1_val[13] _11038_/A vssd1 vssd1 vccd1 vccd1 _11039_/S sky130_fd_sc_hd__and2_1
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09520__B2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09520__A1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10666__B1 _09150_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09460_ _09284_/A _09284_/B _09285_/X vssd1 vssd1 vccd1 vccd1 _09461_/B sky130_fd_sc_hd__a21oi_2
X_06672_ _06672_/A _06672_/B _06962_/B _06672_/D vssd1 vssd1 vccd1 vccd1 _06672_/X
+ sky130_fd_sc_hd__and4_1
X_08411_ _09404_/S _08411_/B vssd1 vssd1 vccd1 vccd1 _08449_/B sky130_fd_sc_hd__nor2_1
XANTENNA__12619__S _12638_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09391_ _09389_/X _09390_/X _09727_/S vssd1 vssd1 vccd1 vccd1 _10018_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_46_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08342_ _08342_/A _08342_/B vssd1 vssd1 vccd1 vccd1 _08393_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11091__B1 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10969__B2 _11093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10969__A1 _11198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08273_ _08284_/A _08284_/B _08262_/Y vssd1 vssd1 vccd1 vccd1 _08282_/B sky130_fd_sc_hd__a21o_1
XANTENNA_fanout134_A _07092_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07224_ _09836_/A _07224_/B vssd1 vssd1 vccd1 vccd1 _07226_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12862__B _12862_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11759__A _12096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07155_ _07155_/A _07155_/B _07155_/C vssd1 vssd1 vccd1 vccd1 _07158_/B sky130_fd_sc_hd__and3_1
XFILLER_0_42_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07086_ reg1_val[9] _07086_/B vssd1 vssd1 vccd1 vccd1 _07086_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_112_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout101 _07088_/Y vssd1 vssd1 vccd1 vccd1 _11476_/A sky130_fd_sc_hd__buf_4
XFILLER_0_100_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout112 _07233_/Y vssd1 vssd1 vccd1 vccd1 _10599_/A sky130_fd_sc_hd__buf_4
XANTENNA__13185__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout123 _07187_/Y vssd1 vssd1 vccd1 vccd1 _08334_/A sky130_fd_sc_hd__buf_12
Xfanout134 _07092_/Y vssd1 vssd1 vccd1 vccd1 _10245_/B2 sky130_fd_sc_hd__buf_8
Xfanout156 _07011_/Y vssd1 vssd1 vccd1 vccd1 _09669_/B2 sky130_fd_sc_hd__buf_8
Xfanout145 _09650_/A vssd1 vssd1 vccd1 vccd1 _08538_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout167 _06962_/Y vssd1 vssd1 vccd1 vccd1 _12322_/A1 sky130_fd_sc_hd__buf_4
Xfanout189 _13248_/B1 vssd1 vssd1 vccd1 vccd1 _13209_/A2 sky130_fd_sc_hd__buf_4
Xfanout178 _12379_/B2 vssd1 vssd1 vccd1 vccd1 _09180_/S sky130_fd_sc_hd__clkbuf_8
X_07988_ _07988_/A _07988_/B _07988_/C vssd1 vssd1 vccd1 vccd1 _08065_/A sky130_fd_sc_hd__or3_2
X_06939_ instruction[20] _06590_/X _06938_/X _06716_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[2]
+ sky130_fd_sc_hd__o211a_4
X_09727_ _09401_/X _09403_/X _09727_/S vssd1 vssd1 vccd1 vccd1 _09727_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_96_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10657__B1 _10539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout47_A _07830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09658_ _09658_/A _09658_/B vssd1 vssd1 vccd1 vccd1 _09676_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _06809_/Y _09587_/X _09588_/Y vssd1 vssd1 vccd1 vccd1 _09589_/Y sky130_fd_sc_hd__o21ai_1
X_08609_ _08609_/A _08609_/B vssd1 vssd1 vccd1 vccd1 _08610_/B sky130_fd_sc_hd__or2_1
X_11620_ _11968_/A vssd1 vssd1 vccd1 vccd1 _11620_/Y sky130_fd_sc_hd__inv_2
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11551_ hold264/A _11650_/B _11649_/B _12376_/C1 vssd1 vssd1 vccd1 vccd1 _11552_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09814__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08308__A _08564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10502_ _10501_/A _10501_/B _10501_/C vssd1 vssd1 vccd1 vccd1 _10503_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11482_ _12093_/A _11482_/B vssd1 vssd1 vccd1 vccd1 _11486_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11909__B1 _11648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13221_ _13221_/A _13221_/B vssd1 vssd1 vccd1 vccd1 _13221_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10433_ _10429_/Y _10432_/Y _11820_/A vssd1 vssd1 vccd1 vccd1 _10433_/X sky130_fd_sc_hd__mux2_1
X_13152_ _13246_/A hold280/X vssd1 vssd1 vccd1 vccd1 _13371_/D sky130_fd_sc_hd__and2_1
XANTENNA__11924__A3 _12049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10364_ _07171_/A _07256_/Y _07262_/X fanout38/X vssd1 vssd1 vccd1 vccd1 _10365_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12103_ _12103_/A _12103_/B vssd1 vssd1 vccd1 vccd1 _12105_/B sky130_fd_sc_hd__xor2_1
XANTENNA__13126__A2 _13254_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13083_ _07128_/Y _13089_/A2 hold124/X vssd1 vssd1 vccd1 vccd1 _13351_/D sky130_fd_sc_hd__o21a_1
X_10295_ _09722_/X _09727_/X _10295_/S vssd1 vssd1 vccd1 vccd1 _10295_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09573__S _09728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12034_ _12111_/A _12034_/B vssd1 vssd1 vccd1 vccd1 _12036_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_18_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12936_ hold50/X hold270/X vssd1 vssd1 vccd1 vccd1 _13168_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_88_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07513__B1 _10476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12867_ _07608_/Y _12871_/A2 hold29/X _13246_/A vssd1 vssd1 vccd1 vccd1 _13294_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10748__A _10748_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11818_ _11732_/A _11732_/B _11730_/A vssd1 vssd1 vccd1 vccd1 _11819_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_55_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11073__B1 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12798_ hold127/X hold167/X hold140/X vssd1 vssd1 vccd1 vccd1 _12798_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_7_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11749_ curr_PC[19] curr_PC[20] _11749_/C vssd1 vssd1 vccd1 vccd1 _11837_/B sky130_fd_sc_hd__and3_1
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06961__A _11813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08241__A1 _06992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09049__A _09936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08241__B2 _08613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08960_ fanout51/X fanout86/X fanout82/X _09661_/B2 vssd1 vssd1 vccd1 vccd1 _08961_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08888__A _09836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07911_ _09669_/B2 fanout84/X fanout80/X _09301_/A vssd1 vssd1 vccd1 vccd1 _07912_/B
+ sky130_fd_sc_hd__o22a_1
X_08891_ _08946_/A _08891_/B vssd1 vssd1 vccd1 vccd1 _08893_/C sky130_fd_sc_hd__or2_1
XANTENNA__07792__A _09667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10422__S _12054_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07842_ _07842_/A _07885_/A vssd1 vssd1 vccd1 vccd1 _07936_/B sky130_fd_sc_hd__nand2_1
X_07773_ _08641_/B _09661_/B2 fanout98/X _08627_/A2 vssd1 vssd1 vccd1 vccd1 _07774_/B
+ sky130_fd_sc_hd__o22a_1
X_09512_ _09512_/A _09512_/B vssd1 vssd1 vccd1 vccd1 _09527_/A sky130_fd_sc_hd__nor2_1
X_06724_ reg2_val[16] _06783_/A _06724_/B1 _06723_/Y vssd1 vssd1 vccd1 vccd1 _07094_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_79_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06655_ reg2_val[24] _06783_/A _06677_/B1 _06654_/Y vssd1 vssd1 vccd1 vccd1 _06995_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_91_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout251_A _06723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09443_ curr_PC[0] curr_PC[1] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _09444_/C sky130_fd_sc_hd__a21oi_1
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06855__B _07078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09257__A0 _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13053__A1 _10243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09374_ _09708_/A _09035_/X _09863_/A _09711_/C _09711_/A vssd1 vssd1 vccd1 vccd1
+ _09375_/B sky130_fd_sc_hd__o32a_2
X_06586_ instruction[0] pred_val vssd1 vssd1 vccd1 vccd1 _06911_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_46_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08325_ _08689_/A _08689_/B vssd1 vssd1 vccd1 vccd1 _08325_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_19_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08256_ _08540_/B _09770_/B2 _09940_/B2 _08515_/A2 vssd1 vssd1 vccd1 vccd1 _08257_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11489__A _11929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07207_ _07228_/B _07208_/C reg1_val[19] vssd1 vssd1 vccd1 vccd1 _07212_/A sky130_fd_sc_hd__o21ai_2
X_08187_ _08188_/A _08188_/B vssd1 vssd1 vccd1 vccd1 _08187_/X sky130_fd_sc_hd__and2_1
XANTENNA__11367__A1 _10159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07138_ _08561_/A2 _07830_/B _09822_/A fanout46/X vssd1 vssd1 vccd1 vccd1 _07139_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13108__A2 _13254_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07069_ _07094_/B _06987_/A _07016_/A vssd1 vssd1 vccd1 vccd1 _07907_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__12316__B1 _12365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12867__A1 _07608_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10080_ _10337_/A _08875_/X _08990_/Y _10225_/A vssd1 vssd1 vccd1 vccd1 _10081_/B
+ sky130_fd_sc_hd__a22o_1
X_10982_ _10983_/B _10983_/A vssd1 vssd1 vccd1 vccd1 _11102_/B sky130_fd_sc_hd__and2b_1
XANTENNA__12095__A2 _08859_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09496__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11671__B _11946_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09422__A _09728_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12721_ _12721_/A _12721_/B _12721_/C vssd1 vssd1 vccd1 vccd1 _12722_/B sky130_fd_sc_hd__and3_2
X_12652_ _12652_/A _12652_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[2] sky130_fd_sc_hd__xnor2_4
XFILLER_0_127_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11603_ _11603_/A _11603_/B vssd1 vssd1 vccd1 vccd1 _11606_/A sky130_fd_sc_hd__xor2_1
X_12583_ _12570_/B _12575_/B _12639_/A vssd1 vssd1 vccd1 vccd1 _12598_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_53_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11534_ _11893_/A _11472_/X _11567_/D vssd1 vssd1 vccd1 vccd1 _11536_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11465_ hold246/A _11464_/X _09238_/Y vssd1 vssd1 vccd1 vccd1 _11465_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_53_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13204_ hold274/A _13203_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13204_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12555__A0 _11134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10416_ _10416_/A _10661_/C vssd1 vssd1 vccd1 vccd1 _10453_/B sky130_fd_sc_hd__xor2_4
X_11396_ _11396_/A _11396_/B vssd1 vssd1 vccd1 vccd1 _11399_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_96_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12007__B fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09420__B1 _11637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12307__B1 _11892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10347_ _07299_/X fanout14/X fanout13/X _10473_/B2 vssd1 vssd1 vccd1 vccd1 _10348_/B
+ sky130_fd_sc_hd__o22a_1
X_13135_ hold260/X _13134_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13135_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ hold130/X _13094_/A2 _13101_/A2 hold135/X _13039_/A vssd1 vssd1 vccd1 vccd1
+ hold153/A sky130_fd_sc_hd__o221a_1
XANTENNA__07982__B1 _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10278_ _10278_/A _10541_/A vssd1 vssd1 vccd1 vccd1 _10278_/Y sky130_fd_sc_hd__nand2_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12017_ _12017_/A _12017_/B vssd1 vssd1 vccd1 vccd1 _12021_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13119__A _13147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07117__A _12438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06956__A _06958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12919_ _12904_/B _13124_/B _12902_/X vssd1 vssd1 vccd1 vccd1 _13129_/A sky130_fd_sc_hd__a21o_1
XANTENNA__06675__B _06675_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10478__A _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08110_ _08110_/A _08157_/A vssd1 vssd1 vccd1 vccd1 _08116_/B sky130_fd_sc_hd__nor2_1
X_09090_ _09281_/B _09090_/B vssd1 vssd1 vccd1 vccd1 _09101_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08041_ _08641_/B fanout76/X fanout72/X _08627_/A2 vssd1 vssd1 vccd1 vccd1 _08042_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10941__A _12093_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09992_ _09992_/A _09992_/B vssd1 vssd1 vccd1 vccd1 _09993_/B sky130_fd_sc_hd__xor2_2
XANTENNA__12849__A1 _11764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10572__A2 _09257_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08943_ _08849_/X _08943_/B vssd1 vssd1 vccd1 vccd1 _08948_/A sky130_fd_sc_hd__and2b_1
XANTENNA__13029__A _13162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08411__A _09404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08874_ _12336_/A _08874_/B vssd1 vssd1 vccd1 vccd1 _08876_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07725__B1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07027__A _09672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07825_ _07828_/A _07828_/B vssd1 vssd1 vccd1 vccd1 _07825_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11772__A _11929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07756_ _07866_/A _07866_/B vssd1 vssd1 vccd1 vccd1 _07756_/X sky130_fd_sc_hd__or2_1
X_06707_ _11652_/S _06707_/B vssd1 vssd1 vccd1 vccd1 _06708_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_79_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09242__A _12795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11285__B1 _10092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09426_ _12416_/C1 _09424_/Y _09425_/X _09257_/S _09728_/S vssd1 vssd1 vccd1 vccd1
+ _09426_/X sky130_fd_sc_hd__o32a_1
X_07687_ _07688_/A _07688_/B vssd1 vssd1 vccd1 vccd1 _07687_/Y sky130_fd_sc_hd__nor2_1
X_06638_ reg1_val[30] _08973_/C vssd1 vssd1 vccd1 vccd1 _06639_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_59_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11588__A1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11037__B1 _12376_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09357_ _09357_/A _09357_/B vssd1 vssd1 vccd1 vccd1 _09362_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_19_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11588__B2 _11671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08308_ _08564_/A _08308_/B vssd1 vssd1 vccd1 vccd1 _08352_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07697__A _09947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08453__A1 _08649_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09288_ _09944_/A _09288_/B vssd1 vssd1 vccd1 vccd1 _09292_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08239_ _08334_/A _08239_/B vssd1 vssd1 vccd1 vccd1 _08314_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08453__B2 _09404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11250_ _11820_/A _11245_/Y _11249_/Y _06946_/X vssd1 vssd1 vccd1 vccd1 _11265_/B
+ sky130_fd_sc_hd__o211a_1
X_11181_ fanout34/X fanout12/X fanout7/X fanout36/X vssd1 vssd1 vccd1 vccd1 _11182_/B
+ sky130_fd_sc_hd__o22a_1
X_10201_ _10201_/A _10201_/B vssd1 vssd1 vccd1 vccd1 _10203_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10132_ _10132_/A _10132_/B vssd1 vssd1 vccd1 vccd1 _10134_/B sky130_fd_sc_hd__xnor2_2
X_10063_ _10065_/A _10065_/B vssd1 vssd1 vccd1 vccd1 _10063_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11276__B1 _07316_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09152__A _12054_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10965_ _11770_/A _10965_/B vssd1 vssd1 vccd1 vccd1 _10966_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12704_ _12705_/A _12705_/B _12705_/C vssd1 vssd1 vccd1 vccd1 _12711_/B sky130_fd_sc_hd__a21o_1
X_10896_ _10897_/A _10897_/B _10897_/C vssd1 vssd1 vccd1 vccd1 _10896_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_57_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12635_ _12628_/B _12630_/B _12628_/A vssd1 vssd1 vccd1 vccd1 _12636_/B sky130_fd_sc_hd__o21ba_2
XFILLER_0_72_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11579__B2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11579__A1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12566_ _12567_/A _12567_/B _12567_/C vssd1 vssd1 vccd1 vccd1 _12572_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_38_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11517_ _11518_/A _11518_/B vssd1 vssd1 vccd1 vccd1 _11616_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12497_ _12497_/A _12497_/B _12497_/C vssd1 vssd1 vccd1 vccd1 _12498_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_80_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11448_ _11813_/S _06850_/Y _11447_/Y vssd1 vssd1 vccd1 vccd1 _11449_/B sky130_fd_sc_hd__o21ai_1
Xhold209 hold209/A vssd1 vssd1 vccd1 vccd1 hold209/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11379_ _11770_/A _11379_/B vssd1 vssd1 vccd1 vccd1 _11381_/B sky130_fd_sc_hd__xnor2_1
X_13118_ hold256/X _13254_/A2 _13117_/X _06577_/A vssd1 vssd1 vccd1 vccd1 hold257/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09327__A _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ hold1/X _13101_/A2 _09302_/A _13101_/B2 _13048_/Y vssd1 vssd1 vccd1 vccd1
+ hold2/A sky130_fd_sc_hd__o221a_1
XFILLER_0_56_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11592__A _11592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07610_ _09671_/A _07610_/B vssd1 vssd1 vccd1 vccd1 _07614_/A sky130_fd_sc_hd__xnor2_4
X_08590_ _08568_/A _08568_/B _08568_/C vssd1 vssd1 vccd1 vccd1 _08739_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_72_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07541_ _07191_/X _10337_/A _12823_/A1 _07202_/Y vssd1 vssd1 vccd1 vccd1 _07542_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07472_ _07121_/Y _07959_/B fanout29/X _07134_/Y vssd1 vssd1 vccd1 vccd1 _07473_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10490__A1 _07198_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10490__B2 _10599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09211_ reg1_val[8] reg1_val[23] _09211_/S vssd1 vssd1 vccd1 vccd1 _09211_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09142_ _09143_/A _09143_/B vssd1 vssd1 vccd1 vccd1 _09142_/X sky130_fd_sc_hd__and2_1
XFILLER_0_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11990__A1 _11990_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09073_ _10749_/A _09073_/B vssd1 vssd1 vccd1 vccd1 _09075_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12870__B _12870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08024_ _08095_/A _08025_/B vssd1 vssd1 vccd1 vccd1 _08024_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09935__A1 _10337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10545__A2 _10415_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09975_ _11582_/A _09975_/B vssd1 vssd1 vccd1 vccd1 _09976_/B sky130_fd_sc_hd__xnor2_2
X_08926_ _08909_/A _08909_/B _08910_/Y vssd1 vssd1 vccd1 vccd1 _09032_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__07980__A _08564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08857_ _09673_/A _08857_/B vssd1 vssd1 vccd1 vccd1 _08867_/A sky130_fd_sc_hd__xnor2_2
X_07808_ _07878_/A _07878_/B vssd1 vssd1 vccd1 vccd1 _07879_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_79_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08788_ _08076_/A _08076_/B _08180_/Y vssd1 vssd1 vccd1 vccd1 _08788_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08123__B1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07739_ _07739_/A _07739_/B vssd1 vssd1 vccd1 vccd1 _07819_/A sky130_fd_sc_hd__nor2_1
X_10750_ _10751_/A _10751_/B vssd1 vssd1 vccd1 vccd1 _10874_/B sky130_fd_sc_hd__and2_1
XFILLER_0_55_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10549__C _10581_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10681_ _10681_/A vssd1 vssd1 vccd1 vccd1 _10681_/Y sky130_fd_sc_hd__inv_2
X_09409_ _09409_/A vssd1 vssd1 vccd1 vccd1 _09409_/Y sky130_fd_sc_hd__inv_2
X_12420_ _12420_/A0 _09422_/B _12438_/B vssd1 vssd1 vccd1 vccd1 _12420_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12351_ _12244_/A _12298_/A _12297_/A vssd1 vssd1 vccd1 vccd1 _12351_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_50_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11302_ _11301_/B _11302_/B vssd1 vssd1 vccd1 vccd1 _11303_/B sky130_fd_sc_hd__and2b_1
X_12282_ _12335_/B _12282_/B vssd1 vssd1 vccd1 vccd1 _12284_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11677__A _12336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11233_ _11234_/A _11271_/B vssd1 vssd1 vccd1 vccd1 _11233_/X sky130_fd_sc_hd__or2_1
XANTENNA__10581__A _10581_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11164_ _11406_/A fanout10/X fanout5/X _11309_/A vssd1 vssd1 vccd1 vccd1 _11165_/B
+ sky130_fd_sc_hd__o22a_1
X_11095_ _11096_/A _11096_/B vssd1 vssd1 vccd1 vccd1 _11095_/Y sky130_fd_sc_hd__nand2b_1
X_10115_ _11393_/A _10115_/B vssd1 vssd1 vccd1 vccd1 _10116_/B sky130_fd_sc_hd__xnor2_2
X_10046_ _10821_/A _10184_/B vssd1 vssd1 vccd1 vccd1 _10046_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_117_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06912__A1 _06944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11997_ _07036_/A _09257_/S _11996_/X _06680_/B vssd1 vssd1 vccd1 vccd1 _11997_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12446__C1 _12446_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10948_ fanout34/X fanout17/X fanout14/X fanout36/X vssd1 vssd1 vccd1 vccd1 _10949_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_58_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06683__A2_N _06810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09610__A _09936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10879_ _10879_/A _10879_/B vssd1 vssd1 vccd1 vccd1 _10892_/A sky130_fd_sc_hd__xor2_1
XANTENNA__13132__A _13147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12618_ _12621_/D _12618_/B vssd1 vssd1 vccd1 vccd1 new_PC[23] sky130_fd_sc_hd__xnor2_4
XFILLER_0_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08417__A1 _08649_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08417__B2 _08657_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12549_ _12708_/B _12550_/B vssd1 vssd1 vccd1 vccd1 _12560_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_53_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_1 _07262_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10491__A _12087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06972_ _07222_/A _07283_/A _06972_/C _07117_/C vssd1 vssd1 vccd1 vccd1 _06974_/B
+ sky130_fd_sc_hd__or4_4
X_09760_ _12356_/B1 _09714_/X _09715_/Y _09759_/X vssd1 vssd1 vccd1 vccd1 _09760_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11488__B1 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09691_ _09531_/A _09531_/B _09530_/A vssd1 vssd1 vccd1 vccd1 _09701_/A sky130_fd_sc_hd__a21o_1
X_08711_ _08711_/A _08711_/B vssd1 vssd1 vccd1 vccd1 _12129_/B sky130_fd_sc_hd__xnor2_2
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08642_ _09302_/A _08652_/A _08652_/B vssd1 vssd1 vccd1 vccd1 _08646_/B sky130_fd_sc_hd__mux2_1
XANTENNA_fanout164_A _11990_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08573_ _08664_/A _08573_/B vssd1 vssd1 vccd1 vccd1 _08608_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07305__A _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12452__A2 _07147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12988__B1 _13257_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07459__A2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07524_ _09943_/B2 _09661_/B2 fanout98/X _09650_/A vssd1 vssd1 vccd1 vccd1 _07525_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07455_ _10479_/A _07455_/B vssd1 vssd1 vccd1 vccd1 _07461_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07959__B _07959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09605__B1 _10049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07386_ _07384_/A _07384_/B _07469_/A vssd1 vssd1 vccd1 vccd1 _07402_/A sky130_fd_sc_hd__o21bai_2
XANTENNA__07040__A _07604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09125_ _09125_/A _09125_/B vssd1 vssd1 vccd1 vccd1 _09126_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07631__A2 _07221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09056_ _09057_/B _09056_/B vssd1 vssd1 vccd1 vccd1 _09058_/A sky130_fd_sc_hd__and2b_1
XANTENNA__11497__A _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09908__A1 _11752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08007_ _08016_/A _08016_/B vssd1 vssd1 vccd1 vccd1 _08009_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__11191__A2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09958_ _09959_/A _09959_/B vssd1 vssd1 vccd1 vccd1 _09958_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout77_A _07270_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08909_ _08909_/A _08909_/B vssd1 vssd1 vccd1 vccd1 _08911_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_99_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09889_ _12322_/A1 _10166_/C hold300/A vssd1 vssd1 vccd1 vccd1 _09889_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__08344__B1 _08334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11920_ _09149_/Y _11891_/Y _11892_/X _11895_/X _11919_/X vssd1 vssd1 vccd1 vccd1
+ _11920_/X sky130_fd_sc_hd__a311o_1
X_11851_ _11851_/A _11851_/B vssd1 vssd1 vccd1 vccd1 _11860_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11782_ _11783_/A _11783_/B vssd1 vssd1 vccd1 vccd1 _11872_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_95_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10802_ _10802_/A vssd1 vssd1 vccd1 vccd1 _10802_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08647__A1 _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10733_ _10734_/A _10734_/B vssd1 vssd1 vccd1 vccd1 _10733_/X sky130_fd_sc_hd__and2_1
X_10664_ _10900_/A _10664_/B vssd1 vssd1 vccd1 vccd1 _11050_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_36_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13383_ _13385_/CLK _13383_/D vssd1 vssd1 vccd1 vccd1 hold266/A sky130_fd_sc_hd__dfxtp_1
X_10595_ _10595_/A1 _08877_/B fanout6/X _07198_/Y vssd1 vssd1 vccd1 vccd1 _10596_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10206__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12403_ _06624_/B _12358_/X _06622_/X vssd1 vssd1 vccd1 vccd1 _12406_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__10206__B2 _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09072__A1 fanout63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09072__B2 fanout61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12334_ _12335_/B _12334_/B vssd1 vssd1 vccd1 vccd1 _12338_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_644 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12265_ _12444_/B _09880_/Y _12264_/X _12446_/C1 vssd1 vssd1 vccd1 vccd1 _12277_/A
+ sky130_fd_sc_hd__o211a_1
X_11216_ _11217_/B _11217_/A vssd1 vssd1 vccd1 vccd1 _11216_/Y sky130_fd_sc_hd__nand2b_1
X_12196_ _12192_/X _12195_/X _12064_/S vssd1 vssd1 vccd1 vccd1 _12196_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11147_ _13310_/Q _11147_/B vssd1 vssd1 vccd1 vccd1 _11251_/B sky130_fd_sc_hd__or2_1
XANTENNA__11854__B fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11078_ fanout34/X fanout14/X fanout12/X fanout36/X vssd1 vssd1 vccd1 vccd1 _11079_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08335__B1 _07274_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07138__A1 _08561_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07138__B2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13127__A _13147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10029_ hold290/A _10170_/C _09425_/C vssd1 vssd1 vccd1 vccd1 _10031_/B sky130_fd_sc_hd__o21a_1
XANTENNA__07689__A2 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07125__A _11584_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10693__A1 _07233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10445__A1 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09835__B1 _07262_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12685__B _12685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10445__B2 _10159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07240_ _09341_/A _07240_/B vssd1 vssd1 vccd1 vccd1 _07241_/B sky130_fd_sc_hd__xnor2_4
X_07171_ _07171_/A vssd1 vssd1 vccd1 vccd1 _07171_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12198__A1 _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09812_ _09650_/A fanout14/X fanout13/X _09943_/B2 vssd1 vssd1 vccd1 vccd1 _09813_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07019__B _07020_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08574__B1 _07166_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11764__B _11946_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06955_ instruction[24] _12359_/A is_load _06783_/B _06954_/X vssd1 vssd1 vccd1 vccd1
+ _06956_/B sky130_fd_sc_hd__a32o_2
XANTENNA__06858__B _07016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout281_A _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09743_ _12438_/A _09743_/B _09743_/C vssd1 vssd1 vccd1 vccd1 _09743_/X sky130_fd_sc_hd__or3_1
X_06886_ _12313_/A _06885_/Y _06867_/Y vssd1 vssd1 vccd1 vccd1 _12359_/B sky130_fd_sc_hd__o21ai_1
X_09674_ _09675_/A _09675_/B vssd1 vssd1 vccd1 vccd1 _09674_/Y sky130_fd_sc_hd__nor2_1
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07035__A _07036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10684__A1 _11820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08625_ _08630_/A _08625_/B vssd1 vssd1 vccd1 vccd1 _08638_/A sky130_fd_sc_hd__xnor2_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ _08556_/A _08556_/B vssd1 vssd1 vccd1 vccd1 _08587_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_76_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09250__A _11138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07507_ _07507_/A _07507_/B vssd1 vssd1 vccd1 vccd1 _07518_/A sky130_fd_sc_hd__xor2_1
XANTENNA__06593__B _06944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08487_ _08454_/A _08524_/A _08525_/A vssd1 vssd1 vccd1 vccd1 _08498_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07438_ _07438_/A _07438_/B vssd1 vssd1 vccd1 vccd1 _07562_/A sky130_fd_sc_hd__or2_2
XFILLER_0_92_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07369_ _07367_/Y _07369_/B vssd1 vssd1 vccd1 vccd1 _07370_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_18_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09054__A1 _07121_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09054__B2 _07417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09108_ _09108_/A _09108_/B vssd1 vssd1 vccd1 vccd1 _09109_/B sky130_fd_sc_hd__xor2_2
X_10380_ _10381_/A _10381_/B vssd1 vssd1 vccd1 vccd1 _10380_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_5_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06812__B1 _06810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09039_ _09708_/A _09039_/B vssd1 vssd1 vccd1 vccd1 _09040_/D sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12050_ _12050_/A _12050_/B _12050_/C vssd1 vssd1 vccd1 vccd1 _12050_/X sky130_fd_sc_hd__and3_2
XANTENNA__11164__A2 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11001_ _11117_/A _11001_/B vssd1 vssd1 vccd1 vccd1 _11004_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10372__B1 fanout74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12952_ hold268/A hold62/X vssd1 vssd1 vccd1 vccd1 _12953_/B sky130_fd_sc_hd__nand2b_1
X_11903_ _11903_/A _11903_/B vssd1 vssd1 vccd1 vccd1 _11905_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12883_ hold266/X hold24/X vssd1 vssd1 vccd1 vccd1 _13211_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__08983__B _08983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ _11637_/A _11814_/Y _11821_/X _11833_/X vssd1 vssd1 vccd1 vccd1 _11834_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13074__C1 _13142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11765_ _11766_/A _11766_/B vssd1 vssd1 vccd1 vccd1 _11767_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_83_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12821__C1 _13147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09293__B2 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09293__A1 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11696_ _11785_/B _11696_/B vssd1 vssd1 vccd1 vccd1 _11698_/C sky130_fd_sc_hd__nand2b_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ _11592_/A _07171_/A fanout38/X _10944_/B2 vssd1 vssd1 vccd1 vccd1 _10717_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10647_ _10647_/A _10647_/B vssd1 vssd1 vccd1 vccd1 _10649_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13366_ _13369_/CLK _13366_/D vssd1 vssd1 vccd1 vccd1 hold248/A sky130_fd_sc_hd__dfxtp_1
X_10578_ _12365_/A _10551_/Y _10552_/X _10577_/X vssd1 vssd1 vccd1 vccd1 _10578_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08504__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12317_ _12259_/X _12260_/Y _12262_/B vssd1 vssd1 vccd1 vccd1 _12366_/C sky130_fd_sc_hd__o21ai_2
X_13297_ _13304_/CLK _13297_/D vssd1 vssd1 vccd1 vccd1 hold293/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12248_ _11972_/B _12114_/B _12350_/A _12247_/X vssd1 vssd1 vccd1 vccd1 _12249_/B
+ sky130_fd_sc_hd__a31oi_4
XANTENNA__11865__A _12335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12179_ _12300_/A _12300_/B vssd1 vssd1 vccd1 vccd1 _12302_/B sky130_fd_sc_hd__nor2_1
XANTENNA__12460__S _12520_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08020__A2 _08457_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06740_ _06927_/A _06817_/B1 _12714_/B _06739_/X vssd1 vssd1 vccd1 vccd1 _11038_/A
+ sky130_fd_sc_hd__a31o_4
X_06671_ _12207_/S _06671_/B vssd1 vssd1 vccd1 vccd1 _06672_/D sky130_fd_sc_hd__or2_2
XANTENNA__09520__A2 _07269_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08410_ _08454_/A _08410_/B vssd1 vssd1 vccd1 vccd1 _08449_/A sky130_fd_sc_hd__xnor2_1
X_09390_ _09180_/X _09200_/X _09403_/S vssd1 vssd1 vccd1 vccd1 _09390_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09808__B1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08341_ _08575_/A _08341_/B vssd1 vssd1 vccd1 vccd1 _08393_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11091__A1 _11476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11091__B2 _11406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10969__A2 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08272_ _08272_/A _08272_/B vssd1 vssd1 vccd1 vccd1 _08284_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_116_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07223_ _07959_/B _10337_/A fanout29/X _12823_/A1 vssd1 vssd1 vccd1 vccd1 _07224_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07154_ reg1_val[26] _07154_/B vssd1 vssd1 vccd1 vccd1 _07155_/C sky130_fd_sc_hd__xor2_2
XFILLER_0_112_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07085_ reg1_val[8] _07105_/D _07248_/A vssd1 vssd1 vccd1 vccd1 _07086_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_42_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12343__A1 _07316_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout124 _10209_/A vssd1 vssd1 vccd1 vccd1 _11381_/A sky130_fd_sc_hd__buf_12
Xfanout135 _08454_/A vssd1 vssd1 vccd1 vccd1 _10749_/A sky130_fd_sc_hd__buf_12
Xfanout146 _07074_/X vssd1 vssd1 vccd1 vccd1 _09650_/A sky130_fd_sc_hd__buf_8
Xfanout179 _09152_/Y vssd1 vssd1 vccd1 vccd1 _12379_/B2 sky130_fd_sc_hd__clkbuf_8
Xfanout168 _12805_/Y vssd1 vssd1 vccd1 vccd1 _13101_/B2 sky130_fd_sc_hd__clkbuf_8
Xfanout157 _11893_/A vssd1 vssd1 vccd1 vccd1 _11630_/A sky130_fd_sc_hd__buf_4
X_07987_ _09670_/A _07987_/B vssd1 vssd1 vccd1 vccd1 _07988_/C sky130_fd_sc_hd__xnor2_1
X_06938_ instruction[27] _06944_/B vssd1 vssd1 vccd1 vccd1 _06938_/X sky130_fd_sc_hd__or2_1
X_09726_ _09248_/A _09725_/X _10297_/S vssd1 vssd1 vccd1 vccd1 _09726_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10657__A1 _10415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06869_ reg1_val[26] _07046_/B vssd1 vssd1 vccd1 vccd1 _06869_/X sky130_fd_sc_hd__and2_1
XFILLER_0_69_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09657_ _10246_/A _09657_/B vssd1 vssd1 vccd1 vccd1 _09658_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ _06809_/Y _09587_/X _11637_/A vssd1 vssd1 vccd1 vccd1 _09588_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08608_ _08608_/A _08608_/B vssd1 vssd1 vccd1 vccd1 _08619_/A sky130_fd_sc_hd__xor2_1
XANTENNA__13071__A2 _12826_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _08580_/A _08539_/B vssd1 vssd1 vccd1 vccd1 _08569_/A sky130_fd_sc_hd__xnor2_2
X_11550_ _11650_/B _11649_/B hold264/A vssd1 vssd1 vccd1 vccd1 _11552_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10501_ _10501_/A _10501_/B _10501_/C vssd1 vssd1 vccd1 vccd1 _10503_/A sky130_fd_sc_hd__and3_1
XFILLER_0_80_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13220_ _13220_/A _13220_/B vssd1 vssd1 vccd1 vccd1 _13221_/B sky130_fd_sc_hd__nand2_1
X_11481_ _12169_/A _07171_/A fanout38/X _06998_/X vssd1 vssd1 vccd1 vccd1 _11482_/B
+ sky130_fd_sc_hd__a22o_1
X_10432_ _11029_/S _10292_/X _10431_/X vssd1 vssd1 vccd1 vccd1 _10432_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_103_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13151_ hold279/X _13248_/B1 _13150_/X _13248_/A2 vssd1 vssd1 vccd1 vccd1 hold280/A
+ sky130_fd_sc_hd__a22o_1
X_10363_ _10363_/A _10363_/B vssd1 vssd1 vccd1 vccd1 _10366_/A sky130_fd_sc_hd__nor2_1
X_12102_ _12102_/A _12102_/B vssd1 vssd1 vccd1 vccd1 _12103_/B sky130_fd_sc_hd__nor2_1
X_13082_ hold89/X _13094_/A2 _13250_/B hold123/X _13142_/A vssd1 vssd1 vccd1 vccd1
+ hold124/A sky130_fd_sc_hd__o221a_1
XFILLER_0_20_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12033_ _12033_/A _12033_/B vssd1 vssd1 vccd1 vccd1 _12034_/B sky130_fd_sc_hd__or2_1
X_10294_ _09719_/X _09721_/X _10294_/S vssd1 vssd1 vccd1 vccd1 _10294_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08538__B1 _09472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12935_ _13163_/A _13164_/A _13163_/B vssd1 vssd1 vccd1 vccd1 _13169_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__11845__B1 _07316_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07513__B2 _10338_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07513__A1 _10595_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12866_ hold28/X _12870_/B vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__or2_1
XFILLER_0_34_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11817_ _11817_/A _11817_/B vssd1 vssd1 vccd1 vccd1 _11819_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_8_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11073__A1 _11764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11073__B2 _11592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12797_ hold167/X hold140/X vssd1 vssd1 vccd1 vccd1 _12797_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_56_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11748_ _11720_/Y _11721_/X _11723_/Y _12365_/A _11747_/X vssd1 vssd1 vccd1 vccd1
+ _11748_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_43_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11679_ _12093_/A _11679_/B vssd1 vssd1 vccd1 vccd1 _11681_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13349_ _13354_/CLK hold105/X vssd1 vssd1 vccd1 vccd1 hold103/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08241__A2 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07910_ _08656_/A _07910_/B _07910_/C vssd1 vssd1 vccd1 vccd1 _07913_/B sky130_fd_sc_hd__or3_1
X_08890_ _08890_/A _08890_/B vssd1 vssd1 vccd1 vccd1 _08891_/B sky130_fd_sc_hd__nor2_1
X_07841_ _07842_/A _07841_/B _07841_/C vssd1 vssd1 vccd1 vccd1 _07885_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_75_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07772_ _08664_/A _07772_/B vssd1 vssd1 vccd1 vccd1 _07777_/A sky130_fd_sc_hd__xnor2_1
X_06723_ _06723_/A _12645_/B vssd1 vssd1 vccd1 vccd1 _06723_/Y sky130_fd_sc_hd__nor2_1
X_09511_ _09511_/A _09511_/B vssd1 vssd1 vccd1 vccd1 _09529_/A sky130_fd_sc_hd__xor2_1
XANTENNA__10939__A _12336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06654_ _06723_/A _12685_/B vssd1 vssd1 vccd1 vccd1 _06654_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_91_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09442_ curr_PC[0] curr_PC[1] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _09762_/B sky130_fd_sc_hd__and3_1
X_06585_ rst vssd1 vssd1 vccd1 vccd1 _06585_/Y sky130_fd_sc_hd__inv_2
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09373_ _09034_/A _09034_/B _09146_/A _09146_/B vssd1 vssd1 vccd1 vccd1 _09711_/C
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout244_A _06958_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13053__A2 _12820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08324_ _08360_/A _08360_/B _08285_/Y vssd1 vssd1 vccd1 vccd1 _08689_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_19_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08255_ _08255_/A _08255_/B vssd1 vssd1 vccd1 vccd1 _08317_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_104_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07206_ reg1_val[18] reg1_val[31] _12359_/A vssd1 vssd1 vccd1 vccd1 _07208_/C sky130_fd_sc_hd__and3_1
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08186_ _08186_/A _08186_/B vssd1 vssd1 vccd1 vccd1 _08188_/B sky130_fd_sc_hd__xnor2_2
X_07137_ _07136_/B _11854_/A _11929_/A vssd1 vssd1 vccd1 vccd1 _07137_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_42_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07068_ _10072_/A _07068_/B vssd1 vssd1 vccd1 vccd1 _07068_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10327__B1 _10276_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10981_ _11102_/A _10981_/B vssd1 vssd1 vccd1 vccd1 _10983_/B sky130_fd_sc_hd__or2_1
XANTENNA__09496__A1 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09496__B2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09709_ _09370_/X _09546_/X _09547_/X vssd1 vssd1 vccd1 vccd1 _09709_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09422__B _09422_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12720_ _12721_/A _12721_/B _12721_/C vssd1 vssd1 vccd1 vccd1 _12722_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12651_ _12649_/Y _12651_/B vssd1 vssd1 vccd1 vccd1 _12652_/B sky130_fd_sc_hd__and2b_1
X_11602_ _11603_/B _11603_/A vssd1 vssd1 vccd1 vccd1 _11698_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_65_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13044__A2 _06577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12582_ _12582_/A _12582_/B vssd1 vssd1 vccd1 vccd1 _12597_/B sky130_fd_sc_hd__or2_1
XFILLER_0_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10584__A _12157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11533_ _11711_/A _11533_/B vssd1 vssd1 vccd1 vccd1 _11567_/D sky130_fd_sc_hd__xor2_4
XFILLER_0_37_188 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11464_ hold292/A _11549_/C _11650_/B vssd1 vssd1 vccd1 vccd1 _11464_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13203_ _13203_/A _13203_/B vssd1 vssd1 vccd1 vccd1 _13203_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10415_ _10415_/A _10415_/B vssd1 vssd1 vccd1 vccd1 _10661_/C sky130_fd_sc_hd__xnor2_4
XFILLER_0_33_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11395_ _11395_/A _11395_/B vssd1 vssd1 vccd1 vccd1 _11396_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_21_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10346_ _10247_/B _10247_/C _10247_/A vssd1 vssd1 vccd1 vccd1 _10355_/A sky130_fd_sc_hd__a21bo_1
X_13134_ _13134_/A _13134_/B vssd1 vssd1 vccd1 vccd1 _13134_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__06785__A2 _06783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07982__A1 _07080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ _10950_/A _13101_/B2 hold131/X vssd1 vssd1 vccd1 vccd1 hold132/A sky130_fd_sc_hd__o21a_1
X_10277_ _10542_/A _10661_/A vssd1 vssd1 vccd1 vccd1 _10541_/A sky130_fd_sc_hd__nor2_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12016_ fanout68/X fanout10/X fanout5/X _12087_/A vssd1 vssd1 vccd1 vccd1 _12017_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07117__B _07147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13316_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09613__A _09922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12918_ _12907_/B _13120_/B _12905_/X vssd1 vssd1 vccd1 vccd1 _13124_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_75_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12849_ _11764_/A _12863_/A2 hold53/X _13210_/A vssd1 vssd1 vccd1 vccd1 _13285_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06691__B _07016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08040_ _08664_/A _08040_/B vssd1 vssd1 vccd1 vccd1 _08046_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09991_ _09991_/A _09991_/B vssd1 vssd1 vccd1 vccd1 _09992_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_3_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07422__B1 _07175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10433__S _11820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08942_ _08942_/A _08942_/B vssd1 vssd1 vccd1 vccd1 _09018_/A sky130_fd_sc_hd__nor2_2
XANTENNA__12849__A2 _12863_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08411__B _08411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout194_A _12205_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08873_ _12336_/A _08874_/B vssd1 vssd1 vccd1 vccd1 _08876_/A sky130_fd_sc_hd__or2_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07725__B2 _07173_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07725__A1 _07166_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12868__B _12870_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07824_ _07824_/A _07824_/B vssd1 vssd1 vccd1 vccd1 _07828_/B sky130_fd_sc_hd__xnor2_2
X_07755_ _07755_/A _07755_/B vssd1 vssd1 vccd1 vccd1 _07866_/B sky130_fd_sc_hd__xnor2_2
X_06706_ reg1_val[19] _07078_/A vssd1 vssd1 vccd1 vccd1 _06707_/B sky130_fd_sc_hd__and2b_1
XANTENNA__09242__B _09242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07686_ _08580_/A _07686_/B vssd1 vssd1 vccd1 vccd1 _07688_/B sky130_fd_sc_hd__xnor2_2
X_06637_ reg1_val[30] _08973_/C vssd1 vssd1 vccd1 vccd1 _12438_/B sky130_fd_sc_hd__and2_1
XFILLER_0_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09425_ hold235/A hold245/A _09425_/C vssd1 vssd1 vccd1 vccd1 _09425_/X sky130_fd_sc_hd__and3_1
XANTENNA__08139__A _08580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13026__A2 _13171_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09356_ _09130_/A _09129_/B _09127_/Y vssd1 vssd1 vccd1 vccd1 _09366_/A sky130_fd_sc_hd__a21o_2
XANTENNA__07978__A _08580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11588__A2 fanout10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08307_ _08515_/A2 _08561_/A2 _09940_/B2 _08540_/B vssd1 vssd1 vccd1 vccd1 _08308_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08453__A2 _08484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09287_ fanout56/X _09943_/B2 _09650_/A fanout68/X vssd1 vssd1 vccd1 vccd1 _09288_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08238_ _08649_/B1 _08289_/B fanout75/X _09404_/S vssd1 vssd1 vccd1 vccd1 _08239_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_90_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10200_ _11484_/A _10200_/B vssd1 vssd1 vccd1 vccd1 _10201_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_43_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08169_ _08169_/A _08169_/B vssd1 vssd1 vccd1 vccd1 _08172_/A sky130_fd_sc_hd__nor2_2
X_11180_ _11180_/A _11180_/B vssd1 vssd1 vccd1 vccd1 _11183_/A sky130_fd_sc_hd__nor2_1
X_10131_ _10132_/B _10132_/A vssd1 vssd1 vccd1 vccd1 _10131_/X sky130_fd_sc_hd__and2b_1
X_10062_ _11179_/A _10062_/B vssd1 vssd1 vccd1 vccd1 _10065_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09433__A _12365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11276__B2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11276__A1 _07051_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06776__B _06810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10964_ _06998_/X fanout32/X fanout30/X _07032_/Y vssd1 vssd1 vccd1 vccd1 _10965_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12703_ _12711_/A _12703_/B vssd1 vssd1 vccd1 vccd1 _12705_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08049__A _10092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10895_ _10897_/A _10897_/B _10897_/C vssd1 vssd1 vccd1 vccd1 _10898_/A sky130_fd_sc_hd__a21oi_1
X_12634_ _12634_/A _12634_/B vssd1 vssd1 vccd1 vccd1 _12636_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_66_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11579__A2 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12565_ _12572_/A _12565_/B vssd1 vssd1 vccd1 vccd1 _12567_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_66_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11516_ _11516_/A _11516_/B vssd1 vssd1 vccd1 vccd1 _11518_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12496_ _12497_/A _12497_/B _12497_/C vssd1 vssd1 vccd1 vccd1 _12504_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_41_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11447_ _11813_/S _11447_/B vssd1 vssd1 vccd1 vccd1 _11447_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_40_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11378_ fanout30/X _07316_/Y _07608_/Y fanout32/X vssd1 vssd1 vccd1 vccd1 _11379_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13117_ hold295/A _13116_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13117_/X sky130_fd_sc_hd__mux2_1
X_10329_ _10661_/A _10661_/B vssd1 vssd1 vccd1 vccd1 _10329_/Y sky130_fd_sc_hd__nor2_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ hold43/A _06577_/A rst vssd1 vssd1 vccd1 vccd1 _13048_/Y sky130_fd_sc_hd__a21oi_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10711__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06967__A _12644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11592__B _12428_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10489__A _12157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12688__B _12689_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12464__A0 _12644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07540_ _07540_/A _07540_/B vssd1 vssd1 vccd1 vccd1 _07556_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_72_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13008__A2 _13171_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09880__A1 _11029_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07471_ _11381_/A _07471_/B vssd1 vssd1 vccd1 vccd1 _07475_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10490__A2 _08877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09210_ reg1_val[9] reg1_val[22] _09211_/S vssd1 vssd1 vccd1 vccd1 _09210_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07891__B1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07798__A _09836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09141_ _09141_/A _09141_/B vssd1 vssd1 vccd1 vccd1 _09143_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09072_ fanout63/X _10473_/B2 _10240_/A fanout61/X vssd1 vssd1 vccd1 vccd1 _09073_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08023_ _08023_/A _08023_/B vssd1 vssd1 vccd1 vccd1 _08025_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11727__C1 _09225_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10952__A _11179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout207_A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_139 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10163__S _10297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09974_ fanout52/X fanout28/X fanout26/X _11476_/A vssd1 vssd1 vccd1 vccd1 _09975_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08925_ _08912_/A _08912_/B _08913_/Y vssd1 vssd1 vccd1 vccd1 _09034_/A sky130_fd_sc_hd__a21bo_2
X_08856_ _09298_/A1 fanout56/X fanout17/X _09298_/B2 vssd1 vssd1 vccd1 vccd1 _08857_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_98_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07807_ _07807_/A _07807_/B vssd1 vssd1 vccd1 vccd1 _07878_/B sky130_fd_sc_hd__xnor2_1
X_08787_ _08783_/A _08783_/B _08786_/Y _11810_/A _11809_/B vssd1 vssd1 vccd1 vccd1
+ _08795_/A sky130_fd_sc_hd__a2111o_2
XFILLER_0_79_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08123__A1 _08649_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08123__B2 _09404_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07738_ _07737_/A _07737_/C _07737_/B vssd1 vssd1 vccd1 vccd1 _07739_/B sky130_fd_sc_hd__a21oi_1
X_07669_ _07669_/A _07669_/B vssd1 vssd1 vccd1 vccd1 _07671_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12207__A0 _09228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10680_ _09568_/X _09574_/X _11246_/S vssd1 vssd1 vccd1 vccd1 _10681_/A sky130_fd_sc_hd__mux2_1
X_09408_ _09393_/X _09407_/X _11247_/A vssd1 vssd1 vccd1 vccd1 _09409_/A sky130_fd_sc_hd__mux2_1
XANTENNA_fanout22_A _12428_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09339_ _09834_/A _09339_/B vssd1 vssd1 vccd1 vccd1 _09343_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12350_ _12350_/A _12350_/B vssd1 vssd1 vccd1 vccd1 _12350_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11301_ _11302_/B _11301_/B vssd1 vssd1 vccd1 vccd1 _11303_/A sky130_fd_sc_hd__and2b_1
XANTENNA__10862__A _12017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12281_ fanout12/X fanout10/X fanout5/X _12335_/A vssd1 vssd1 vccd1 vccd1 _12282_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_62_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11232_ _11433_/A _11232_/B vssd1 vssd1 vccd1 vccd1 _11271_/B sky130_fd_sc_hd__xnor2_4
X_11163_ _11052_/B _11124_/Y _11893_/A vssd1 vssd1 vccd1 vccd1 _11234_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__10581__B _10581_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10114_ fanout47/X _11309_/A _11198_/A fanout45/X vssd1 vssd1 vccd1 vccd1 _10115_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11094_ _11094_/A _11094_/B vssd1 vssd1 vccd1 vccd1 _11096_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12289__A3 _12158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10045_ curr_PC[4] curr_PC[5] _10045_/C vssd1 vssd1 vccd1 vccd1 _10184_/B sky130_fd_sc_hd__and3_1
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
X_11996_ _11995_/A _09228_/X _11995_/Y _12421_/A1 vssd1 vssd1 vccd1 vccd1 _11996_/X
+ sky130_fd_sc_hd__o211a_1
X_10947_ _10947_/A _10947_/B vssd1 vssd1 vccd1 vccd1 _10956_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12617_ _12609_/B _12614_/B _12607_/X vssd1 vssd1 vccd1 vccd1 _12618_/B sky130_fd_sc_hd__a21o_1
X_10878_ _10878_/A _10878_/B vssd1 vssd1 vccd1 vccd1 _10879_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_54_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07411__A _09779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11928__A_N _11929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08417__A2 _10221_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12548_ reg1_val[13] curr_PC[13] _12638_/S vssd1 vssd1 vccd1 vccd1 _12550_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_53_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11868__A _11868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ _12655_/B _12480_/B vssd1 vssd1 vccd1 vccd1 _12490_/A sky130_fd_sc_hd__nand2_1
XANTENNA_2 _07268_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09378__B1 _09150_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12382__C1 _12631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08242__A _08664_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06971_ _07165_/A _07172_/A _07149_/A _07959_/A vssd1 vssd1 vccd1 vccd1 _07133_/A
+ sky130_fd_sc_hd__or4_4
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11488__B2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11488__A1 _12233_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08710_ _09037_/A _08710_/B vssd1 vssd1 vccd1 vccd1 _12364_/B sky130_fd_sc_hd__xor2_2
X_09690_ _09690_/A _09690_/B vssd1 vssd1 vccd1 vccd1 _09703_/A sky130_fd_sc_hd__xor2_4
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08641_ _12808_/A _08641_/B vssd1 vssd1 vccd1 vccd1 _08652_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09550__B1 _09371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09073__A _10749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10012__A _12438_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08572_ _07983_/A _07121_/Y _07282_/Y _12642_/A vssd1 vssd1 vccd1 vccd1 _08573_/B
+ sky130_fd_sc_hd__a22o_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12638__S _12638_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07523_ _07526_/A _07526_/B vssd1 vssd1 vccd1 vccd1 _07734_/B sky130_fd_sc_hd__or2_1
X_07454_ _10245_/B2 fanout98/X _10245_/A1 fanout84/X vssd1 vssd1 vccd1 vccd1 _07455_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_119_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07321__A _09947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07385_ _07468_/A _07468_/B vssd1 vssd1 vccd1 vccd1 _07469_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07616__B1 _10240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09124_ _09125_/B _09125_/A vssd1 vssd1 vccd1 vccd1 _09124_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_115_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09055_ _09779_/A _09055_/B vssd1 vssd1 vccd1 vccd1 _09056_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_114_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08006_ _08006_/A _08006_/B vssd1 vssd1 vccd1 vccd1 _08016_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11176__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10923__B1 _11648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08041__B1 fanout72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09957_ _09957_/A _09957_/B vssd1 vssd1 vccd1 vccd1 _09959_/B sky130_fd_sc_hd__xnor2_4
X_08908_ _07667_/A _07667_/B _07665_/X vssd1 vssd1 vccd1 vccd1 _08909_/B sky130_fd_sc_hd__a21oi_2
X_09888_ hold221/A hold237/A hold301/A hold293/A vssd1 vssd1 vccd1 vccd1 _10166_/C
+ sky130_fd_sc_hd__or4_2
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08839_ _08840_/A _08840_/B vssd1 vssd1 vccd1 vccd1 _08839_/Y sky130_fd_sc_hd__nor2_1
X_11850_ _11763_/A _11763_/B _11762_/A vssd1 vssd1 vccd1 vccd1 _11851_/B sky130_fd_sc_hd__o21a_1
X_11781_ _11781_/A _11781_/B vssd1 vssd1 vccd1 vccd1 _11783_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12548__S _12638_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10801_ _09723_/X _09729_/X _11246_/S vssd1 vssd1 vccd1 vccd1 _10802_/A sky130_fd_sc_hd__mux2_1
XANTENNA__08647__A2 _07166_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10732_ _11770_/A _10732_/B vssd1 vssd1 vccd1 vccd1 _10734_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10663_ _09554_/B _10138_/C _10661_/X _10662_/Y _10660_/Y vssd1 vssd1 vccd1 vccd1
+ _10664_/B sky130_fd_sc_hd__o311ai_4
X_13382_ _13385_/CLK _13382_/D vssd1 vssd1 vccd1 vccd1 hold268/A sky130_fd_sc_hd__dfxtp_1
X_12402_ _12398_/Y _12400_/X _12401_/Y vssd1 vssd1 vccd1 vccd1 _12402_/Y sky130_fd_sc_hd__a21oi_1
X_10594_ _10482_/A _10481_/B _10481_/A vssd1 vssd1 vccd1 vccd1 _10597_/A sky130_fd_sc_hd__a21boi_2
XANTENNA__10206__A2 fanout86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09072__A2 _10473_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12333_ fanout10/X fanout7/X fanout5/X fanout12/X vssd1 vssd1 vccd1 vccd1 _12334_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_50_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12264_ _12259_/X _12262_/X _12263_/Y vssd1 vssd1 vccd1 vccd1 _12264_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_50_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11215_ _11215_/A _11215_/B vssd1 vssd1 vccd1 vccd1 _11217_/B sky130_fd_sc_hd__xnor2_2
X_12195_ _12193_/Y _12195_/B vssd1 vssd1 vccd1 vccd1 _12195_/X sky130_fd_sc_hd__and2b_1
XANTENNA__08032__B1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11146_ _11146_/A _11146_/B vssd1 vssd1 vccd1 vccd1 _11146_/X sky130_fd_sc_hd__or2_1
XANTENNA__07109__C _07109_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11077_ _11194_/A _11077_/B vssd1 vssd1 vccd1 vccd1 _11087_/A sky130_fd_sc_hd__and2_1
XFILLER_0_37_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10028_ hold196/A _10028_/B vssd1 vssd1 vccd1 vccd1 _10028_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08335__B2 _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07138__A2 _07830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12419__B1 _11648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10693__A2 _12422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11979_ _06860_/A _11896_/X _11913_/S vssd1 vssd1 vccd1 vccd1 _11979_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_85_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09835__B2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09835__A1 _07959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06964__B _12359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07846__B1 _09479_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07141__A _11134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08237__A _10207_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06980__A _07097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07170_ _07170_/A _07170_/B vssd1 vssd1 vccd1 vccd1 _07170_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_42_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07074__A1 _09944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10933__C _10933_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09220__C1 _12446_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10905__B1 _09150_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09811_ _09811_/A _09811_/B vssd1 vssd1 vccd1 vccd1 _09819_/A sky130_fd_sc_hd__xor2_1
X_09742_ _09586_/A _09586_/B _06809_/A vssd1 vssd1 vccd1 vccd1 _09743_/C sky130_fd_sc_hd__a21boi_1
X_06954_ instruction[40] _06610_/X _06952_/X _06953_/Y vssd1 vssd1 vccd1 vccd1 _06954_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12222__A _12335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07316__A _10476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout274_A _13019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06885_ _06874_/A _06884_/X _06868_/Y vssd1 vssd1 vccd1 vccd1 _06885_/Y sky130_fd_sc_hd__a21boi_1
X_09673_ _09673_/A _09673_/B vssd1 vssd1 vccd1 vccd1 _09675_/B sky130_fd_sc_hd__xnor2_2
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _08624_/A _08624_/B vssd1 vssd1 vccd1 vccd1 _08725_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_77_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ _08556_/A _08556_/B vssd1 vssd1 vccd1 vccd1 _08568_/A sky130_fd_sc_hd__or2_1
XFILLER_0_77_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07506_ _07571_/A _07571_/B vssd1 vssd1 vccd1 vccd1 _07506_/X sky130_fd_sc_hd__and2_1
XFILLER_0_119_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10436__A2 _11990_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08486_ _08524_/A _08524_/B vssd1 vssd1 vccd1 vccd1 _08525_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08147__A _08334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_13_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13296_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07437_ _07424_/B _07437_/B vssd1 vssd1 vccd1 vccd1 _07438_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_45_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07368_ _07368_/A _07368_/B vssd1 vssd1 vccd1 vccd1 _07369_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_17_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09054__A2 fanout42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13199__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11397__B1 fanout38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09107_ _09108_/A _09108_/B vssd1 vssd1 vccd1 vccd1 _09107_/Y sky130_fd_sc_hd__nand2_1
X_07299_ _07298_/A _07298_/B _10060_/A vssd1 vssd1 vccd1 vccd1 _07299_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_103_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11149__B1 _11648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09038_ _08710_/B _09036_/Y _09035_/X vssd1 vssd1 vccd1 vccd1 _09039_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11000_ _11000_/A _11000_/B vssd1 vssd1 vccd1 vccd1 _11001_/B sky130_fd_sc_hd__or2_1
XANTENNA__09706__A _09707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10372__A1 _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10372__B2 fanout65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12951_ _13202_/A _13203_/A _13202_/B vssd1 vssd1 vccd1 vccd1 _13207_/A sky130_fd_sc_hd__a21bo_1
X_12882_ hold77/X hold254/X vssd1 vssd1 vccd1 vccd1 _12882_/X sky130_fd_sc_hd__and2b_1
X_11902_ reg1_val[22] curr_PC[22] vssd1 vssd1 vccd1 vccd1 _11903_/B sky130_fd_sc_hd__or2_1
X_11833_ _11827_/Y _11828_/X _11832_/X _11825_/X vssd1 vssd1 vccd1 vccd1 _11833_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11764_ _11764_/A _11946_/C _11764_/C vssd1 vssd1 vccd1 vccd1 _11766_/B sky130_fd_sc_hd__and3_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06620__A2_N _06766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09293__A2 _07092_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11695_ _11695_/A _11695_/B vssd1 vssd1 vccd1 vccd1 _11696_/B sky130_fd_sc_hd__or2_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _10715_/A _10715_/B vssd1 vssd1 vccd1 vccd1 _10719_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_83_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10646_ _10646_/A _10646_/B vssd1 vssd1 vccd1 vccd1 _10647_/B sky130_fd_sc_hd__and2_1
XANTENNA__09587__S _12054_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06635__A2_N _06783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10577_ _12446_/C1 _10564_/X _10576_/X _10556_/X vssd1 vssd1 vccd1 vccd1 _10577_/X
+ sky130_fd_sc_hd__a211o_1
X_13365_ _13365_/CLK _13365_/D vssd1 vssd1 vccd1 vccd1 hold290/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08253__B1 _08501_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13296_ _13296_/CLK _13296_/D vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__dfxtp_1
X_12316_ _12364_/A _09040_/A _08810_/B _12365_/A _12315_/Y vssd1 vssd1 vccd1 vccd1
+ _12331_/B sky130_fd_sc_hd__o311a_1
XFILLER_0_11_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12247_ _12116_/Y _12350_/A _12246_/X vssd1 vssd1 vccd1 vccd1 _12247_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09753__B1 _09422_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09616__A _09779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12178_ _12178_/A _12178_/B vssd1 vssd1 vccd1 vccd1 _12299_/A sky130_fd_sc_hd__or2_2
X_11129_ _11022_/A _11019_/X _11039_/S vssd1 vssd1 vccd1 vccd1 _11129_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07136__A _11929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12977__A _13001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11863__A1 _11770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06670_ reg1_val[26] _07046_/B vssd1 vssd1 vccd1 vccd1 _06671_/B sky130_fd_sc_hd__and2b_1
XANTENNA__12696__B _12696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06694__B _12670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09808__A1 fanout53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09808__B2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10418__A2 _10453_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08340_ _08657_/B _10338_/B2 _08457_/A2 _08649_/A2 vssd1 vssd1 vccd1 vccd1 _08341_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11091__A2 _07362_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08271_ _08327_/A _08327_/B _08268_/A vssd1 vssd1 vccd1 vccd1 _08284_/A sky130_fd_sc_hd__a21o_1
X_07222_ _07222_/A _07222_/B vssd1 vssd1 vccd1 vccd1 _10225_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_61_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07153_ _07155_/A _07155_/B vssd1 vssd1 vccd1 vccd1 _11398_/A sky130_fd_sc_hd__and2_4
XFILLER_0_6_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07084_ _07248_/A _07105_/D vssd1 vssd1 vccd1 vccd1 _07089_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_42_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10960__A _11582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12328__C1 _12422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12343__A2 _11946_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11551__B1 _12376_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout125 _07183_/X vssd1 vssd1 vccd1 vccd1 _10092_/A sky130_fd_sc_hd__clkbuf_16
Xfanout136 _10060_/A vssd1 vssd1 vccd1 vccd1 _08454_/A sky130_fd_sc_hd__buf_12
Xfanout147 _09943_/B2 vssd1 vssd1 vccd1 vccd1 _08598_/B sky130_fd_sc_hd__buf_6
Xfanout114 _07221_/X vssd1 vssd1 vccd1 vccd1 _09770_/B2 sky130_fd_sc_hd__buf_6
Xfanout169 _12805_/Y vssd1 vssd1 vccd1 vccd1 _13089_/A2 sky130_fd_sc_hd__buf_2
Xfanout158 _12364_/A vssd1 vssd1 vccd1 vccd1 _11893_/A sky130_fd_sc_hd__clkbuf_4
X_07986_ _08641_/B fanout80/X fanout76/X _08627_/A2 vssd1 vssd1 vccd1 vccd1 _07987_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_38_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06937_ instruction[19] _06590_/X _06936_/X _06716_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[1]
+ sky130_fd_sc_hd__o211a_4
X_09725_ _09395_/X _09397_/X _09725_/S vssd1 vssd1 vccd1 vccd1 _09725_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10657__A2 _10415_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09656_ fanout56/X _10245_/B2 _10245_/A1 fanout68/X vssd1 vssd1 vccd1 vccd1 _09657_/B
+ sky130_fd_sc_hd__o22a_1
X_06868_ reg1_val[27] _07049_/A vssd1 vssd1 vccd1 vccd1 _06868_/Y sky130_fd_sc_hd__nand2_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ _08677_/A _08677_/B vssd1 vssd1 vccd1 vccd1 _08607_/X sky130_fd_sc_hd__and2_1
XFILLER_0_96_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06799_ _06815_/A _06817_/B1 _12660_/B _06797_/X vssd1 vssd1 vccd1 vccd1 _07165_/A
+ sky130_fd_sc_hd__a31o_4
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ _06820_/X _09586_/Y _12054_/S vssd1 vssd1 vccd1 vccd1 _09587_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10200__A _11484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _08538_/A1 _08649_/B1 _09472_/A _08598_/B vssd1 vssd1 vccd1 vccd1 _08539_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_65_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08469_ _08469_/A _08469_/B vssd1 vssd1 vccd1 vccd1 _08470_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10500_ _10500_/A _12087_/B vssd1 vssd1 vccd1 vccd1 _10501_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_80_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11480_ _11600_/B _11480_/B vssd1 vssd1 vccd1 vccd1 _11492_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11909__A2 _12447_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10431_ _11247_/A _10431_/B vssd1 vssd1 vccd1 vccd1 _10431_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13150_ hold294/A _13149_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13150_/X sky130_fd_sc_hd__mux2_1
X_10362_ _10362_/A _10362_/B vssd1 vssd1 vccd1 vccd1 _10363_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_33_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12101_ _12101_/A _12101_/B _12101_/C vssd1 vssd1 vccd1 vccd1 _12102_/B sky130_fd_sc_hd__nor3_1
X_13081_ _11584_/A _13089_/A2 hold90/X vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__o21a_1
X_10293_ _11247_/A _10292_/X _09251_/A vssd1 vssd1 vccd1 vccd1 _10293_/X sky130_fd_sc_hd__o21a_1
X_12032_ _12033_/A _12033_/B vssd1 vssd1 vccd1 vccd1 _12111_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08538__A1 _08538_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08538__B2 _08598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold190 hold190/A vssd1 vssd1 vccd1 vccd1 hold190/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11542__B1 _09225_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12934_ hold106/X hold285/A vssd1 vssd1 vccd1 vccd1 _13163_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__11845__A1 _07051_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11845__B2 fanout43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07513__A2 _08411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12865_ _07316_/Y _12871_/A2 hold59/X _13246_/A vssd1 vssd1 vccd1 vccd1 _13293_/D
+ sky130_fd_sc_hd__o211a_1
X_11816_ reg1_val[21] curr_PC[21] vssd1 vssd1 vccd1 vccd1 _11817_/B sky130_fd_sc_hd__or2_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10110__A _11484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12796_ _12796_/A _12796_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[31] sky130_fd_sc_hd__xnor2_4
XFILLER_0_56_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11073__A2 _07417_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _11747_/A _11747_/B _11747_/C _11747_/D vssd1 vssd1 vccd1 vccd1 _11747_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_55_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08474__B1 _09940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11678_ _12233_/B _07175_/Y fanout17/X _07171_/Y vssd1 vssd1 vccd1 vccd1 _11679_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_70_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10629_ _11179_/A _10629_/B vssd1 vssd1 vccd1 vccd1 _10631_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13348_ _13354_/CLK hold115/X vssd1 vssd1 vccd1 vccd1 hold113/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10033__B1 _09422_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09974__B1 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12471__S _12471_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13279_ _13392_/CLK _13279_/D vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09346__A _11770_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07201__A1 _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07840_ _09673_/A _07840_/B vssd1 vssd1 vccd1 vccd1 _07841_/C sky130_fd_sc_hd__xor2_1
XANTENNA__12089__A1 _12009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07771_ _06993_/A fanout63/X fanout61/X _06993_/Y vssd1 vssd1 vccd1 vccd1 _07772_/B
+ sky130_fd_sc_hd__o22a_1
X_06722_ instruction[0] instruction[1] instruction[2] instruction[26] pred_val vssd1
+ vssd1 vccd1 vccd1 _12645_/B sky130_fd_sc_hd__o311a_4
XFILLER_0_79_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09510_ _09510_/A _09510_/B vssd1 vssd1 vccd1 vccd1 _09511_/B sky130_fd_sc_hd__xor2_1
XANTENNA__12500__A _12670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09081__A _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06653_ instruction[34] _06675_/B vssd1 vssd1 vccd1 vccd1 _12685_/B sky130_fd_sc_hd__and2_4
XANTENNA__06712__B1 _06783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13038__B1 _12820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09441_ _09260_/X _09440_/Y _10821_/A vssd1 vssd1 vccd1 vccd1 dest_val[1] sky130_fd_sc_hd__mux2_8
XFILLER_0_93_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06584_ _12438_/A vssd1 vssd1 vccd1 vccd1 _06584_/Y sky130_fd_sc_hd__inv_2
X_09372_ _09708_/A _09372_/B _09863_/A _08710_/B vssd1 vssd1 vccd1 vccd1 _09375_/A
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_86_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08323_ _08323_/A _08323_/B vssd1 vssd1 vccd1 vccd1 _08360_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout237_A _06993_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08254_ _08580_/A _08254_/B vssd1 vssd1 vccd1 vccd1 _08255_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_27_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07205_ reg1_val[14] reg1_val[15] _07141_/C _07109_/C _07248_/A vssd1 vssd1 vccd1
+ vccd1 _07228_/B sky130_fd_sc_hd__o41a_2
X_08185_ _08185_/A _08185_/B vssd1 vssd1 vccd1 vccd1 _08188_/A sky130_fd_sc_hd__nor2_1
X_07136_ _11929_/A _07136_/B vssd1 vssd1 vccd1 vccd1 _07136_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_70_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07067_ _09947_/A _07073_/B vssd1 vssd1 vccd1 vccd1 _07068_/B sky130_fd_sc_hd__or2_1
XANTENNA__07983__B _07983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06599__B _06944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10327__B2 _10276_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10327__A1 _10136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11725__S _11813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ _09708_/A _09863_/A _10004_/A _10137_/A vssd1 vssd1 vccd1 vccd1 _09708_/X
+ sky130_fd_sc_hd__or4_1
X_07969_ _07969_/A _07969_/B vssd1 vssd1 vccd1 vccd1 _07970_/C sky130_fd_sc_hd__nor2_1
X_10980_ _10980_/A _10980_/B _10980_/C vssd1 vssd1 vccd1 vccd1 _10981_/B sky130_fd_sc_hd__and3_1
XANTENNA__11827__A1 _11990_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout52_A _07079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09496__A2 fanout78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09639_ _09850_/B _09639_/B vssd1 vssd1 vccd1 vccd1 _09688_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_84_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12650_ reg1_val[2] _12650_/B vssd1 vssd1 vccd1 vccd1 _12651_/B sky130_fd_sc_hd__nand2_1
X_11601_ _11698_/A _11601_/B vssd1 vssd1 vccd1 vccd1 _11603_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_108_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12581_ _12598_/A _12581_/B vssd1 vssd1 vccd1 vccd1 _12597_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_108_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11532_ max_cap3/X _11122_/X _11527_/X _11531_/X vssd1 vssd1 vccd1 vccd1 _11533_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_52_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11463_ _11646_/B _11557_/B hold177/A vssd1 vssd1 vccd1 vccd1 _11463_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13202_ _13202_/A _13202_/B vssd1 vssd1 vccd1 vccd1 _13203_/B sky130_fd_sc_hd__nand2_1
X_10414_ _10538_/B _10414_/B vssd1 vssd1 vccd1 vccd1 _10415_/B sky130_fd_sc_hd__or2_4
X_11394_ _11395_/A _11395_/B vssd1 vssd1 vccd1 vccd1 _11396_/A sky130_fd_sc_hd__and2_1
XANTENNA__10566__A1 _11990_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13133_ _13133_/A _13133_/B vssd1 vssd1 vccd1 vccd1 _13134_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_61_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10345_ _10215_/A _10215_/B _10212_/A vssd1 vssd1 vccd1 vccd1 _10356_/A sky130_fd_sc_hd__o21bai_1
X_13064_ _13341_/Q _13094_/A2 _13101_/A2 hold130/X _13259_/A vssd1 vssd1 vccd1 vccd1
+ hold131/A sky130_fd_sc_hd__o221a_1
X_10276_ _10276_/A _10276_/B vssd1 vssd1 vccd1 vccd1 _10661_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__07982__A2 _07080_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12015_ _12336_/A _12015_/B vssd1 vssd1 vccd1 vccd1 _12024_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07117__C _07117_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap3 _10664_/B vssd1 vssd1 vccd1 vccd1 max_cap3/X sky130_fd_sc_hd__clkbuf_2
X_12917_ _13115_/A _13116_/A _13115_/B vssd1 vssd1 vccd1 vccd1 _13120_/B sky130_fd_sc_hd__a21bo_1
X_12848_ hold52/X _12862_/B vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__or2_1
XFILLER_0_75_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ _12790_/B _12779_/B vssd1 vssd1 vccd1 vccd1 _12782_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_126_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11754__B1 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09990_ _09991_/A _09991_/B vssd1 vssd1 vccd1 vccd1 _09990_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_12_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07422__B2 _07148_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07422__A1 _07554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08941_ _08940_/B _08941_/B vssd1 vssd1 vccd1 vccd1 _08942_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_110_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08872_ reg1_val[30] _08872_/B vssd1 vssd1 vccd1 vccd1 _08874_/B sky130_fd_sc_hd__xnor2_2
X_07823_ _07823_/A _07823_/B vssd1 vssd1 vccd1 vccd1 _07828_/A sky130_fd_sc_hd__xor2_2
XANTENNA__07725__A2 _07959_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout187_A _13257_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07754_ _07754_/A _07754_/B vssd1 vssd1 vccd1 vccd1 _07866_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06705_ _07078_/A reg1_val[19] vssd1 vssd1 vccd1 vccd1 _11652_/S sky130_fd_sc_hd__and2b_1
XFILLER_0_67_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11285__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07685_ _09943_/B2 fanout98/X fanout84/X _08538_/A1 vssd1 vssd1 vccd1 vccd1 _07686_/B
+ sky130_fd_sc_hd__o22a_1
X_06636_ _06634_/Y _06724_/B1 _06783_/A reg2_val[30] vssd1 vssd1 vccd1 vccd1 _08973_/C
+ sky130_fd_sc_hd__a2bb2o_4
X_09424_ hold245/A _09425_/C hold235/A vssd1 vssd1 vccd1 vccd1 _09424_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09355_ _09355_/A _09355_/B vssd1 vssd1 vccd1 vccd1 _09368_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_117_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10245__B1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08306_ _08306_/A _08306_/B vssd1 vssd1 vccd1 vccd1 _08352_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_7_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09286_ _09286_/A _09286_/B vssd1 vssd1 vccd1 vccd1 _09336_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08237_ _10207_/A _08237_/B vssd1 vssd1 vccd1 vccd1 _08314_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08168_ _08005_/A _08004_/B _08004_/C vssd1 vssd1 vccd1 vccd1 _08169_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_113_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07119_ _07215_/B _07133_/A _07133_/B _06827_/B vssd1 vssd1 vccd1 vccd1 _07121_/B
+ sky130_fd_sc_hd__a211o_1
X_08099_ _08099_/A _08099_/B vssd1 vssd1 vccd1 vccd1 _08155_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06767__A3 _12685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10130_ _10130_/A _10130_/B vssd1 vssd1 vccd1 vccd1 _10132_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10061_ _12009_/A fanout78/X fanout74/X fanout58/X vssd1 vssd1 vccd1 vccd1 _10062_/B
+ sky130_fd_sc_hd__o22a_1
X_10963_ _10963_/A _10963_/B vssd1 vssd1 vccd1 vccd1 _10966_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11276__A2 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12702_ reg1_val[12] _12702_/B vssd1 vssd1 vccd1 vccd1 _12703_/B sky130_fd_sc_hd__or2_1
X_10894_ _10894_/A _10894_/B vssd1 vssd1 vccd1 vccd1 _10897_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12633_ _12633_/A _12633_/B vssd1 vssd1 vccd1 vccd1 _12634_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_26_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12564_ _12719_/B _12564_/B vssd1 vssd1 vccd1 vccd1 _12565_/B sky130_fd_sc_hd__or2_1
XFILLER_0_93_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11515_ _11516_/B _11516_/A vssd1 vssd1 vccd1 vccd1 _11612_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_110_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12495_ _12504_/A _12495_/B vssd1 vssd1 vccd1 vccd1 _12497_/C sky130_fd_sc_hd__nand2_1
X_11446_ _06728_/B _11346_/X _06726_/X vssd1 vssd1 vccd1 vccd1 _11447_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_40_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11377_ _12050_/A _11567_/B _11893_/A vssd1 vssd1 vccd1 vccd1 _11377_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13116_ _13116_/A _13116_/B vssd1 vssd1 vccd1 vccd1 _13116_/Y sky130_fd_sc_hd__xnor2_1
X_10328_ _10276_/A _10276_/B _10327_/X vssd1 vssd1 vccd1 vccd1 _10328_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07409__A _07604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _07010_/B _12820_/B _13046_/X vssd1 vssd1 vccd1 vccd1 _13333_/D sky130_fd_sc_hd__a21oi_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ _10259_/A _10259_/B vssd1 vssd1 vccd1 vccd1 _10260_/B sky130_fd_sc_hd__nor2_2
XANTENNA__10711__A1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10711__B2 _11671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10172__C1 _12416_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12050__A _12050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10475__B1 _08411_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12985__A _13001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07470_ _07202_/Y _10337_/A _07238_/Y _07191_/X vssd1 vssd1 vccd1 vccd1 _07471_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07891__A1 _09934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07891__B2 _09822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09093__B1 _09301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09140_ _09141_/B _09141_/A vssd1 vssd1 vccd1 vccd1 _09140_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_16_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_210 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09071_ _09944_/A _09071_/B vssd1 vssd1 vccd1 vccd1 _09075_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08022_ _08094_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08095_/A sky130_fd_sc_hd__or2_1
XFILLER_0_97_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout5 fanout6/X vssd1 vssd1 vccd1 vccd1 fanout5/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_12_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09973_ _09973_/A _09973_/B vssd1 vssd1 vccd1 vccd1 _09976_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07319__A _09672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09148__A1 _10049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08924_ _09040_/A _09040_/B _09040_/C vssd1 vssd1 vccd1 vccd1 _08924_/X sky130_fd_sc_hd__and3_1
XANTENNA__12152__B1 _12631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10702__A1 _11752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08855_ _08943_/B _08855_/B vssd1 vssd1 vccd1 vccd1 _08868_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_98_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07806_ _07806_/A _07806_/B vssd1 vssd1 vccd1 vccd1 _07878_/A sky130_fd_sc_hd__xnor2_1
X_08786_ _08790_/A _08786_/B vssd1 vssd1 vccd1 vccd1 _08786_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07737_ _07737_/A _07737_/B _07737_/C vssd1 vssd1 vccd1 vccd1 _07739_/A sky130_fd_sc_hd__and3_1
XANTENNA__08123__A2 _08199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06893__A _06992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07668_ _07502_/A _07502_/B _07500_/Y vssd1 vssd1 vccd1 vccd1 _07669_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__07331__B1 _10240_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06619_ _06723_/A _12714_/B vssd1 vssd1 vccd1 vccd1 _06619_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_82_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09407_ _09399_/X _09406_/X _11138_/A vssd1 vssd1 vccd1 vccd1 _09407_/X sky130_fd_sc_hd__mux2_1
X_07599_ _07599_/A _07599_/B vssd1 vssd1 vccd1 vccd1 _07601_/C sky130_fd_sc_hd__xor2_1
X_09338_ _07830_/B _07198_/Y _10599_/A fanout46/X vssd1 vssd1 vccd1 vccd1 _09339_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_124_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout15_A fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11300_ _12096_/A _11300_/B vssd1 vssd1 vccd1 vccd1 _11301_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_90_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09269_ _09270_/B _09269_/B vssd1 vssd1 vccd1 vccd1 _09512_/A sky130_fd_sc_hd__and2b_1
X_12280_ _12335_/B _12235_/A _12234_/B _12233_/X vssd1 vssd1 vccd1 vccd1 _12292_/A
+ sky130_fd_sc_hd__o31a_1
XANTENNA__08613__A _08613_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11231_ _10283_/B _10780_/X _11229_/X _11230_/X vssd1 vssd1 vccd1 vccd1 _11232_/B
+ sky130_fd_sc_hd__a31o_2
XANTENNA__07229__A _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10581__C _10581_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11162_ _11158_/X _11161_/Y _11752_/S vssd1 vssd1 vccd1 vccd1 dest_val[14] sky130_fd_sc_hd__mux2_8
X_10113_ _10113_/A _10113_/B vssd1 vssd1 vccd1 vccd1 _10116_/A sky130_fd_sc_hd__nor2_2
X_11093_ _11093_/A _12087_/B vssd1 vssd1 vccd1 vccd1 _11094_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_101_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12143__A0 _09228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
X_10044_ curr_PC[3] curr_PC[4] _09762_/B curr_PC[5] vssd1 vssd1 vccd1 vccd1 _10044_/X
+ sky130_fd_sc_hd__a31o_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11995_ _11995_/A _11995_/B vssd1 vssd1 vccd1 vccd1 _11995_/Y sky130_fd_sc_hd__nand2_1
X_10946_ _10947_/A _10947_/B vssd1 vssd1 vccd1 vccd1 _11055_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07899__A _09341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10877_ _10877_/A _10877_/B vssd1 vssd1 vccd1 vccd1 _10878_/B sky130_fd_sc_hd__and2_1
XFILLER_0_42_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12616_ _12633_/A _12616_/B vssd1 vssd1 vccd1 vccd1 _12621_/D sky130_fd_sc_hd__xnor2_4
XFILLER_0_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12547_ _12553_/B _12547_/B vssd1 vssd1 vccd1 vccd1 new_PC[12] sky130_fd_sc_hd__and2_4
XFILLER_0_81_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11868__B _12335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_3 _11567_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12478_ reg1_val[3] curr_PC[3] _12520_/S vssd1 vssd1 vccd1 vccd1 _12480_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11429_ _11429_/A _11429_/B vssd1 vssd1 vccd1 vccd1 _11431_/C sky130_fd_sc_hd__xor2_2
XANTENNA__09378__A1 _10049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07389__B1 _10500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07139__A _09834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11884__A _11884_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10932__B2 _12446_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10932__A1 _09221_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06978__A _07262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06970_ _11138_/A _10297_/S _09728_/S _12808_/A vssd1 vssd1 vccd1 vccd1 _06970_/X
+ sky130_fd_sc_hd__and4_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11488__A2 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08640_ _08640_/A _08640_/B vssd1 vssd1 vccd1 vccd1 _08652_/A sky130_fd_sc_hd__xor2_2
XANTENNA__09550__B2 _09371_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08571_ _08585_/A _08585_/B vssd1 vssd1 vccd1 vccd1 _08571_/Y sky130_fd_sc_hd__nand2_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12988__A2 _13000_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07522_ _08564_/A _07522_/B vssd1 vssd1 vccd1 vccd1 _07526_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07453_ _07463_/B _07531_/A _07463_/A vssd1 vssd1 vccd1 vccd1 _07466_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_119_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07384_ _07384_/A _07384_/B vssd1 vssd1 vccd1 vccd1 _07468_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09123_ _08998_/A _08998_/B _08996_/X vssd1 vssd1 vccd1 vccd1 _09125_/B sky130_fd_sc_hd__o21ba_1
XANTENNA__12070__C1 _12376_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07616__A1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07616__B2 _09661_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09054_ _07121_/Y fanout42/X _07282_/Y _07417_/B vssd1 vssd1 vccd1 vccd1 _09055_/B
+ sky130_fd_sc_hd__a22o_1
X_08005_ _08005_/A _08169_/A vssd1 vssd1 vccd1 vccd1 _08016_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11176__B2 fanout28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11176__A1 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08041__A1 _08641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08041__B2 _08627_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09956_ _09957_/A _09957_/B vssd1 vssd1 vccd1 vccd1 _09956_/Y sky130_fd_sc_hd__nor2_1
X_09887_ _11820_/A _12446_/C1 _09221_/Y vssd1 vssd1 vccd1 vccd1 _09887_/X sky130_fd_sc_hd__a21o_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08907_ _08907_/A _08907_/B vssd1 vssd1 vccd1 vccd1 _08909_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__10687__B1 _12205_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08838_ _09944_/A _08838_/B vssd1 vssd1 vccd1 vccd1 _08840_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07552__B1 _07172_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08769_ _08769_/A _08769_/B vssd1 vssd1 vccd1 vccd1 _11630_/C sky130_fd_sc_hd__xor2_1
X_11780_ _11781_/A _11781_/B vssd1 vssd1 vccd1 vccd1 _11872_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_95_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10800_ _10800_/A _11820_/A _10798_/X vssd1 vssd1 vccd1 vccd1 _10800_/X sky130_fd_sc_hd__or3b_1
XANTENNA__07304__B1 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10731_ _11946_/B fanout32/X fanout30/X _07013_/X vssd1 vssd1 vccd1 vccd1 _10732_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12401_ _12398_/Y _12400_/X _09149_/Y vssd1 vssd1 vccd1 vccd1 _12401_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10662_ _10143_/A _10143_/B _10661_/X vssd1 vssd1 vccd1 vccd1 _10662_/Y sky130_fd_sc_hd__o21bai_2
XFILLER_0_35_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13381_ _13385_/CLK _13381_/D vssd1 vssd1 vccd1 vccd1 hold274/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10593_ _10593_/A _10593_/B vssd1 vssd1 vccd1 vccd1 _10612_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12332_ _08973_/B _06961_/X _12309_/X _12331_/X _12631_/S vssd1 vssd1 vccd1 vccd1
+ dest_val[28] sky130_fd_sc_hd__o221a_4
XFILLER_0_35_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12263_ _12259_/X _12262_/X _12064_/S vssd1 vssd1 vccd1 vccd1 _12263_/Y sky130_fd_sc_hd__o21ai_1
X_11214_ _11214_/A _11214_/B vssd1 vssd1 vccd1 vccd1 _11215_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_120_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12194_ reg1_val[26] curr_PC[26] vssd1 vssd1 vccd1 vccd1 _12195_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08032__B2 _08561_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08032__A1 _08561_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11145_ hold272/A _12271_/A1 _11255_/B _12376_/C1 vssd1 vssd1 vccd1 vccd1 _11146_/B
+ sky130_fd_sc_hd__a31o_1
X_11076_ _11076_/A _11076_/B vssd1 vssd1 vccd1 vccd1 _11077_/B sky130_fd_sc_hd__or2_1
XANTENNA__07791__B1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10027_ hold300/A _10166_/C _11538_/A vssd1 vssd1 vccd1 vccd1 _10028_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__08335__A2 _07195_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07543__B1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11978_ _06860_/A _11897_/X _06861_/Y _12359_/A vssd1 vssd1 vccd1 vccd1 _11978_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10929_ _07195_/A _12422_/A _10925_/X _10926_/Y _10928_/Y vssd1 vssd1 vccd1 vccd1
+ _10929_/X sky130_fd_sc_hd__a221o_1
XANTENNA__09835__A2 _07256_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07846__A1 _10338_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07141__B _11242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07846__B2 _08457_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09048__B1 fanout16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12355__B1 _11892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11158__A1 _12365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09810_ _09811_/A _09811_/B vssd1 vssd1 vccd1 vccd1 _09931_/B sky130_fd_sc_hd__and2_1
XANTENNA__08574__A2 _07134_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06953_ instruction[6] is_load vssd1 vssd1 vccd1 vccd1 _06953_/Y sky130_fd_sc_hd__nor2_1
X_09741_ _10165_/S _09740_/X _09251_/A vssd1 vssd1 vccd1 vccd1 _12319_/B sky130_fd_sc_hd__o21a_2
XANTENNA__09523__A1 _09325_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06884_ _06672_/D _06883_/X _06869_/X vssd1 vssd1 vccd1 vccd1 _06884_/X sky130_fd_sc_hd__a21o_1
X_09672_ _09672_/A _09672_/B vssd1 vssd1 vccd1 vccd1 _09673_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07316__B _10476_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10958__A _11929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08623_ _08603_/X _08621_/Y _08620_/Y _08611_/Y vssd1 vssd1 vccd1 vccd1 _08624_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout267_A _06783_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08554_ _08554_/A _08554_/B vssd1 vssd1 vccd1 vccd1 _08556_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09287__B1 _09650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07332__A _10749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07505_ _07505_/A _07505_/B vssd1 vssd1 vccd1 vccd1 _07571_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_92_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08485_ _08485_/A _08485_/B vssd1 vssd1 vccd1 vccd1 _08524_/B sky130_fd_sc_hd__xor2_1
XANTENNA__10841__B1 fanout45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07436_ _07440_/A _07440_/B vssd1 vssd1 vccd1 vccd1 _07436_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_9_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07367_ _07368_/A _07368_/B vssd1 vssd1 vccd1 vccd1 _07367_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_17_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11397__B2 _07032_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11397__A1 _06998_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09106_ _11946_/C _09106_/B vssd1 vssd1 vccd1 vccd1 _09108_/B sky130_fd_sc_hd__xnor2_2
X_07298_ _07298_/A _07298_/B vssd1 vssd1 vccd1 vccd1 _07298_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_60_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09037_ _09037_/A _09549_/A vssd1 vssd1 vccd1 vccd1 _09372_/B sky130_fd_sc_hd__or2_1
XFILLER_0_5_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09706__B _09707_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10372__A2 _08289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout82_A _10476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07773__B1 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09939_ _09939_/A _09939_/B vssd1 vssd1 vccd1 vccd1 _09942_/A sky130_fd_sc_hd__nand2_1
X_12950_ hold34/X hold274/A vssd1 vssd1 vccd1 vccd1 _13202_/B sky130_fd_sc_hd__nand2b_1
X_12881_ hold278/X hold64/X vssd1 vssd1 vccd1 vccd1 _13220_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11901_ reg1_val[22] curr_PC[22] vssd1 vssd1 vccd1 vccd1 _11903_/A sky130_fd_sc_hd__nand2_1
X_11832_ _10159_/A _10682_/X _10695_/Y _09222_/Y _11831_/X vssd1 vssd1 vccd1 vccd1
+ _11832_/X sky130_fd_sc_hd__o221a_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08338__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _11763_/A _11763_/B vssd1 vssd1 vccd1 vccd1 _11766_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12821__A1 _07282_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11694_ _11695_/A _11695_/B vssd1 vssd1 vccd1 vccd1 _11785_/B sky130_fd_sc_hd__and2_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _12096_/A _10714_/B vssd1 vssd1 vccd1 vccd1 _10715_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_126_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10645_ _10645_/A _10645_/B _10645_/C vssd1 vssd1 vccd1 vccd1 _10646_/B sky130_fd_sc_hd__or3_1
XFILLER_0_106_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13364_ _13365_/CLK _13364_/D vssd1 vssd1 vccd1 vccd1 hold256/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08253__A1 _08538_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10576_ _09221_/Y _10563_/X _10575_/X _12379_/B2 _10574_/Y vssd1 vssd1 vccd1 vccd1
+ _10576_/X sky130_fd_sc_hd__a221o_1
X_12315_ _12364_/A _09040_/A _08810_/B vssd1 vssd1 vccd1 vccd1 _12315_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09450__B1 _07238_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08253__B2 _08598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13295_ _13296_/CLK _13295_/D vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10108__A _11398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12246_ _12110_/Y _12178_/A _12178_/B vssd1 vssd1 vccd1 vccd1 _12246_/X sky130_fd_sc_hd__o21ba_1
X_12177_ _12177_/A _12177_/B _12177_/C vssd1 vssd1 vccd1 vccd1 _12178_/B sky130_fd_sc_hd__and3_1
XANTENNA__09753__A1 _11138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11128_ _11630_/A _11128_/B _08751_/A vssd1 vssd1 vccd1 vccd1 _11128_/X sky130_fd_sc_hd__or3b_1
XANTENNA__07764__B1 fanout72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07417__A _07959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11059_ _11060_/B _11060_/A vssd1 vssd1 vccd1 vccd1 _11207_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_64_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09632__A _09836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10666__A3 _11050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13065__A1 _10950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09808__A2 _08199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08248__A _08575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12993__A _13001_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08270_ _08270_/A _08270_/B vssd1 vssd1 vccd1 vccd1 _08327_/B sky130_fd_sc_hd__and2_1
XFILLER_0_116_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07221_ _07222_/A _07221_/B vssd1 vssd1 vccd1 vccd1 _07221_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_6_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07152_ reg1_val[24] _07585_/B1 _07167_/B reg1_val[25] vssd1 vssd1 vccd1 vccd1 _07155_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_27_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07083_ reg1_val[6] reg1_val[7] _07083_/C _07083_/D vssd1 vssd1 vccd1 vccd1 _07105_/D
+ sky130_fd_sc_hd__or4_2
XFILLER_0_112_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11548__S _12064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout104 _09479_/B1 vssd1 vssd1 vccd1 vccd1 _10240_/A sky130_fd_sc_hd__buf_6
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09744__A1 _12054_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12233__A _12233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout115 _07217_/Y vssd1 vssd1 vccd1 vccd1 _10221_/B2 sky130_fd_sc_hd__buf_8
Xfanout126 _07183_/X vssd1 vssd1 vccd1 vccd1 _11182_/A sky130_fd_sc_hd__clkbuf_8
Xfanout137 _10207_/A vssd1 vssd1 vccd1 vccd1 _10623_/A sky130_fd_sc_hd__buf_12
XANTENNA__07327__A _09944_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout148 _07068_/Y vssd1 vssd1 vccd1 vccd1 _09943_/B2 sky130_fd_sc_hd__buf_8
Xfanout159 _11892_/A vssd1 vssd1 vccd1 vccd1 _12364_/A sky130_fd_sc_hd__buf_4
X_07985_ _08664_/A _07985_/B _07985_/C vssd1 vssd1 vccd1 vccd1 _07988_/B sky130_fd_sc_hd__and3_1
X_06936_ instruction[26] _06944_/B vssd1 vssd1 vccd1 vccd1 _06936_/X sky130_fd_sc_hd__or2_1
X_09724_ _09720_/X _09723_/X _11246_/S vssd1 vssd1 vccd1 vccd1 _09724_/X sky130_fd_sc_hd__mux2_1
X_06867_ reg1_val[28] _06867_/B vssd1 vssd1 vccd1 vccd1 _06867_/Y sky130_fd_sc_hd__nand2_1
X_09655_ _09655_/A _09655_/B vssd1 vssd1 vccd1 vccd1 _09658_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_96_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08606_ _08677_/A _08677_/B vssd1 vssd1 vccd1 vccd1 _08678_/B sky130_fd_sc_hd__or2_1
X_06798_ _06815_/A _06817_/B1 _12660_/B _06797_/X vssd1 vssd1 vccd1 vccd1 _07166_/A
+ sky130_fd_sc_hd__a31oi_4
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ _09586_/A _09586_/B vssd1 vssd1 vccd1 vccd1 _09586_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08537_ _08543_/B _08543_/A vssd1 vssd1 vccd1 vccd1 _08537_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_108_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08468_ _08468_/A _08468_/B vssd1 vssd1 vccd1 vccd1 _08470_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07419_ _07420_/A _07420_/B vssd1 vssd1 vccd1 vccd1 _07425_/A sky130_fd_sc_hd__nor2_1
X_10430_ _09183_/X _09214_/X _11246_/S vssd1 vssd1 vccd1 vccd1 _10431_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_45_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08399_ _08399_/A _08399_/B vssd1 vssd1 vccd1 vccd1 _08431_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_122_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10042__A1 _09225_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_1_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10361_ _10362_/A _10362_/B vssd1 vssd1 vccd1 vccd1 _10363_/A sky130_fd_sc_hd__and2_1
XANTENNA__10042__B2 _12379_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12100_ _12101_/A _12101_/B _12101_/C vssd1 vssd1 vccd1 vccd1 _12102_/A sky130_fd_sc_hd__o21a_1
X_13080_ hold103/A _12805_/A _13250_/B hold89/X _13259_/A vssd1 vssd1 vccd1 vccd1
+ hold90/A sky130_fd_sc_hd__o221a_1
X_10292_ _11246_/S _09199_/X _11247_/C vssd1 vssd1 vccd1 vccd1 _10292_/X sky130_fd_sc_hd__o21a_1
Xhold180 hold180/A vssd1 vssd1 vccd1 vccd1 hold180/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12031_ _12108_/B _12031_/B vssd1 vssd1 vccd1 vccd1 _12033_/B sky130_fd_sc_hd__and2_1
XANTENNA__08538__A2 _08649_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold191 hold191/A vssd1 vssd1 vccd1 vccd1 hold191/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09499__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12933_ _13158_/A _13159_/A _13158_/B vssd1 vssd1 vccd1 vccd1 _13164_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__11845__A2 fanout41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10598__A _10599_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06795__B _07117_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12864_ hold58/X _12870_/B vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__or2_1
X_11815_ reg1_val[21] curr_PC[21] vssd1 vssd1 vccd1 vccd1 _11817_/A sky130_fd_sc_hd__nand2_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _12795_/A _12795_/B vssd1 vssd1 vccd1 vccd1 _12796_/B sky130_fd_sc_hd__xnor2_2
X_11746_ _11740_/Y _11741_/X _11745_/X vssd1 vssd1 vccd1 vccd1 _11747_/D sky130_fd_sc_hd__o21ai_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08474__A1 _08627_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07700__A _08575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08474__B2 _08641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11677_ _12336_/A _11677_/B vssd1 vssd1 vccd1 vccd1 _11681_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10628_ _12233_/B fanout75/X fanout17/X _08289_/B vssd1 vssd1 vccd1 vccd1 _10629_/B
+ sky130_fd_sc_hd__o22a_1
X_10559_ reg1_val[9] curr_PC[9] vssd1 vssd1 vccd1 vccd1 _10560_/B sky130_fd_sc_hd__nand2_1
X_13347_ _13354_/CLK _13347_/D vssd1 vssd1 vccd1 vccd1 hold133/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09974__A1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09974__B2 _11476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13278_ _13390_/CLK _13278_/D vssd1 vssd1 vccd1 vccd1 hold106/A sky130_fd_sc_hd__dfxtp_1
X_12229_ _12230_/A _12230_/B vssd1 vssd1 vccd1 vccd1 _12284_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08531__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07147__A _12359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12089__A2 _12335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11892__A _11892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07770_ _07781_/A _07781_/B vssd1 vssd1 vccd1 vccd1 _07770_/X sky130_fd_sc_hd__and2b_1
XANTENNA__06986__A _07036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06721_ _06719_/X _06721_/B vssd1 vssd1 vccd1 vccd1 _11449_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_91_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09440_ _09377_/Y _09378_/X _09439_/X vssd1 vssd1 vccd1 vccd1 _09440_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_94_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06652_ _12143_/S _06652_/B vssd1 vssd1 vccd1 vccd1 _06672_/A sky130_fd_sc_hd__or2_2
XANTENNA__13038__B2 _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06583_ reg1_val[31] vssd1 vssd1 vccd1 vccd1 _12795_/A sky130_fd_sc_hd__clkinv_4
X_09371_ _09371_/A _09371_/B vssd1 vssd1 vccd1 vccd1 _10004_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_86_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08322_ _08320_/A _08320_/B _08321_/X vssd1 vssd1 vccd1 vccd1 _08360_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08253_ _08538_/A1 _10221_/B2 _08501_/B1 _08598_/B vssd1 vssd1 vccd1 vccd1 _08254_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout132_A _07098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07204_ _11381_/A _07204_/B vssd1 vssd1 vccd1 vccd1 _07226_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09414__B1 _09242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08184_ _08087_/A _08086_/B _08086_/C vssd1 vssd1 vccd1 vccd1 _08185_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_113_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07135_ _08613_/B _08613_/C vssd1 vssd1 vccd1 vccd1 _07135_/X sky130_fd_sc_hd__or2_1
X_07066_ _09947_/A _07073_/B vssd1 vssd1 vccd1 vccd1 _10072_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08441__A _08564_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10327__A2 _10136_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10910__S _11813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ _07968_/A _07968_/B vssd1 vssd1 vccd1 vccd1 _07969_/B sky130_fd_sc_hd__and2_1
X_06919_ _06783_/A _06610_/X _09239_/B instruction[4] _06917_/Y vssd1 vssd1 vccd1
+ vccd1 _12804_/B sky130_fd_sc_hd__a221o_1
X_09707_ _09707_/A _09707_/B vssd1 vssd1 vccd1 vccd1 _10137_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_4_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07899_ _09341_/A _07899_/B vssd1 vssd1 vccd1 vccd1 _08000_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11307__A _12017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout45_A fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09638_ _09638_/A _09638_/B vssd1 vssd1 vccd1 vccd1 _09639_/B sky130_fd_sc_hd__or2_1
XFILLER_0_78_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09569_ _09565_/X _09568_/X _11246_/S vssd1 vssd1 vccd1 vccd1 _09569_/X sky130_fd_sc_hd__mux2_1
X_11600_ _11600_/A _11600_/B _11598_/Y vssd1 vssd1 vccd1 vccd1 _11601_/B sky130_fd_sc_hd__or3b_1
X_12580_ _12633_/A _12580_/B vssd1 vssd1 vccd1 vccd1 _12581_/B sky130_fd_sc_hd__or2_1
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06649__A2_N _06766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11531_ _11121_/X _11527_/X _11530_/X vssd1 vssd1 vccd1 vccd1 _11531_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07520__A _09947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11462_ hold177/A _11646_/B _11557_/B vssd1 vssd1 vccd1 vccd1 _11462_/X sky130_fd_sc_hd__and3_1
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13201_ _13210_/A _13201_/B vssd1 vssd1 vccd1 vccd1 _13381_/D sky130_fd_sc_hd__and2_1
X_11393_ _11393_/A _11393_/B vssd1 vssd1 vccd1 vccd1 _11395_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10413_ _10413_/A _10413_/B _10413_/C vssd1 vssd1 vccd1 vccd1 _10414_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_33_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10344_ _10468_/B _10344_/B vssd1 vssd1 vccd1 vccd1 _10368_/A sky130_fd_sc_hd__and2_1
X_13132_ _13147_/A hold261/X vssd1 vssd1 vccd1 vccd1 _13367_/D sky130_fd_sc_hd__and2_1
XFILLER_0_21_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10275_ _10275_/A _10275_/B vssd1 vssd1 vccd1 vccd1 _10276_/B sky130_fd_sc_hd__xnor2_4
X_13063_ _07254_/B _12826_/B hold83/X vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12014_ fanout17/X fanout23/X fanout15/X _12233_/B vssd1 vssd1 vccd1 vccd1 _12015_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap4 _10004_/Y vssd1 vssd1 vccd1 vccd1 max_cap4/X sky130_fd_sc_hd__buf_1
XANTENNA__08144__B1 _09479_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12916_ hold92/X hold295/A vssd1 vssd1 vccd1 vccd1 _13115_/B sky130_fd_sc_hd__nand2b_1
X_12847_ _11592_/A _12863_/A2 hold97/X _13019_/A vssd1 vssd1 vccd1 vccd1 _13284_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09910__A _10049_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _12787_/A _12778_/B vssd1 vssd1 vccd1 vccd1 _12782_/A sky130_fd_sc_hd__or2_1
XFILLER_0_29_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11729_ reg1_val[20] curr_PC[20] vssd1 vssd1 vccd1 vccd1 _11730_/B sky130_fd_sc_hd__or2_1
XFILLER_0_83_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10791__A _11813_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11754__A1 _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11754__B2 _12009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07422__A2 _07173_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11506__A1 _11406_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08940_ _08941_/B _08940_/B vssd1 vssd1 vccd1 vccd1 _08942_/A sky130_fd_sc_hd__and2b_1
X_08871_ reg1_val[28] reg1_val[29] _08870_/C _12779_/B _07248_/A vssd1 vssd1 vccd1
+ vccd1 _08872_/B sky130_fd_sc_hd__o41a_1
XANTENNA__07186__A1 _11134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07822_ _07822_/A _07822_/B vssd1 vssd1 vccd1 vccd1 _07872_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09092__A _09673_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07753_ _07754_/A _07754_/B vssd1 vssd1 vccd1 vccd1 _07753_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06704_ reg2_val[19] _06766_/B _06724_/B1 _06703_/Y vssd1 vssd1 vccd1 vccd1 _07078_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07684_ _08454_/A _07684_/B vssd1 vssd1 vccd1 vccd1 _07688_/A sky130_fd_sc_hd__xnor2_2
X_09423_ hold9/A _12359_/A vssd1 vssd1 vccd1 vccd1 _09423_/X sky130_fd_sc_hd__and2_1
X_06635_ reg2_val[30] _06783_/A _06724_/B1 _06634_/Y vssd1 vssd1 vccd1 vccd1 _08860_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_09354_ _09354_/A _09354_/B vssd1 vssd1 vccd1 vccd1 _09355_/B sky130_fd_sc_hd__and2_1
XANTENNA__10245__A1 _10245_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08305_ _08580_/A _08305_/B vssd1 vssd1 vccd1 vccd1 _08306_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_90_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08989__A2 _12428_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07110__A1 _11134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10245__B2 _10245_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11442__B1 _12356_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09285_ _09286_/A _09286_/B vssd1 vssd1 vccd1 vccd1 _09285_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_117_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08236_ _08576_/A2 _08411_/B _10476_/A _09472_/A vssd1 vssd1 vccd1 vccd1 _08237_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08167_ _08165_/A _08165_/B _08166_/Y vssd1 vssd1 vccd1 vccd1 _08177_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__11745__A1 _10159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11745__B2 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07118_ _11029_/S _06970_/X _06969_/Y _06972_/C vssd1 vssd1 vccd1 vccd1 _07121_/A
+ sky130_fd_sc_hd__a211o_1
X_08098_ _08098_/A _08098_/B vssd1 vssd1 vccd1 vccd1 _08155_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07049_ _07049_/A _07215_/B vssd1 vssd1 vccd1 vccd1 _07049_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__06621__B1 _06766_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10060_ _10060_/A _10060_/B vssd1 vssd1 vccd1 vccd1 _10065_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08126__B1 fanout80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10962_ _10962_/A _10962_/B vssd1 vssd1 vccd1 vccd1 _10963_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_85_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12701_ reg1_val[12] _12702_/B vssd1 vssd1 vccd1 vccd1 _12711_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_97_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10893_ _10894_/A _10894_/B vssd1 vssd1 vccd1 vccd1 _11006_/B sky130_fd_sc_hd__nand2_1
X_12632_ _12633_/A _12633_/B vssd1 vssd1 vccd1 vccd1 _12634_/A sky130_fd_sc_hd__and2_1
XANTENNA__07250__A _10749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12563_ _12719_/B _12564_/B vssd1 vssd1 vccd1 vccd1 _12572_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_93_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11514_ _11514_/A _11514_/B vssd1 vssd1 vccd1 vccd1 _11516_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12494_ _12665_/B _12494_/B vssd1 vssd1 vccd1 vccd1 _12495_/B sky130_fd_sc_hd__or2_1
XFILLER_0_81_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11445_ _11630_/A _11444_/B _11444_/C vssd1 vssd1 vccd1 vccd1 _11445_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_111_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11376_ _11374_/Y _11564_/B _11752_/S vssd1 vssd1 vccd1 vccd1 _11471_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_0_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13115_ _13115_/A _13115_/B vssd1 vssd1 vccd1 vccd1 _13116_/B sky130_fd_sc_hd__nand2_1
X_10327_ _10136_/A _10136_/B _10276_/A _10276_/B vssd1 vssd1 vccd1 vccd1 _10327_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10258_ _10257_/B _10257_/C _10257_/A vssd1 vssd1 vccd1 vccd1 _10259_/B sky130_fd_sc_hd__a21oi_1
X_13046_ hold39/X _06577_/A _13254_/A2 hold43/X rst vssd1 vssd1 vccd1 vccd1 _13046_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10711__A2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10189_ _10130_/A _10130_/B _10131_/X vssd1 vssd1 vccd1 vccd1 _10275_/A sky130_fd_sc_hd__o21bai_4
XANTENNA__10475__A1 _07608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13162__A _13162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07891__A2 _08199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09093__B2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09093__A1 _09669_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09070_ fanout68/X _07068_/Y _09650_/A fanout65/X vssd1 vssd1 vccd1 vccd1 _09071_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08021_ _08564_/A _08021_/B vssd1 vssd1 vccd1 vccd1 _08094_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout6 fanout6/A vssd1 vssd1 vccd1 vccd1 fanout6/X sky130_fd_sc_hd__buf_4
XANTENNA__09087__A _09667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09972_ _09973_/A _09973_/B vssd1 vssd1 vccd1 vccd1 _09972_/X sky130_fd_sc_hd__and2_1
XFILLER_0_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08923_ _09549_/A _10138_/A vssd1 vssd1 vccd1 vccd1 _09040_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_110_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08854_ _08854_/A _08854_/B vssd1 vssd1 vccd1 vccd1 _08855_/B sky130_fd_sc_hd__nand2_1
X_07805_ _07805_/A _07805_/B vssd1 vssd1 vccd1 vccd1 _07807_/B sky130_fd_sc_hd__xnor2_1
X_08785_ _08183_/X _08776_/B _08697_/X vssd1 vssd1 vccd1 vccd1 _08786_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__13101__B1 _11946_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07736_ _07537_/A _07537_/C _07537_/B vssd1 vssd1 vccd1 vccd1 _07737_/C sky130_fd_sc_hd__a21o_1
XANTENNA__11663__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06893__B _12808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07331__B2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07331__A1 _09661_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07667_ _07667_/A _07667_/B vssd1 vssd1 vccd1 vccd1 _07669_/A sky130_fd_sc_hd__xnor2_4
X_06618_ instruction[39] _06675_/B vssd1 vssd1 vccd1 vccd1 _12714_/B sky130_fd_sc_hd__and2_4
X_09406_ _09402_/X _10022_/B _10294_/S vssd1 vssd1 vccd1 vccd1 _09406_/X sky130_fd_sc_hd__mux2_1
X_07598_ _11844_/A _07598_/B vssd1 vssd1 vccd1 vccd1 _07599_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09337_ _09050_/Y _09053_/B _09058_/A vssd1 vssd1 vccd1 vccd1 _09351_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_63_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09268_ _09922_/A _09268_/B vssd1 vssd1 vccd1 vccd1 _09269_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08219_ _08222_/A _08222_/B vssd1 vssd1 vccd1 vccd1 _08219_/X sky130_fd_sc_hd__and2b_1
X_09199_ _09191_/X _09198_/X _10295_/S vssd1 vssd1 vccd1 vccd1 _09199_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11230_ _10782_/X _11229_/X _11623_/A vssd1 vssd1 vccd1 vccd1 _11230_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_30_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11161_ _11268_/B _11161_/B vssd1 vssd1 vccd1 vccd1 _11161_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10112_ _10112_/A _10112_/B vssd1 vssd1 vccd1 vccd1 _10113_/B sky130_fd_sc_hd__nor2_1
X_11092_ _12336_/A _11092_/B vssd1 vssd1 vccd1 vccd1 _11094_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
X_10043_ _12365_/A _10009_/Y _10010_/X _10042_/X _10008_/Y vssd1 vssd1 vccd1 vccd1
+ _10043_/X sky130_fd_sc_hd__a311o_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
X_11994_ hold254/A _12271_/A1 _12068_/B _11993_/Y _12376_/C1 vssd1 vssd1 vccd1 vccd1
+ _11994_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_98_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10945_ _12224_/A _10945_/B vssd1 vssd1 vccd1 vccd1 _10947_/B sky130_fd_sc_hd__xor2_1
X_10876_ _10877_/A _10877_/B vssd1 vssd1 vccd1 vccd1 _10878_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12615_ reg1_val[23] curr_PC[23] _12638_/S vssd1 vssd1 vccd1 vccd1 _12616_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12546_ _12546_/A _12546_/B _12546_/C vssd1 vssd1 vccd1 vccd1 _12547_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_53_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12477_ _12483_/B _12477_/B vssd1 vssd1 vccd1 vccd1 new_PC[2] sky130_fd_sc_hd__and2_4
X_11428_ _11429_/A _11429_/B vssd1 vssd1 vccd1 vccd1 _11524_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_4 instruction[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11359_ _11359_/A _11359_/B vssd1 vssd1 vccd1 vccd1 _11359_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07389__A1 _08199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07389__B2 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06978__B _07270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ _13162_/A hold225/X vssd1 vssd1 vccd1 vccd1 hold226/A sky130_fd_sc_hd__and2_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10696__B2 _10159_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10696__A1 _09222_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09550__A2 _09146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08570_ _08594_/A _08570_/B vssd1 vssd1 vccd1 vccd1 _08585_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09370__A _09371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07521_ _08540_/B fanout84/X fanout80/X _08515_/A2 vssd1 vssd1 vccd1 vccd1 _07522_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11405__A _12336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07452_ _07530_/A _07530_/B vssd1 vssd1 vccd1 vccd1 _07531_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_9_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07383_ _10623_/A _07383_/B vssd1 vssd1 vccd1 vccd1 _07468_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07077__B1 _07078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09122_ _09122_/A _09122_/B vssd1 vssd1 vccd1 vccd1 _09125_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_32_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07616__A2 _10473_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09053_ _09053_/A _09053_/B vssd1 vssd1 vccd1 vccd1 _09057_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_102_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08004_ _08005_/A _08004_/B _08004_/C vssd1 vssd1 vccd1 vccd1 _08169_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_12_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11176__A2 fanout17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap240 _09671_/A vssd1 vssd1 vccd1 vccd1 _08656_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_6_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10384__B1 fanout34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10923__A2 _11990_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08041__A2 fanout76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09955_ _11179_/A _09955_/B vssd1 vssd1 vccd1 vccd1 _09957_/B sky130_fd_sc_hd__xnor2_4
X_09886_ _09883_/X _09885_/X _11247_/A vssd1 vssd1 vccd1 vccd1 _09886_/X sky130_fd_sc_hd__mux2_2
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08906_ _08906_/A _08906_/B vssd1 vssd1 vccd1 vccd1 _08907_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_99_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08837_ fanout59/X _09943_/B2 _09650_/A fanout57/X vssd1 vssd1 vccd1 vccd1 _08838_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07552__B2 _07830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07552__A1 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08768_ _08769_/A _08769_/B vssd1 vssd1 vccd1 vccd1 _08768_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__12833__C1 _13162_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07719_ _08334_/A _07719_/B vssd1 vssd1 vccd1 vccd1 _07755_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07304__A1 fanout86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08699_ _08077_/X _08183_/X _08776_/B _08696_/Y _08698_/X vssd1 vssd1 vccd1 vccd1
+ _08711_/B sky130_fd_sc_hd__o311a_2
XFILLER_0_95_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10730_ _11182_/A _10730_/B vssd1 vssd1 vccd1 vccd1 _10734_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07304__B2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08501__B1 _08501_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10661_ _10661_/A _10661_/B _10661_/C _10779_/A vssd1 vssd1 vccd1 vccd1 _10661_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_125_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12400_ _12050_/X _12306_/X _12399_/X _11892_/A vssd1 vssd1 vccd1 vccd1 _12400_/X
+ sky130_fd_sc_hd__a31o_1
X_13380_ _13385_/CLK _13380_/D vssd1 vssd1 vccd1 vccd1 hold262/A sky130_fd_sc_hd__dfxtp_1
X_10592_ _10591_/B _10592_/B vssd1 vssd1 vccd1 vccd1 _10593_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_8_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12331_ _12331_/A _12331_/B _12331_/C _12330_/X vssd1 vssd1 vccd1 vccd1 _12331_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_63_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12262_ _12260_/Y _12262_/B vssd1 vssd1 vccd1 vccd1 _12262_/X sky130_fd_sc_hd__and2b_1
XANTENNA__11050__A _11050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11213_ _11214_/B vssd1 vssd1 vccd1 vccd1 _11213_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_121_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12193_ reg1_val[26] curr_PC[26] vssd1 vssd1 vccd1 vccd1 _12193_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08032__A2 _08289_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11144_ _12271_/A1 _11255_/B hold272/A vssd1 vssd1 vccd1 vccd1 _11146_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11075_ _11076_/A _11076_/B vssd1 vssd1 vccd1 vccd1 _11194_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07791__A1 _07217_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07791__B2 _07221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10026_ _10165_/S _10025_/Y _10021_/X vssd1 vssd1 vccd1 vccd1 _10026_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07543__B2 _07166_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07543__A1 _07134_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12419__A2 _12447_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11977_ _11977_/A _11977_/B vssd1 vssd1 vccd1 vccd1 _11977_/X sky130_fd_sc_hd__or2_2
X_10928_ _12144_/A1 _10927_/X _06748_/B vssd1 vssd1 vccd1 vccd1 _10928_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07846__A2 _08484_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10859_ _11309_/A _07362_/B fanout16/X _11198_/A vssd1 vssd1 vccd1 vccd1 _10860_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09048__A1 _09822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09048__B2 _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12052__B1 _09149_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09599__A2 _12420_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08534__A _08575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12529_ _12689_/B _12529_/B vssd1 vssd1 vccd1 vccd1 _12530_/B sky130_fd_sc_hd__or2_1
XFILLER_0_14_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08559__B1 _09940_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09220__A1 _12064_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10905__A2 _11050_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06952_ instruction[17] _09242_/B _09221_/B _06783_/A vssd1 vssd1 vccd1 vccd1 _06952_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_94_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09740_ _11246_/S _09739_/X _11247_/C vssd1 vssd1 vccd1 vccd1 _09740_/X sky130_fd_sc_hd__o21a_1
.ends

