magic
tech sky130B
magscale 1 2
timestamp 1716925469
<< obsli1 >>
rect 1104 2159 218868 147441
<< obsm1 >>
rect 750 348 218928 147472
<< metal2 >>
rect 3698 149200 3754 150000
rect 9770 149200 9826 150000
rect 15842 149200 15898 150000
rect 21914 149200 21970 150000
rect 27986 149200 28042 150000
rect 34058 149200 34114 150000
rect 40130 149200 40186 150000
rect 46202 149200 46258 150000
rect 52274 149200 52330 150000
rect 58346 149200 58402 150000
rect 64418 149200 64474 150000
rect 70490 149200 70546 150000
rect 76562 149200 76618 150000
rect 82634 149200 82690 150000
rect 88706 149200 88762 150000
rect 94778 149200 94834 150000
rect 100850 149200 100906 150000
rect 106922 149200 106978 150000
rect 112994 149200 113050 150000
rect 119066 149200 119122 150000
rect 125138 149200 125194 150000
rect 131210 149200 131266 150000
rect 137282 149200 137338 150000
rect 143354 149200 143410 150000
rect 149426 149200 149482 150000
rect 155498 149200 155554 150000
rect 161570 149200 161626 150000
rect 167642 149200 167698 150000
rect 173714 149200 173770 150000
rect 179786 149200 179842 150000
rect 185858 149200 185914 150000
rect 191930 149200 191986 150000
rect 198002 149200 198058 150000
rect 204074 149200 204130 150000
rect 210146 149200 210202 150000
rect 216218 149200 216274 150000
rect 3698 0 3754 800
rect 9770 0 9826 800
rect 15842 0 15898 800
rect 21914 0 21970 800
rect 27986 0 28042 800
rect 34058 0 34114 800
rect 40130 0 40186 800
rect 46202 0 46258 800
rect 52274 0 52330 800
rect 58346 0 58402 800
rect 64418 0 64474 800
rect 70490 0 70546 800
rect 76562 0 76618 800
rect 82634 0 82690 800
rect 88706 0 88762 800
rect 94778 0 94834 800
rect 100850 0 100906 800
rect 106922 0 106978 800
rect 112994 0 113050 800
rect 119066 0 119122 800
rect 125138 0 125194 800
rect 131210 0 131266 800
rect 137282 0 137338 800
rect 143354 0 143410 800
rect 149426 0 149482 800
rect 155498 0 155554 800
rect 161570 0 161626 800
rect 167642 0 167698 800
rect 173714 0 173770 800
rect 179786 0 179842 800
rect 185858 0 185914 800
rect 191930 0 191986 800
rect 198002 0 198058 800
rect 204074 0 204130 800
rect 210146 0 210202 800
rect 216218 0 216274 800
<< obsm2 >>
rect 756 149144 3642 149200
rect 3810 149144 9714 149200
rect 9882 149144 15786 149200
rect 15954 149144 21858 149200
rect 22026 149144 27930 149200
rect 28098 149144 34002 149200
rect 34170 149144 40074 149200
rect 40242 149144 46146 149200
rect 46314 149144 52218 149200
rect 52386 149144 58290 149200
rect 58458 149144 64362 149200
rect 64530 149144 70434 149200
rect 70602 149144 76506 149200
rect 76674 149144 82578 149200
rect 82746 149144 88650 149200
rect 88818 149144 94722 149200
rect 94890 149144 100794 149200
rect 100962 149144 106866 149200
rect 107034 149144 112938 149200
rect 113106 149144 119010 149200
rect 119178 149144 125082 149200
rect 125250 149144 131154 149200
rect 131322 149144 137226 149200
rect 137394 149144 143298 149200
rect 143466 149144 149370 149200
rect 149538 149144 155442 149200
rect 155610 149144 161514 149200
rect 161682 149144 167586 149200
rect 167754 149144 173658 149200
rect 173826 149144 179730 149200
rect 179898 149144 185802 149200
rect 185970 149144 191874 149200
rect 192042 149144 197946 149200
rect 198114 149144 204018 149200
rect 204186 149144 210090 149200
rect 210258 149144 216162 149200
rect 216330 149144 218850 149200
rect 756 856 218850 149144
rect 756 342 3642 856
rect 3810 342 9714 856
rect 9882 342 15786 856
rect 15954 342 21858 856
rect 22026 342 27930 856
rect 28098 342 34002 856
rect 34170 342 40074 856
rect 40242 342 46146 856
rect 46314 342 52218 856
rect 52386 342 58290 856
rect 58458 342 64362 856
rect 64530 342 70434 856
rect 70602 342 76506 856
rect 76674 342 82578 856
rect 82746 342 88650 856
rect 88818 342 94722 856
rect 94890 342 100794 856
rect 100962 342 106866 856
rect 107034 342 112938 856
rect 113106 342 119010 856
rect 119178 342 125082 856
rect 125250 342 131154 856
rect 131322 342 137226 856
rect 137394 342 143298 856
rect 143466 342 149370 856
rect 149538 342 155442 856
rect 155610 342 161514 856
rect 161682 342 167586 856
rect 167754 342 173658 856
rect 173826 342 179730 856
rect 179898 342 185802 856
rect 185970 342 191874 856
rect 192042 342 197946 856
rect 198114 342 204018 856
rect 204186 342 210090 856
rect 210258 342 216162 856
rect 216330 342 218850 856
<< metal3 >>
rect 0 146616 800 146736
rect 219200 146344 220000 146464
rect 0 142264 800 142384
rect 219200 142264 220000 142384
rect 219200 138184 220000 138304
rect 0 137912 800 138032
rect 219200 134104 220000 134224
rect 0 133560 800 133680
rect 219200 130024 220000 130144
rect 0 129208 800 129328
rect 219200 125944 220000 126064
rect 0 124856 800 124976
rect 219200 121864 220000 121984
rect 0 120504 800 120624
rect 219200 117784 220000 117904
rect 0 116152 800 116272
rect 219200 113704 220000 113824
rect 0 111800 800 111920
rect 219200 109624 220000 109744
rect 0 107448 800 107568
rect 219200 105544 220000 105664
rect 0 103096 800 103216
rect 219200 101464 220000 101584
rect 0 98744 800 98864
rect 219200 97384 220000 97504
rect 0 94392 800 94512
rect 219200 93304 220000 93424
rect 0 90040 800 90160
rect 219200 89224 220000 89344
rect 0 85688 800 85808
rect 219200 85144 220000 85264
rect 0 81336 800 81456
rect 219200 81064 220000 81184
rect 0 76984 800 77104
rect 219200 76984 220000 77104
rect 219200 72904 220000 73024
rect 0 72632 800 72752
rect 219200 68824 220000 68944
rect 0 68280 800 68400
rect 219200 64744 220000 64864
rect 0 63928 800 64048
rect 219200 60664 220000 60784
rect 0 59576 800 59696
rect 219200 56584 220000 56704
rect 0 55224 800 55344
rect 219200 52504 220000 52624
rect 0 50872 800 50992
rect 219200 48424 220000 48544
rect 0 46520 800 46640
rect 219200 44344 220000 44464
rect 0 42168 800 42288
rect 219200 40264 220000 40384
rect 0 37816 800 37936
rect 219200 36184 220000 36304
rect 0 33464 800 33584
rect 219200 32104 220000 32224
rect 0 29112 800 29232
rect 219200 28024 220000 28144
rect 0 24760 800 24880
rect 219200 23944 220000 24064
rect 0 20408 800 20528
rect 219200 19864 220000 19984
rect 0 16056 800 16176
rect 219200 15784 220000 15904
rect 0 11704 800 11824
rect 219200 11704 220000 11824
rect 219200 7624 220000 7744
rect 0 7352 800 7472
rect 219200 3544 220000 3664
rect 0 3000 800 3120
<< obsm3 >>
rect 798 146816 219200 147457
rect 880 146544 219200 146816
rect 880 146536 219120 146544
rect 798 146264 219120 146536
rect 798 142464 219200 146264
rect 880 142184 219120 142464
rect 798 138384 219200 142184
rect 798 138112 219120 138384
rect 880 138104 219120 138112
rect 880 137832 219200 138104
rect 798 134304 219200 137832
rect 798 134024 219120 134304
rect 798 133760 219200 134024
rect 880 133480 219200 133760
rect 798 130224 219200 133480
rect 798 129944 219120 130224
rect 798 129408 219200 129944
rect 880 129128 219200 129408
rect 798 126144 219200 129128
rect 798 125864 219120 126144
rect 798 125056 219200 125864
rect 880 124776 219200 125056
rect 798 122064 219200 124776
rect 798 121784 219120 122064
rect 798 120704 219200 121784
rect 880 120424 219200 120704
rect 798 117984 219200 120424
rect 798 117704 219120 117984
rect 798 116352 219200 117704
rect 880 116072 219200 116352
rect 798 113904 219200 116072
rect 798 113624 219120 113904
rect 798 112000 219200 113624
rect 880 111720 219200 112000
rect 798 109824 219200 111720
rect 798 109544 219120 109824
rect 798 107648 219200 109544
rect 880 107368 219200 107648
rect 798 105744 219200 107368
rect 798 105464 219120 105744
rect 798 103296 219200 105464
rect 880 103016 219200 103296
rect 798 101664 219200 103016
rect 798 101384 219120 101664
rect 798 98944 219200 101384
rect 880 98664 219200 98944
rect 798 97584 219200 98664
rect 798 97304 219120 97584
rect 798 94592 219200 97304
rect 880 94312 219200 94592
rect 798 93504 219200 94312
rect 798 93224 219120 93504
rect 798 90240 219200 93224
rect 880 89960 219200 90240
rect 798 89424 219200 89960
rect 798 89144 219120 89424
rect 798 85888 219200 89144
rect 880 85608 219200 85888
rect 798 85344 219200 85608
rect 798 85064 219120 85344
rect 798 81536 219200 85064
rect 880 81264 219200 81536
rect 880 81256 219120 81264
rect 798 80984 219120 81256
rect 798 77184 219200 80984
rect 880 76904 219120 77184
rect 798 73104 219200 76904
rect 798 72832 219120 73104
rect 880 72824 219120 72832
rect 880 72552 219200 72824
rect 798 69024 219200 72552
rect 798 68744 219120 69024
rect 798 68480 219200 68744
rect 880 68200 219200 68480
rect 798 64944 219200 68200
rect 798 64664 219120 64944
rect 798 64128 219200 64664
rect 880 63848 219200 64128
rect 798 60864 219200 63848
rect 798 60584 219120 60864
rect 798 59776 219200 60584
rect 880 59496 219200 59776
rect 798 56784 219200 59496
rect 798 56504 219120 56784
rect 798 55424 219200 56504
rect 880 55144 219200 55424
rect 798 52704 219200 55144
rect 798 52424 219120 52704
rect 798 51072 219200 52424
rect 880 50792 219200 51072
rect 798 48624 219200 50792
rect 798 48344 219120 48624
rect 798 46720 219200 48344
rect 880 46440 219200 46720
rect 798 44544 219200 46440
rect 798 44264 219120 44544
rect 798 42368 219200 44264
rect 880 42088 219200 42368
rect 798 40464 219200 42088
rect 798 40184 219120 40464
rect 798 38016 219200 40184
rect 880 37736 219200 38016
rect 798 36384 219200 37736
rect 798 36104 219120 36384
rect 798 33664 219200 36104
rect 880 33384 219200 33664
rect 798 32304 219200 33384
rect 798 32024 219120 32304
rect 798 29312 219200 32024
rect 880 29032 219200 29312
rect 798 28224 219200 29032
rect 798 27944 219120 28224
rect 798 24960 219200 27944
rect 880 24680 219200 24960
rect 798 24144 219200 24680
rect 798 23864 219120 24144
rect 798 20608 219200 23864
rect 880 20328 219200 20608
rect 798 20064 219200 20328
rect 798 19784 219120 20064
rect 798 16256 219200 19784
rect 880 15984 219200 16256
rect 880 15976 219120 15984
rect 798 15704 219120 15976
rect 798 11904 219200 15704
rect 880 11624 219120 11904
rect 798 7824 219200 11624
rect 798 7552 219120 7824
rect 880 7544 219120 7552
rect 880 7272 219200 7544
rect 798 3744 219200 7272
rect 798 3464 219120 3744
rect 798 3200 219200 3464
rect 880 2920 219200 3200
rect 798 444 219200 2920
<< metal4 >>
rect 4208 2128 4528 147472
rect 19568 2128 19888 147472
rect 34928 2128 35248 147472
rect 50288 2128 50608 147472
rect 65648 2128 65968 147472
rect 81008 2128 81328 147472
rect 96368 2128 96688 147472
rect 111728 2128 112048 147472
rect 127088 2128 127408 147472
rect 142448 2128 142768 147472
rect 157808 2128 158128 147472
rect 173168 2128 173488 147472
rect 188528 2128 188848 147472
rect 203888 2128 204208 147472
<< obsm4 >>
rect 2635 2048 4128 147117
rect 4608 2048 19488 147117
rect 19968 2048 34848 147117
rect 35328 2048 50208 147117
rect 50688 2048 65568 147117
rect 66048 2048 80928 147117
rect 81408 2048 96288 147117
rect 96768 2048 111648 147117
rect 112128 2048 127008 147117
rect 127488 2048 142368 147117
rect 142848 2048 157728 147117
rect 158208 2048 173088 147117
rect 173568 2048 188448 147117
rect 188928 2048 203808 147117
rect 204288 2048 217245 147117
rect 2635 443 217245 2048
<< labels >>
rlabel metal3 s 0 11704 800 11824 6 custom_settings[0]
port 1 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 custom_settings[10]
port 2 nsew signal input
rlabel metal3 s 0 59576 800 59696 6 custom_settings[11]
port 3 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 custom_settings[12]
port 4 nsew signal input
rlabel metal3 s 0 68280 800 68400 6 custom_settings[13]
port 5 nsew signal input
rlabel metal3 s 0 72632 800 72752 6 custom_settings[14]
port 6 nsew signal input
rlabel metal3 s 0 76984 800 77104 6 custom_settings[15]
port 7 nsew signal input
rlabel metal3 s 0 81336 800 81456 6 custom_settings[16]
port 8 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 custom_settings[17]
port 9 nsew signal input
rlabel metal3 s 0 90040 800 90160 6 custom_settings[18]
port 10 nsew signal input
rlabel metal3 s 0 94392 800 94512 6 custom_settings[19]
port 11 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 custom_settings[1]
port 12 nsew signal input
rlabel metal3 s 0 98744 800 98864 6 custom_settings[20]
port 13 nsew signal input
rlabel metal3 s 0 103096 800 103216 6 custom_settings[21]
port 14 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 custom_settings[22]
port 15 nsew signal input
rlabel metal3 s 0 111800 800 111920 6 custom_settings[23]
port 16 nsew signal input
rlabel metal3 s 0 116152 800 116272 6 custom_settings[24]
port 17 nsew signal input
rlabel metal3 s 0 120504 800 120624 6 custom_settings[25]
port 18 nsew signal input
rlabel metal3 s 0 124856 800 124976 6 custom_settings[26]
port 19 nsew signal input
rlabel metal3 s 0 129208 800 129328 6 custom_settings[27]
port 20 nsew signal input
rlabel metal3 s 0 133560 800 133680 6 custom_settings[28]
port 21 nsew signal input
rlabel metal3 s 0 137912 800 138032 6 custom_settings[29]
port 22 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 custom_settings[2]
port 23 nsew signal input
rlabel metal3 s 0 142264 800 142384 6 custom_settings[30]
port 24 nsew signal input
rlabel metal3 s 0 146616 800 146736 6 custom_settings[31]
port 25 nsew signal input
rlabel metal3 s 0 24760 800 24880 6 custom_settings[3]
port 26 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 custom_settings[4]
port 27 nsew signal input
rlabel metal3 s 0 33464 800 33584 6 custom_settings[5]
port 28 nsew signal input
rlabel metal3 s 0 37816 800 37936 6 custom_settings[6]
port 29 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 custom_settings[7]
port 30 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 custom_settings[8]
port 31 nsew signal input
rlabel metal3 s 0 50872 800 50992 6 custom_settings[9]
port 32 nsew signal input
rlabel metal2 s 3698 149200 3754 150000 6 io_in[0]
port 33 nsew signal input
rlabel metal2 s 64418 149200 64474 150000 6 io_in[10]
port 34 nsew signal input
rlabel metal2 s 70490 149200 70546 150000 6 io_in[11]
port 35 nsew signal input
rlabel metal2 s 76562 149200 76618 150000 6 io_in[12]
port 36 nsew signal input
rlabel metal2 s 82634 149200 82690 150000 6 io_in[13]
port 37 nsew signal input
rlabel metal2 s 88706 149200 88762 150000 6 io_in[14]
port 38 nsew signal input
rlabel metal2 s 94778 149200 94834 150000 6 io_in[15]
port 39 nsew signal input
rlabel metal2 s 100850 149200 100906 150000 6 io_in[16]
port 40 nsew signal input
rlabel metal2 s 106922 149200 106978 150000 6 io_in[17]
port 41 nsew signal input
rlabel metal2 s 112994 149200 113050 150000 6 io_in[18]
port 42 nsew signal input
rlabel metal2 s 119066 149200 119122 150000 6 io_in[19]
port 43 nsew signal input
rlabel metal2 s 9770 149200 9826 150000 6 io_in[1]
port 44 nsew signal input
rlabel metal2 s 125138 149200 125194 150000 6 io_in[20]
port 45 nsew signal input
rlabel metal2 s 131210 149200 131266 150000 6 io_in[21]
port 46 nsew signal input
rlabel metal2 s 137282 149200 137338 150000 6 io_in[22]
port 47 nsew signal input
rlabel metal2 s 143354 149200 143410 150000 6 io_in[23]
port 48 nsew signal input
rlabel metal2 s 149426 149200 149482 150000 6 io_in[24]
port 49 nsew signal input
rlabel metal2 s 155498 149200 155554 150000 6 io_in[25]
port 50 nsew signal input
rlabel metal2 s 161570 149200 161626 150000 6 io_in[26]
port 51 nsew signal input
rlabel metal2 s 167642 149200 167698 150000 6 io_in[27]
port 52 nsew signal input
rlabel metal2 s 173714 149200 173770 150000 6 io_in[28]
port 53 nsew signal input
rlabel metal2 s 179786 149200 179842 150000 6 io_in[29]
port 54 nsew signal input
rlabel metal2 s 15842 149200 15898 150000 6 io_in[2]
port 55 nsew signal input
rlabel metal2 s 185858 149200 185914 150000 6 io_in[30]
port 56 nsew signal input
rlabel metal2 s 191930 149200 191986 150000 6 io_in[31]
port 57 nsew signal input
rlabel metal2 s 198002 149200 198058 150000 6 io_in[32]
port 58 nsew signal input
rlabel metal2 s 204074 149200 204130 150000 6 io_in[33]
port 59 nsew signal input
rlabel metal2 s 210146 149200 210202 150000 6 io_in[34]
port 60 nsew signal input
rlabel metal2 s 216218 149200 216274 150000 6 io_in[35]
port 61 nsew signal input
rlabel metal2 s 21914 149200 21970 150000 6 io_in[3]
port 62 nsew signal input
rlabel metal2 s 27986 149200 28042 150000 6 io_in[4]
port 63 nsew signal input
rlabel metal2 s 34058 149200 34114 150000 6 io_in[5]
port 64 nsew signal input
rlabel metal2 s 40130 149200 40186 150000 6 io_in[6]
port 65 nsew signal input
rlabel metal2 s 46202 149200 46258 150000 6 io_in[7]
port 66 nsew signal input
rlabel metal2 s 52274 149200 52330 150000 6 io_in[8]
port 67 nsew signal input
rlabel metal2 s 58346 149200 58402 150000 6 io_in[9]
port 68 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 io_oeb[0]
port 69 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 io_oeb[10]
port 70 nsew signal output
rlabel metal2 s 70490 0 70546 800 6 io_oeb[11]
port 71 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 io_oeb[12]
port 72 nsew signal output
rlabel metal2 s 82634 0 82690 800 6 io_oeb[13]
port 73 nsew signal output
rlabel metal2 s 88706 0 88762 800 6 io_oeb[14]
port 74 nsew signal output
rlabel metal2 s 94778 0 94834 800 6 io_oeb[15]
port 75 nsew signal output
rlabel metal2 s 100850 0 100906 800 6 io_oeb[16]
port 76 nsew signal output
rlabel metal2 s 106922 0 106978 800 6 io_oeb[17]
port 77 nsew signal output
rlabel metal2 s 112994 0 113050 800 6 io_oeb[18]
port 78 nsew signal output
rlabel metal2 s 119066 0 119122 800 6 io_oeb[19]
port 79 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 io_oeb[1]
port 80 nsew signal output
rlabel metal2 s 125138 0 125194 800 6 io_oeb[20]
port 81 nsew signal output
rlabel metal2 s 131210 0 131266 800 6 io_oeb[21]
port 82 nsew signal output
rlabel metal2 s 137282 0 137338 800 6 io_oeb[22]
port 83 nsew signal output
rlabel metal2 s 143354 0 143410 800 6 io_oeb[23]
port 84 nsew signal output
rlabel metal2 s 149426 0 149482 800 6 io_oeb[24]
port 85 nsew signal output
rlabel metal2 s 155498 0 155554 800 6 io_oeb[25]
port 86 nsew signal output
rlabel metal2 s 161570 0 161626 800 6 io_oeb[26]
port 87 nsew signal output
rlabel metal2 s 167642 0 167698 800 6 io_oeb[27]
port 88 nsew signal output
rlabel metal2 s 173714 0 173770 800 6 io_oeb[28]
port 89 nsew signal output
rlabel metal2 s 179786 0 179842 800 6 io_oeb[29]
port 90 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 io_oeb[2]
port 91 nsew signal output
rlabel metal2 s 185858 0 185914 800 6 io_oeb[30]
port 92 nsew signal output
rlabel metal2 s 191930 0 191986 800 6 io_oeb[31]
port 93 nsew signal output
rlabel metal2 s 198002 0 198058 800 6 io_oeb[32]
port 94 nsew signal output
rlabel metal2 s 204074 0 204130 800 6 io_oeb[33]
port 95 nsew signal output
rlabel metal2 s 210146 0 210202 800 6 io_oeb[34]
port 96 nsew signal output
rlabel metal2 s 216218 0 216274 800 6 io_oeb[35]
port 97 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 io_oeb[3]
port 98 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 io_oeb[4]
port 99 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 io_oeb[5]
port 100 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 io_oeb[6]
port 101 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 io_oeb[7]
port 102 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 io_oeb[8]
port 103 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 io_oeb[9]
port 104 nsew signal output
rlabel metal3 s 219200 3544 220000 3664 6 io_out[0]
port 105 nsew signal output
rlabel metal3 s 219200 44344 220000 44464 6 io_out[10]
port 106 nsew signal output
rlabel metal3 s 219200 48424 220000 48544 6 io_out[11]
port 107 nsew signal output
rlabel metal3 s 219200 52504 220000 52624 6 io_out[12]
port 108 nsew signal output
rlabel metal3 s 219200 56584 220000 56704 6 io_out[13]
port 109 nsew signal output
rlabel metal3 s 219200 60664 220000 60784 6 io_out[14]
port 110 nsew signal output
rlabel metal3 s 219200 64744 220000 64864 6 io_out[15]
port 111 nsew signal output
rlabel metal3 s 219200 68824 220000 68944 6 io_out[16]
port 112 nsew signal output
rlabel metal3 s 219200 72904 220000 73024 6 io_out[17]
port 113 nsew signal output
rlabel metal3 s 219200 76984 220000 77104 6 io_out[18]
port 114 nsew signal output
rlabel metal3 s 219200 81064 220000 81184 6 io_out[19]
port 115 nsew signal output
rlabel metal3 s 219200 7624 220000 7744 6 io_out[1]
port 116 nsew signal output
rlabel metal3 s 219200 85144 220000 85264 6 io_out[20]
port 117 nsew signal output
rlabel metal3 s 219200 89224 220000 89344 6 io_out[21]
port 118 nsew signal output
rlabel metal3 s 219200 93304 220000 93424 6 io_out[22]
port 119 nsew signal output
rlabel metal3 s 219200 97384 220000 97504 6 io_out[23]
port 120 nsew signal output
rlabel metal3 s 219200 101464 220000 101584 6 io_out[24]
port 121 nsew signal output
rlabel metal3 s 219200 105544 220000 105664 6 io_out[25]
port 122 nsew signal output
rlabel metal3 s 219200 109624 220000 109744 6 io_out[26]
port 123 nsew signal output
rlabel metal3 s 219200 113704 220000 113824 6 io_out[27]
port 124 nsew signal output
rlabel metal3 s 219200 117784 220000 117904 6 io_out[28]
port 125 nsew signal output
rlabel metal3 s 219200 121864 220000 121984 6 io_out[29]
port 126 nsew signal output
rlabel metal3 s 219200 11704 220000 11824 6 io_out[2]
port 127 nsew signal output
rlabel metal3 s 219200 125944 220000 126064 6 io_out[30]
port 128 nsew signal output
rlabel metal3 s 219200 130024 220000 130144 6 io_out[31]
port 129 nsew signal output
rlabel metal3 s 219200 134104 220000 134224 6 io_out[32]
port 130 nsew signal output
rlabel metal3 s 219200 138184 220000 138304 6 io_out[33]
port 131 nsew signal output
rlabel metal3 s 219200 142264 220000 142384 6 io_out[34]
port 132 nsew signal output
rlabel metal3 s 219200 146344 220000 146464 6 io_out[35]
port 133 nsew signal output
rlabel metal3 s 219200 15784 220000 15904 6 io_out[3]
port 134 nsew signal output
rlabel metal3 s 219200 19864 220000 19984 6 io_out[4]
port 135 nsew signal output
rlabel metal3 s 219200 23944 220000 24064 6 io_out[5]
port 136 nsew signal output
rlabel metal3 s 219200 28024 220000 28144 6 io_out[6]
port 137 nsew signal output
rlabel metal3 s 219200 32104 220000 32224 6 io_out[7]
port 138 nsew signal output
rlabel metal3 s 219200 36184 220000 36304 6 io_out[8]
port 139 nsew signal output
rlabel metal3 s 219200 40264 220000 40384 6 io_out[9]
port 140 nsew signal output
rlabel metal3 s 0 7352 800 7472 6 rst_n
port 141 nsew signal input
rlabel metal4 s 4208 2128 4528 147472 6 vccd1
port 142 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 147472 6 vccd1
port 142 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 147472 6 vccd1
port 142 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 147472 6 vccd1
port 142 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 147472 6 vccd1
port 142 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 147472 6 vccd1
port 142 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 147472 6 vccd1
port 142 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 147472 6 vssd1
port 143 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 147472 6 vssd1
port 143 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 147472 6 vssd1
port 143 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 147472 6 vssd1
port 143 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 147472 6 vssd1
port 143 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 147472 6 vssd1
port 143 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 147472 6 vssd1
port 143 nsew ground bidirectional
rlabel metal3 s 0 3000 800 3120 6 wb_clk_i
port 144 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 220000 150000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 107885482
string GDS_FILE /run/media/tholin/8a6b8802-051e-45a8-8492-771202e4c08a/ci2406-rej-pommedeterrible-tholin/openlane/VLIW/runs/24_05_28_20_01/results/signoff/vliw.magic.gds
string GDS_START 1681446
<< end >>

