magic
tech sky130B
magscale 1 2
timestamp 1717501102
<< viali >>
rect 2881 36193 2915 36227
rect 8125 36193 8159 36227
rect 13369 36193 13403 36227
rect 18613 36193 18647 36227
rect 20729 36193 20763 36227
rect 27169 36193 27203 36227
rect 29929 36193 29963 36227
rect 32597 36193 32631 36227
rect 34897 36193 34931 36227
rect 36737 36193 36771 36227
rect 2145 36125 2179 36159
rect 3617 36125 3651 36159
rect 4169 36125 4203 36159
rect 6101 36125 6135 36159
rect 6469 36125 6503 36159
rect 7021 36125 7055 36159
rect 8769 36125 8803 36159
rect 9781 36125 9815 36159
rect 11253 36125 11287 36159
rect 12449 36125 12483 36159
rect 13921 36125 13955 36159
rect 14473 36125 14507 36159
rect 16405 36125 16439 36159
rect 16957 36125 16991 36159
rect 17601 36125 17635 36159
rect 19073 36125 19107 36159
rect 19809 36125 19843 36159
rect 20453 36125 20487 36159
rect 22293 36125 22327 36159
rect 24501 36125 24535 36159
rect 25973 36125 26007 36159
rect 28365 36125 28399 36159
rect 29101 36125 29135 36159
rect 29653 36125 29687 36159
rect 31585 36125 31619 36159
rect 32137 36125 32171 36159
rect 34161 36125 34195 36159
rect 35909 36125 35943 36159
rect 5733 36057 5767 36091
rect 10885 36057 10919 36091
rect 16037 36057 16071 36091
rect 22753 36057 22787 36091
rect 24869 36057 24903 36091
rect 26525 36057 26559 36091
rect 1501 35989 1535 36023
rect 4721 35989 4755 36023
rect 9229 35989 9263 36023
rect 11805 35989 11839 36023
rect 15025 35989 15059 36023
rect 19257 35989 19291 36023
rect 28457 35989 28491 36023
rect 31033 35989 31067 36023
rect 33609 35989 33643 36023
rect 36185 35989 36219 36023
rect 22477 35785 22511 35819
rect 4077 35717 4111 35751
rect 4997 35717 5031 35751
rect 9321 35717 9355 35751
rect 14197 35717 14231 35751
rect 19441 35717 19475 35751
rect 20821 35717 20855 35751
rect 31033 35717 31067 35751
rect 35725 35717 35759 35751
rect 2697 35649 2731 35683
rect 3709 35649 3743 35683
rect 6009 35649 6043 35683
rect 6745 35649 6779 35683
rect 8953 35649 8987 35683
rect 10149 35649 10183 35683
rect 11989 35649 12023 35683
rect 14749 35649 14783 35683
rect 15301 35649 15335 35683
rect 17233 35649 17267 35683
rect 19993 35649 20027 35683
rect 20361 35649 20395 35683
rect 22753 35649 22787 35683
rect 24777 35649 24811 35683
rect 27537 35649 27571 35683
rect 28089 35649 28123 35683
rect 28917 35649 28951 35683
rect 30481 35649 30515 35683
rect 33517 35649 33551 35683
rect 33701 35649 33735 35683
rect 35173 35649 35207 35683
rect 2421 35581 2455 35615
rect 7205 35581 7239 35615
rect 10425 35581 10459 35615
rect 12449 35581 12483 35615
rect 15577 35581 15611 35615
rect 17693 35581 17727 35615
rect 21925 35581 21959 35615
rect 23121 35581 23155 35615
rect 25053 35581 25087 35615
rect 26617 35581 26651 35615
rect 29377 35581 29411 35615
rect 32321 35581 32355 35615
rect 33977 35581 34011 35615
rect 37013 35581 37047 35615
rect 36645 35513 36679 35547
rect 26065 35445 26099 35479
rect 27261 35445 27295 35479
rect 28549 35445 28583 35479
rect 31401 35445 31435 35479
rect 36369 35445 36403 35479
rect 36553 35445 36587 35479
rect 4445 35241 4479 35275
rect 9229 35241 9263 35275
rect 12173 35241 12207 35275
rect 14841 35241 14875 35275
rect 19257 35241 19291 35275
rect 29377 35241 29411 35275
rect 3341 35173 3375 35207
rect 3985 35173 4019 35207
rect 9965 35173 9999 35207
rect 16497 35173 16531 35207
rect 33057 35173 33091 35207
rect 37013 35173 37047 35207
rect 9873 35105 9907 35139
rect 11529 35105 11563 35139
rect 14197 35105 14231 35139
rect 19073 35105 19107 35139
rect 36185 35105 36219 35139
rect 1961 35037 1995 35071
rect 5825 35037 5859 35071
rect 7297 35037 7331 35071
rect 8769 35037 8803 35071
rect 11345 35037 11379 35071
rect 13553 35037 13587 35071
rect 16221 35037 16255 35071
rect 18245 35037 18279 35071
rect 20637 35037 20671 35071
rect 21005 35037 21039 35071
rect 22569 35037 22603 35071
rect 22845 35037 22879 35071
rect 24685 35037 24719 35071
rect 26249 35037 26283 35071
rect 26525 35037 26559 35071
rect 27997 35037 28031 35071
rect 29837 35037 29871 35071
rect 31493 35037 31527 35071
rect 31677 35037 31711 35071
rect 31944 35037 31978 35071
rect 34529 35037 34563 35071
rect 34805 35037 34839 35071
rect 36737 35037 36771 35071
rect 2206 34969 2240 35003
rect 4261 34969 4295 35003
rect 5580 34969 5614 35003
rect 7052 34969 7086 35003
rect 8524 34969 8558 35003
rect 11100 34969 11134 35003
rect 13286 34969 13320 35003
rect 15976 34969 16010 35003
rect 16773 34969 16807 35003
rect 18000 34969 18034 35003
rect 20370 34969 20404 35003
rect 22302 34969 22336 35003
rect 23112 34969 23146 35003
rect 26004 34969 26038 35003
rect 26792 34969 26826 35003
rect 28264 34969 28298 35003
rect 30104 34969 30138 35003
rect 34284 34969 34318 35003
rect 35357 34969 35391 35003
rect 36093 34969 36127 35003
rect 37381 34969 37415 35003
rect 3801 34901 3835 34935
rect 5917 34901 5951 34935
rect 7389 34901 7423 34935
rect 12081 34901 12115 34935
rect 14749 34901 14783 34935
rect 16313 34901 16347 34935
rect 16865 34901 16899 34935
rect 18429 34901 18463 34935
rect 21189 34901 21223 34935
rect 24225 34901 24259 34935
rect 24869 34901 24903 34935
rect 27905 34901 27939 34935
rect 31217 34901 31251 34935
rect 33149 34901 33183 34935
rect 36921 34901 36955 34935
rect 1961 34697 1995 34731
rect 2789 34697 2823 34731
rect 8769 34697 8803 34731
rect 8953 34697 8987 34731
rect 9689 34697 9723 34731
rect 11529 34697 11563 34731
rect 12173 34697 12207 34731
rect 17785 34697 17819 34731
rect 18981 34697 19015 34731
rect 19901 34697 19935 34731
rect 24041 34697 24075 34731
rect 24777 34697 24811 34731
rect 26249 34697 26283 34731
rect 27629 34697 27663 34731
rect 28549 34697 28583 34731
rect 5641 34629 5675 34663
rect 9413 34629 9447 34663
rect 15577 34629 15611 34663
rect 20453 34629 20487 34663
rect 20821 34629 20855 34663
rect 28365 34629 28399 34663
rect 2145 34561 2179 34595
rect 3902 34561 3936 34595
rect 4169 34561 4203 34595
rect 6009 34561 6043 34595
rect 6377 34561 6411 34595
rect 7389 34561 7423 34595
rect 10149 34561 10183 34595
rect 10609 34561 10643 34595
rect 12725 34561 12759 34595
rect 14401 34561 14435 34595
rect 14657 34561 14691 34595
rect 15209 34561 15243 34595
rect 17049 34561 17083 34595
rect 21833 34561 21867 34595
rect 22569 34561 22603 34595
rect 23397 34561 23431 34595
rect 24225 34561 24259 34595
rect 25513 34561 25547 34595
rect 27077 34561 27111 34595
rect 27813 34561 27847 34595
rect 30481 34561 30515 34595
rect 31953 34561 31987 34595
rect 33250 34561 33284 34595
rect 33517 34561 33551 34595
rect 34069 34561 34103 34595
rect 36573 34561 36607 34595
rect 36829 34561 36863 34595
rect 1501 34493 1535 34527
rect 8217 34493 8251 34527
rect 11989 34493 12023 34527
rect 16865 34493 16899 34527
rect 17693 34493 17727 34527
rect 18337 34493 18371 34527
rect 18521 34493 18555 34527
rect 19257 34493 19291 34527
rect 19993 34493 20027 34527
rect 22477 34493 22511 34527
rect 23121 34493 23155 34527
rect 24869 34493 24903 34527
rect 25329 34493 25363 34527
rect 26157 34493 26191 34527
rect 26709 34493 26743 34527
rect 29009 34493 29043 34527
rect 30021 34493 30055 34527
rect 31493 34493 31527 34527
rect 34345 34493 34379 34527
rect 1869 34425 1903 34459
rect 2697 34425 2731 34459
rect 9137 34425 9171 34459
rect 11713 34425 11747 34459
rect 18797 34425 18831 34459
rect 20177 34425 20211 34459
rect 25053 34425 25087 34459
rect 26433 34425 26467 34459
rect 28733 34425 28767 34459
rect 35449 34425 35483 34459
rect 7021 34357 7055 34391
rect 8033 34357 8067 34391
rect 13277 34357 13311 34391
rect 32137 34357 32171 34391
rect 3617 34153 3651 34187
rect 5917 34153 5951 34187
rect 6285 34153 6319 34187
rect 7665 34153 7699 34187
rect 8585 34153 8619 34187
rect 10609 34153 10643 34187
rect 12081 34153 12115 34187
rect 13185 34153 13219 34187
rect 15117 34153 15151 34187
rect 21925 34153 21959 34187
rect 23029 34153 23063 34187
rect 25421 34153 25455 34187
rect 26065 34153 26099 34187
rect 27445 34153 27479 34187
rect 30113 34153 30147 34187
rect 32781 34153 32815 34187
rect 35357 34153 35391 34187
rect 7573 34085 7607 34119
rect 13093 34085 13127 34119
rect 14105 34085 14139 34119
rect 22017 34085 22051 34119
rect 27629 34085 27663 34119
rect 30021 34085 30055 34119
rect 35633 34085 35667 34119
rect 37105 34085 37139 34119
rect 2973 34017 3007 34051
rect 4261 34017 4295 34051
rect 5273 34017 5307 34051
rect 6929 34017 6963 34051
rect 8033 34017 8067 34051
rect 9965 34017 9999 34051
rect 12725 34017 12759 34051
rect 13277 34017 13311 34051
rect 15669 34017 15703 34051
rect 22385 34017 22419 34051
rect 22753 34017 22787 34051
rect 26617 34017 26651 34051
rect 28733 34017 28767 34051
rect 29653 34017 29687 34051
rect 31125 34017 31159 34051
rect 32045 34017 32079 34051
rect 34713 34017 34747 34051
rect 35909 34017 35943 34051
rect 2697 33949 2731 33983
rect 3801 33949 3835 33983
rect 7205 33949 7239 33983
rect 13921 33949 13955 33983
rect 14657 33949 14691 33983
rect 28089 33949 28123 33983
rect 29377 33949 29411 33983
rect 31585 33949 31619 33983
rect 31769 33949 31803 33983
rect 33241 33949 33275 33983
rect 36185 33949 36219 33983
rect 2329 33881 2363 33915
rect 27905 33881 27939 33915
rect 33609 33881 33643 33915
rect 36553 33881 36587 33915
rect 18337 33813 18371 33847
rect 27077 33813 27111 33847
rect 28641 33813 28675 33847
rect 35449 33813 35483 33847
rect 5365 33609 5399 33643
rect 6377 33609 6411 33643
rect 13277 33609 13311 33643
rect 14657 33609 14691 33643
rect 28917 33609 28951 33643
rect 31217 33609 31251 33643
rect 27997 33541 28031 33575
rect 28825 33541 28859 33575
rect 30481 33541 30515 33575
rect 32965 33541 32999 33575
rect 35112 33541 35146 33575
rect 2697 33473 2731 33507
rect 2881 33473 2915 33507
rect 4721 33473 4755 33507
rect 6837 33473 6871 33507
rect 13921 33473 13955 33507
rect 14565 33473 14599 33507
rect 29561 33473 29595 33507
rect 29929 33473 29963 33507
rect 31309 33473 31343 33507
rect 32413 33473 32447 33507
rect 32597 33473 32631 33507
rect 35357 33473 35391 33507
rect 35449 33473 35483 33507
rect 35705 33473 35739 33507
rect 2421 33405 2455 33439
rect 3341 33405 3375 33439
rect 6009 33405 6043 33439
rect 15117 33405 15151 33439
rect 15393 33405 15427 33439
rect 30665 33405 30699 33439
rect 31953 33405 31987 33439
rect 6561 33337 6595 33371
rect 14749 33337 14783 33371
rect 33977 33337 34011 33371
rect 5457 33269 5491 33303
rect 33609 33269 33643 33303
rect 36829 33269 36863 33303
rect 32505 33065 32539 33099
rect 33057 33065 33091 33099
rect 32873 32997 32907 33031
rect 35081 32997 35115 33031
rect 1593 32929 1627 32963
rect 29653 32929 29687 32963
rect 31217 32929 31251 32963
rect 31769 32929 31803 32963
rect 34253 32929 34287 32963
rect 2605 32861 2639 32895
rect 2973 32861 3007 32895
rect 5089 32861 5123 32895
rect 30481 32861 30515 32895
rect 31861 32861 31895 32895
rect 32597 32861 32631 32895
rect 33333 32861 33367 32895
rect 36001 32861 36035 32895
rect 36277 32861 36311 32895
rect 4537 32793 4571 32827
rect 31033 32793 31067 32827
rect 34805 32793 34839 32827
rect 37197 32793 37231 32827
rect 3525 32725 3559 32759
rect 30297 32725 30331 32759
rect 35265 32725 35299 32759
rect 35357 32725 35391 32759
rect 4997 32521 5031 32555
rect 31953 32521 31987 32555
rect 3065 32453 3099 32487
rect 32689 32453 32723 32487
rect 36185 32453 36219 32487
rect 36737 32453 36771 32487
rect 2605 32385 2639 32419
rect 4261 32385 4295 32419
rect 34161 32385 34195 32419
rect 35633 32385 35667 32419
rect 35817 32385 35851 32419
rect 1593 32317 1627 32351
rect 4445 32317 4479 32351
rect 30665 32317 30699 32351
rect 31217 32317 31251 32351
rect 31401 32317 31435 32351
rect 33701 32317 33735 32351
rect 35173 32317 35207 32351
rect 32321 32249 32355 32283
rect 32229 32181 32263 32215
rect 31493 31977 31527 32011
rect 36829 31977 36863 32011
rect 31401 31909 31435 31943
rect 36921 31909 36955 31943
rect 37013 31909 37047 31943
rect 2421 31841 2455 31875
rect 30757 31841 30791 31875
rect 32137 31841 32171 31875
rect 33241 31841 33275 31875
rect 33977 31841 34011 31875
rect 35449 31841 35483 31875
rect 37381 31841 37415 31875
rect 2697 31773 2731 31807
rect 2973 31773 3007 31807
rect 3525 31773 3559 31807
rect 3801 31773 3835 31807
rect 8125 31773 8159 31807
rect 8769 31773 8803 31807
rect 32321 31773 32355 31807
rect 32873 31773 32907 31807
rect 34529 31773 34563 31807
rect 34805 31773 34839 31807
rect 35705 31773 35739 31807
rect 33793 31705 33827 31739
rect 4445 31637 4479 31671
rect 35357 31637 35391 31671
rect 3617 31433 3651 31467
rect 34161 31433 34195 31467
rect 36829 31433 36863 31467
rect 36277 31365 36311 31399
rect 2605 31297 2639 31331
rect 4261 31297 4295 31331
rect 32781 31297 32815 31331
rect 35449 31297 35483 31331
rect 35771 31297 35805 31331
rect 1593 31229 1627 31263
rect 2881 31229 2915 31263
rect 33517 31229 33551 31263
rect 35173 31229 35207 31263
rect 33425 31161 33459 31195
rect 3525 31093 3559 31127
rect 2881 30889 2915 30923
rect 3801 30889 3835 30923
rect 33793 30889 33827 30923
rect 4629 30821 4663 30855
rect 35081 30821 35115 30855
rect 2421 30753 2455 30787
rect 4997 30753 5031 30787
rect 33241 30753 33275 30787
rect 34529 30753 34563 30787
rect 2697 30685 2731 30719
rect 3433 30685 3467 30719
rect 4445 30685 4479 30719
rect 33885 30685 33919 30719
rect 35357 30685 35391 30719
rect 36001 30685 36035 30719
rect 36277 30685 36311 30719
rect 34805 30617 34839 30651
rect 37197 30617 37231 30651
rect 4537 30549 4571 30583
rect 35265 30549 35299 30583
rect 36829 30345 36863 30379
rect 3433 30277 3467 30311
rect 34621 30277 34655 30311
rect 35694 30277 35728 30311
rect 3085 30209 3119 30243
rect 3341 30209 3375 30243
rect 33977 30209 34011 30243
rect 35265 30209 35299 30243
rect 35449 30209 35483 30243
rect 4077 30141 4111 30175
rect 1961 30005 1995 30039
rect 34713 30005 34747 30039
rect 1961 29801 1995 29835
rect 3801 29801 3835 29835
rect 6285 29801 6319 29835
rect 10885 29801 10919 29835
rect 35081 29801 35115 29835
rect 37381 29801 37415 29835
rect 6929 29665 6963 29699
rect 35357 29665 35391 29699
rect 36461 29665 36495 29699
rect 3341 29597 3375 29631
rect 4353 29597 4387 29631
rect 11529 29597 11563 29631
rect 36001 29597 36035 29631
rect 36185 29597 36219 29631
rect 3096 29529 3130 29563
rect 4353 29257 4387 29291
rect 32781 29257 32815 29291
rect 4813 29189 4847 29223
rect 5365 29189 5399 29223
rect 2697 29121 2731 29155
rect 30389 29121 30423 29155
rect 34437 29121 34471 29155
rect 35817 29121 35851 29155
rect 1593 29053 1627 29087
rect 2973 29053 3007 29087
rect 3617 29053 3651 29087
rect 4169 29053 4203 29087
rect 20453 29053 20487 29087
rect 32137 29053 32171 29087
rect 35633 29053 35667 29087
rect 36921 29053 36955 29087
rect 4537 28985 4571 29019
rect 4997 28985 5031 29019
rect 19901 28985 19935 29019
rect 28457 28985 28491 29019
rect 29101 28985 29135 29019
rect 34713 28985 34747 29019
rect 34989 28985 35023 29019
rect 3525 28917 3559 28951
rect 4905 28917 4939 28951
rect 34897 28917 34931 28951
rect 3341 28713 3375 28747
rect 19901 28713 19935 28747
rect 31033 28713 31067 28747
rect 32689 28713 32723 28747
rect 36829 28713 36863 28747
rect 35449 28577 35483 28611
rect 1961 28509 1995 28543
rect 3893 28509 3927 28543
rect 19257 28509 19291 28543
rect 31217 28509 31251 28543
rect 34805 28509 34839 28543
rect 35705 28509 35739 28543
rect 2228 28441 2262 28475
rect 4445 28373 4479 28407
rect 35357 28373 35391 28407
rect 3617 28101 3651 28135
rect 36185 28101 36219 28135
rect 2605 28033 2639 28067
rect 4169 28033 4203 28067
rect 34989 28033 35023 28067
rect 35817 28033 35851 28067
rect 1593 27965 1627 27999
rect 35633 27965 35667 27999
rect 3801 27557 3835 27591
rect 4629 27557 4663 27591
rect 35173 27557 35207 27591
rect 2421 27489 2455 27523
rect 4997 27489 5031 27523
rect 34529 27489 34563 27523
rect 34805 27489 34839 27523
rect 2697 27421 2731 27455
rect 2881 27421 2915 27455
rect 3525 27421 3559 27455
rect 4445 27421 4479 27455
rect 36001 27421 36035 27455
rect 36277 27421 36311 27455
rect 37289 27353 37323 27387
rect 4537 27285 4571 27319
rect 35265 27285 35299 27319
rect 35357 27285 35391 27319
rect 3341 27081 3375 27115
rect 4813 27081 4847 27115
rect 13461 27081 13495 27115
rect 16773 27081 16807 27115
rect 36829 27081 36863 27115
rect 3433 27013 3467 27047
rect 5549 27013 5583 27047
rect 35694 27013 35728 27047
rect 1961 26945 1995 26979
rect 2228 26945 2262 26979
rect 3985 26945 4019 26979
rect 14585 26945 14619 26979
rect 14841 26945 14875 26979
rect 17601 26945 17635 26979
rect 35265 26945 35299 26979
rect 35449 26945 35483 26979
rect 4169 26877 4203 26911
rect 4905 26877 4939 26911
rect 17233 26877 17267 26911
rect 16957 26809 16991 26843
rect 17417 26741 17451 26775
rect 17877 26741 17911 26775
rect 34713 26741 34747 26775
rect 4445 26537 4479 26571
rect 31493 26537 31527 26571
rect 4537 26469 4571 26503
rect 1961 26401 1995 26435
rect 5273 26401 5307 26435
rect 35357 26401 35391 26435
rect 36461 26401 36495 26435
rect 3801 26333 3835 26367
rect 4721 26333 4755 26367
rect 4905 26333 4939 26367
rect 30849 26333 30883 26367
rect 36001 26333 36035 26367
rect 36185 26333 36219 26367
rect 2228 26265 2262 26299
rect 7021 26265 7055 26299
rect 7389 26265 7423 26299
rect 17325 26265 17359 26299
rect 34989 26265 35023 26299
rect 3341 26197 3375 26231
rect 8309 25993 8343 26027
rect 20361 25993 20395 26027
rect 2697 25857 2731 25891
rect 9597 25857 9631 25891
rect 35909 25857 35943 25891
rect 1593 25789 1627 25823
rect 2973 25789 3007 25823
rect 3617 25789 3651 25823
rect 4169 25789 4203 25823
rect 4813 25789 4847 25823
rect 5365 25789 5399 25823
rect 19717 25789 19751 25823
rect 34437 25789 34471 25823
rect 35633 25789 35667 25823
rect 36921 25789 36955 25823
rect 4537 25721 4571 25755
rect 4997 25721 5031 25755
rect 9965 25721 9999 25755
rect 34713 25721 34747 25755
rect 34989 25721 35023 25755
rect 3525 25653 3559 25687
rect 4353 25653 4387 25687
rect 4905 25653 4939 25687
rect 34897 25653 34931 25687
rect 3341 25449 3375 25483
rect 31585 25449 31619 25483
rect 36829 25449 36863 25483
rect 1961 25245 1995 25279
rect 2228 25245 2262 25279
rect 3801 25245 3835 25279
rect 30941 25245 30975 25279
rect 34805 25245 34839 25279
rect 35449 25245 35483 25279
rect 35705 25245 35739 25279
rect 4445 25109 4479 25143
rect 35357 25109 35391 25143
rect 35633 24905 35667 24939
rect 3617 24837 3651 24871
rect 2605 24769 2639 24803
rect 4169 24769 4203 24803
rect 34989 24769 35023 24803
rect 35817 24769 35851 24803
rect 36185 24769 36219 24803
rect 1593 24701 1627 24735
rect 4813 24701 4847 24735
rect 4445 24633 4479 24667
rect 4353 24565 4387 24599
rect 35173 24293 35207 24327
rect 3341 24157 3375 24191
rect 3801 24157 3835 24191
rect 36001 24157 36035 24191
rect 36277 24157 36311 24191
rect 3096 24089 3130 24123
rect 34529 24089 34563 24123
rect 34805 24089 34839 24123
rect 37289 24089 37323 24123
rect 1961 24021 1995 24055
rect 4445 24021 4479 24055
rect 35265 24021 35299 24055
rect 35357 24021 35391 24055
rect 3341 23817 3375 23851
rect 4077 23817 4111 23851
rect 36829 23817 36863 23851
rect 2228 23749 2262 23783
rect 35694 23749 35728 23783
rect 4721 23681 4755 23715
rect 34805 23681 34839 23715
rect 1961 23613 1995 23647
rect 3433 23613 3467 23647
rect 35449 23613 35483 23647
rect 4169 23477 4203 23511
rect 35357 23477 35391 23511
rect 29009 23273 29043 23307
rect 2421 23137 2455 23171
rect 3525 23137 3559 23171
rect 36461 23137 36495 23171
rect 2697 23069 2731 23103
rect 2881 23069 2915 23103
rect 28365 23069 28399 23103
rect 35449 23069 35483 23103
rect 36001 23069 36035 23103
rect 36185 23069 36219 23103
rect 36093 22729 36127 22763
rect 2605 22593 2639 22627
rect 1593 22525 1627 22559
rect 3433 22525 3467 22559
rect 4077 22525 4111 22559
rect 36461 22525 36495 22559
rect 3801 22457 3835 22491
rect 2881 22389 2915 22423
rect 3617 22389 3651 22423
rect 37105 22389 37139 22423
rect 35633 22117 35667 22151
rect 36001 22049 36035 22083
rect 3341 21981 3375 22015
rect 4445 21981 4479 22015
rect 20729 21981 20763 22015
rect 36185 21981 36219 22015
rect 3096 21913 3130 21947
rect 20462 21913 20496 21947
rect 36553 21913 36587 21947
rect 1961 21845 1995 21879
rect 3801 21845 3835 21879
rect 19349 21845 19383 21879
rect 21097 21845 21131 21879
rect 35541 21845 35575 21879
rect 29653 21641 29687 21675
rect 29929 21641 29963 21675
rect 2329 21573 2363 21607
rect 36921 21573 36955 21607
rect 2697 21505 2731 21539
rect 2881 21505 2915 21539
rect 3525 21505 3559 21539
rect 28273 21505 28307 21539
rect 28529 21505 28563 21539
rect 35909 21505 35943 21539
rect 4077 21437 4111 21471
rect 3801 21369 3835 21403
rect 3617 21301 3651 21335
rect 36829 21097 36863 21131
rect 4629 21029 4663 21063
rect 4997 20961 5031 20995
rect 34805 20961 34839 20995
rect 35449 20961 35483 20995
rect 2697 20893 2731 20927
rect 2973 20893 3007 20927
rect 3801 20893 3835 20927
rect 4353 20893 4387 20927
rect 35705 20893 35739 20927
rect 2329 20825 2363 20859
rect 35357 20825 35391 20859
rect 3525 20757 3559 20791
rect 4537 20757 4571 20791
rect 3433 20553 3467 20587
rect 20269 20553 20303 20587
rect 2228 20417 2262 20451
rect 20729 20417 20763 20451
rect 21097 20417 21131 20451
rect 35633 20417 35667 20451
rect 35817 20417 35851 20451
rect 1961 20349 1995 20383
rect 3985 20349 4019 20383
rect 35081 20349 35115 20383
rect 36093 20349 36127 20383
rect 3341 20281 3375 20315
rect 20453 20281 20487 20315
rect 25789 20009 25823 20043
rect 35449 20009 35483 20043
rect 1593 19873 1627 19907
rect 2973 19873 3007 19907
rect 35817 19873 35851 19907
rect 37197 19873 37231 19907
rect 2605 19805 2639 19839
rect 24409 19805 24443 19839
rect 26065 19805 26099 19839
rect 35541 19805 35575 19839
rect 36185 19805 36219 19839
rect 24676 19737 24710 19771
rect 3525 19669 3559 19703
rect 1685 19465 1719 19499
rect 3341 19465 3375 19499
rect 20361 19465 20395 19499
rect 1777 19397 1811 19431
rect 2228 19329 2262 19363
rect 3893 19329 3927 19363
rect 21649 19329 21683 19363
rect 35817 19329 35851 19363
rect 1961 19261 1995 19295
rect 27537 19261 27571 19295
rect 34989 19261 35023 19295
rect 36921 19261 36955 19295
rect 3525 19193 3559 19227
rect 3433 19125 3467 19159
rect 26985 19125 27019 19159
rect 35633 19125 35667 19159
rect 1869 18921 1903 18955
rect 35449 18853 35483 18887
rect 37105 18853 37139 18887
rect 3341 18785 3375 18819
rect 35265 18785 35299 18819
rect 4353 18717 4387 18751
rect 36829 18717 36863 18751
rect 3096 18649 3130 18683
rect 36584 18649 36618 18683
rect 37381 18649 37415 18683
rect 1961 18581 1995 18615
rect 3801 18581 3835 18615
rect 34713 18581 34747 18615
rect 36921 18581 36955 18615
rect 3617 18377 3651 18411
rect 22477 18377 22511 18411
rect 24133 18377 24167 18411
rect 34989 18377 35023 18411
rect 36737 18377 36771 18411
rect 2504 18309 2538 18343
rect 34345 18309 34379 18343
rect 34437 18309 34471 18343
rect 36185 18309 36219 18343
rect 1593 18241 1627 18275
rect 2237 18241 2271 18275
rect 23949 18241 23983 18275
rect 35541 18241 35575 18275
rect 35817 18241 35851 18275
rect 3709 18173 3743 18207
rect 4169 18173 4203 18207
rect 21833 18173 21867 18207
rect 3801 18105 3835 18139
rect 34713 18105 34747 18139
rect 2145 18037 2179 18071
rect 4537 18037 4571 18071
rect 34897 18037 34931 18071
rect 27537 17833 27571 17867
rect 3525 17765 3559 17799
rect 27445 17765 27479 17799
rect 1593 17697 1627 17731
rect 3801 17697 3835 17731
rect 2605 17629 2639 17663
rect 2881 17629 2915 17663
rect 8217 17629 8251 17663
rect 33977 17629 34011 17663
rect 35265 17629 35299 17663
rect 35449 17629 35483 17663
rect 35705 17629 35739 17663
rect 27077 17561 27111 17595
rect 4445 17493 4479 17527
rect 7573 17493 7607 17527
rect 27905 17493 27939 17527
rect 34529 17493 34563 17527
rect 34713 17493 34747 17527
rect 36829 17493 36863 17527
rect 34989 17289 35023 17323
rect 2329 17221 2363 17255
rect 2697 17153 2731 17187
rect 3994 17153 4028 17187
rect 4261 17153 4295 17187
rect 35817 17153 35851 17187
rect 4905 17085 4939 17119
rect 35633 17085 35667 17119
rect 36277 17085 36311 17119
rect 2881 16949 2915 16983
rect 4353 16949 4387 16983
rect 20913 16949 20947 16983
rect 34529 16745 34563 16779
rect 20545 16677 20579 16711
rect 21373 16677 21407 16711
rect 21925 16677 21959 16711
rect 35081 16677 35115 16711
rect 3433 16609 3467 16643
rect 4721 16609 4755 16643
rect 15485 16609 15519 16643
rect 20269 16609 20303 16643
rect 20821 16609 20855 16643
rect 21097 16609 21131 16643
rect 34805 16609 34839 16643
rect 37197 16609 37231 16643
rect 1593 16541 1627 16575
rect 2605 16541 2639 16575
rect 4353 16541 4387 16575
rect 36001 16541 36035 16575
rect 36277 16541 36311 16575
rect 4966 16473 5000 16507
rect 15730 16473 15764 16507
rect 2881 16405 2915 16439
rect 3801 16405 3835 16439
rect 6101 16405 6135 16439
rect 16865 16405 16899 16439
rect 20361 16405 20395 16439
rect 21557 16405 21591 16439
rect 22293 16405 22327 16439
rect 35265 16405 35299 16439
rect 35357 16405 35391 16439
rect 4261 16201 4295 16235
rect 13277 16201 13311 16235
rect 13645 16201 13679 16235
rect 36829 16201 36863 16235
rect 2329 16133 2363 16167
rect 3801 16133 3835 16167
rect 4537 16133 4571 16167
rect 12817 16133 12851 16167
rect 35694 16133 35728 16167
rect 2697 16065 2731 16099
rect 2881 16065 2915 16099
rect 20177 16065 20211 16099
rect 20444 16065 20478 16099
rect 21833 16065 21867 16099
rect 22089 16065 22123 16099
rect 35265 16065 35299 16099
rect 35449 16065 35483 16099
rect 3525 15929 3559 15963
rect 4077 15929 4111 15963
rect 13093 15929 13127 15963
rect 21557 15861 21591 15895
rect 23213 15861 23247 15895
rect 23581 15861 23615 15895
rect 34713 15861 34747 15895
rect 3341 15657 3375 15691
rect 12633 15657 12667 15691
rect 21925 15657 21959 15691
rect 3157 15589 3191 15623
rect 11897 15589 11931 15623
rect 21833 15589 21867 15623
rect 21465 15521 21499 15555
rect 35357 15521 35391 15555
rect 2697 15453 2731 15487
rect 4445 15453 4479 15487
rect 12265 15453 12299 15487
rect 22017 15453 22051 15487
rect 36001 15453 36035 15487
rect 36185 15453 36219 15487
rect 2329 15385 2363 15419
rect 2881 15385 2915 15419
rect 36553 15385 36587 15419
rect 4077 15317 4111 15351
rect 4261 15317 4295 15351
rect 11805 15317 11839 15351
rect 22661 15317 22695 15351
rect 34989 15317 35023 15351
rect 22109 15113 22143 15147
rect 1593 15045 1627 15079
rect 36921 15045 36955 15079
rect 2605 14977 2639 15011
rect 35817 14977 35851 15011
rect 2881 14909 2915 14943
rect 3525 14909 3559 14943
rect 4077 14909 4111 14943
rect 34437 14909 34471 14943
rect 35081 14909 35115 14943
rect 3801 14841 3835 14875
rect 34713 14841 34747 14875
rect 3617 14773 3651 14807
rect 4353 14773 4387 14807
rect 34897 14773 34931 14807
rect 35633 14773 35667 14807
rect 1961 14569 1995 14603
rect 35357 14569 35391 14603
rect 3341 14433 3375 14467
rect 4353 14433 4387 14467
rect 35449 14433 35483 14467
rect 3085 14365 3119 14399
rect 34805 14365 34839 14399
rect 35705 14365 35739 14399
rect 3801 14229 3835 14263
rect 36829 14229 36863 14263
rect 34989 14025 35023 14059
rect 2697 13889 2731 13923
rect 2881 13889 2915 13923
rect 25329 13889 25363 13923
rect 35633 13889 35667 13923
rect 35817 13889 35851 13923
rect 2421 13821 2455 13855
rect 3525 13821 3559 13855
rect 4077 13821 4111 13855
rect 4353 13821 4387 13855
rect 25973 13821 26007 13855
rect 36277 13821 36311 13855
rect 3801 13753 3835 13787
rect 3617 13685 3651 13719
rect 2881 13481 2915 13515
rect 35173 13413 35207 13447
rect 1593 13345 1627 13379
rect 3433 13345 3467 13379
rect 6561 13345 6595 13379
rect 23213 13345 23247 13379
rect 37197 13345 37231 13379
rect 2605 13277 2639 13311
rect 3801 13277 3835 13311
rect 11069 13277 11103 13311
rect 25789 13277 25823 13311
rect 36001 13277 36035 13311
rect 36277 13277 36311 13311
rect 34805 13209 34839 13243
rect 4445 13141 4479 13175
rect 7205 13141 7239 13175
rect 10425 13141 10459 13175
rect 23765 13141 23799 13175
rect 25973 13141 26007 13175
rect 34529 13141 34563 13175
rect 35265 13141 35299 13175
rect 35357 13141 35391 13175
rect 3341 12937 3375 12971
rect 36829 12937 36863 12971
rect 14442 12869 14476 12903
rect 35694 12869 35728 12903
rect 1961 12801 1995 12835
rect 2228 12801 2262 12835
rect 4077 12801 4111 12835
rect 14197 12801 14231 12835
rect 35265 12801 35299 12835
rect 35449 12801 35483 12835
rect 3433 12597 3467 12631
rect 15577 12597 15611 12631
rect 34713 12597 34747 12631
rect 3433 12257 3467 12291
rect 35357 12257 35391 12291
rect 2697 12189 2731 12223
rect 2881 12189 2915 12223
rect 36001 12189 36035 12223
rect 36185 12189 36219 12223
rect 2329 12121 2363 12155
rect 36553 12121 36587 12155
rect 34989 12053 35023 12087
rect 1593 11781 1627 11815
rect 36921 11781 36955 11815
rect 2605 11713 2639 11747
rect 3525 11713 3559 11747
rect 35909 11713 35943 11747
rect 4077 11645 4111 11679
rect 34437 11645 34471 11679
rect 35081 11645 35115 11679
rect 3709 11577 3743 11611
rect 34713 11577 34747 11611
rect 2881 11509 2915 11543
rect 3617 11509 3651 11543
rect 4353 11509 4387 11543
rect 34897 11509 34931 11543
rect 35633 11509 35667 11543
rect 35357 11305 35391 11339
rect 3341 11237 3375 11271
rect 1961 11169 1995 11203
rect 4353 11169 4387 11203
rect 35449 11169 35483 11203
rect 2228 11101 2262 11135
rect 34805 11101 34839 11135
rect 35705 11101 35739 11135
rect 3801 10965 3835 10999
rect 36829 10965 36863 10999
rect 28917 10761 28951 10795
rect 34989 10761 35023 10795
rect 2697 10625 2731 10659
rect 2881 10625 2915 10659
rect 17233 10625 17267 10659
rect 27905 10625 27939 10659
rect 29469 10625 29503 10659
rect 35817 10625 35851 10659
rect 2421 10557 2455 10591
rect 3433 10557 3467 10591
rect 4077 10557 4111 10591
rect 35541 10557 35575 10591
rect 36093 10557 36127 10591
rect 3709 10489 3743 10523
rect 3617 10421 3651 10455
rect 4353 10421 4387 10455
rect 17877 10421 17911 10455
rect 27353 10421 27387 10455
rect 2881 10217 2915 10251
rect 7573 10217 7607 10251
rect 22937 10217 22971 10251
rect 35173 10149 35207 10183
rect 1593 10081 1627 10115
rect 7021 10081 7055 10115
rect 23581 10081 23615 10115
rect 35265 10081 35299 10115
rect 37197 10081 37231 10115
rect 2605 10013 2639 10047
rect 3525 10013 3559 10047
rect 3801 10013 3835 10047
rect 17049 10013 17083 10047
rect 17325 10013 17359 10047
rect 32965 10013 32999 10047
rect 36001 10013 36035 10047
rect 36185 10013 36219 10047
rect 31217 9945 31251 9979
rect 34529 9945 34563 9979
rect 34805 9945 34839 9979
rect 4445 9877 4479 9911
rect 17141 9877 17175 9911
rect 31033 9877 31067 9911
rect 35357 9877 35391 9911
rect 3341 9673 3375 9707
rect 36829 9673 36863 9707
rect 2228 9605 2262 9639
rect 35694 9605 35728 9639
rect 1961 9537 1995 9571
rect 4077 9537 4111 9571
rect 35265 9537 35299 9571
rect 35449 9537 35483 9571
rect 3433 9333 3467 9367
rect 34713 9333 34747 9367
rect 3433 8993 3467 9027
rect 35357 8993 35391 9027
rect 2697 8925 2731 8959
rect 2881 8925 2915 8959
rect 36001 8925 36035 8959
rect 36185 8925 36219 8959
rect 2329 8857 2363 8891
rect 36553 8857 36587 8891
rect 34989 8789 35023 8823
rect 1593 8517 1627 8551
rect 36921 8517 36955 8551
rect 2605 8449 2639 8483
rect 35909 8449 35943 8483
rect 3341 8381 3375 8415
rect 34437 8381 34471 8415
rect 35081 8381 35115 8415
rect 3065 8313 3099 8347
rect 3709 8313 3743 8347
rect 34713 8313 34747 8347
rect 2881 8245 2915 8279
rect 34897 8245 34931 8279
rect 35633 8245 35667 8279
rect 11897 8041 11931 8075
rect 35357 8041 35391 8075
rect 3341 7973 3375 8007
rect 1961 7905 1995 7939
rect 3801 7905 3835 7939
rect 19809 7905 19843 7939
rect 35449 7905 35483 7939
rect 2228 7837 2262 7871
rect 34529 7837 34563 7871
rect 34805 7837 34839 7871
rect 35705 7837 35739 7871
rect 10425 7769 10459 7803
rect 12541 7769 12575 7803
rect 37289 7769 37323 7803
rect 4445 7701 4479 7735
rect 19257 7701 19291 7735
rect 33885 7701 33919 7735
rect 36829 7701 36863 7735
rect 37013 7701 37047 7735
rect 9965 7497 9999 7531
rect 28457 7497 28491 7531
rect 34989 7497 35023 7531
rect 3096 7429 3130 7463
rect 9597 7429 9631 7463
rect 28641 7429 28675 7463
rect 3341 7361 3375 7395
rect 7849 7361 7883 7395
rect 35541 7361 35575 7395
rect 35817 7361 35851 7395
rect 4353 7293 4387 7327
rect 4997 7293 5031 7327
rect 5641 7293 5675 7327
rect 5917 7293 5951 7327
rect 33517 7293 33551 7327
rect 34805 7293 34839 7327
rect 36185 7293 36219 7327
rect 5273 7225 5307 7259
rect 1961 7157 1995 7191
rect 3709 7157 3743 7191
rect 4445 7157 4479 7191
rect 5181 7157 5215 7191
rect 29929 7157 29963 7191
rect 34161 7157 34195 7191
rect 34253 7157 34287 7191
rect 4721 6885 4755 6919
rect 35173 6885 35207 6919
rect 3341 6817 3375 6851
rect 3801 6817 3835 6851
rect 4445 6817 4479 6851
rect 33793 6817 33827 6851
rect 37197 6817 37231 6851
rect 3085 6749 3119 6783
rect 33057 6749 33091 6783
rect 34529 6749 34563 6783
rect 35357 6749 35391 6783
rect 36001 6749 36035 6783
rect 36185 6749 36219 6783
rect 4997 6681 5031 6715
rect 34805 6681 34839 6715
rect 1961 6613 1995 6647
rect 4537 6613 4571 6647
rect 5365 6613 5399 6647
rect 32413 6613 32447 6647
rect 33149 6613 33183 6647
rect 33885 6613 33919 6647
rect 35265 6613 35299 6647
rect 4261 6409 4295 6443
rect 33149 6409 33183 6443
rect 36829 6409 36863 6443
rect 1593 6341 1627 6375
rect 35694 6341 35728 6375
rect 2605 6273 2639 6307
rect 3433 6273 3467 6307
rect 35265 6273 35299 6307
rect 35449 6273 35483 6307
rect 3617 6205 3651 6239
rect 18521 6205 18555 6239
rect 32597 6205 32631 6239
rect 33333 6205 33367 6239
rect 34529 6205 34563 6239
rect 34713 6205 34747 6239
rect 2881 6069 2915 6103
rect 14013 6069 14047 6103
rect 19165 6069 19199 6103
rect 33885 6069 33919 6103
rect 3525 5865 3559 5899
rect 30205 5865 30239 5899
rect 13553 5797 13587 5831
rect 14473 5797 14507 5831
rect 15393 5797 15427 5831
rect 35541 5797 35575 5831
rect 2421 5729 2455 5763
rect 2881 5729 2915 5763
rect 13461 5729 13495 5763
rect 31033 5729 31067 5763
rect 34069 5729 34103 5763
rect 35449 5729 35483 5763
rect 2697 5661 2731 5695
rect 10977 5661 11011 5695
rect 12357 5661 12391 5695
rect 13093 5661 13127 5695
rect 31677 5661 31711 5695
rect 33057 5661 33091 5695
rect 34529 5661 34563 5695
rect 35357 5661 35391 5695
rect 36185 5661 36219 5695
rect 11805 5593 11839 5627
rect 13921 5593 13955 5627
rect 14105 5593 14139 5627
rect 14841 5593 14875 5627
rect 15669 5593 15703 5627
rect 15945 5593 15979 5627
rect 32413 5593 32447 5627
rect 35909 5593 35943 5627
rect 36553 5593 36587 5627
rect 10701 5525 10735 5559
rect 11621 5525 11655 5559
rect 12541 5525 12575 5559
rect 14565 5525 14599 5559
rect 15209 5525 15243 5559
rect 29101 5525 29135 5559
rect 29745 5525 29779 5559
rect 31585 5525 31619 5559
rect 32321 5525 32355 5559
rect 34713 5525 34747 5559
rect 37105 5525 37139 5559
rect 3525 5321 3559 5355
rect 11713 5321 11747 5355
rect 14933 5321 14967 5355
rect 15853 5321 15887 5355
rect 35265 5321 35299 5355
rect 16129 5253 16163 5287
rect 34713 5253 34747 5287
rect 2697 5185 2731 5219
rect 2881 5185 2915 5219
rect 12357 5185 12391 5219
rect 13921 5185 13955 5219
rect 31401 5185 31435 5219
rect 33048 5185 33082 5219
rect 34345 5185 34379 5219
rect 35817 5185 35851 5219
rect 2421 5117 2455 5151
rect 10149 5117 10183 5151
rect 11253 5117 11287 5151
rect 13093 5117 13127 5151
rect 13737 5117 13771 5151
rect 14473 5117 14507 5151
rect 15485 5117 15519 5151
rect 16957 5117 16991 5151
rect 17141 5117 17175 5151
rect 27169 5117 27203 5151
rect 28181 5117 28215 5151
rect 28917 5117 28951 5151
rect 29469 5117 29503 5151
rect 29653 5117 29687 5151
rect 30481 5117 30515 5151
rect 32229 5117 32263 5151
rect 32781 5117 32815 5151
rect 36093 5117 36127 5151
rect 10517 5049 10551 5083
rect 13185 5049 13219 5083
rect 17509 5049 17543 5083
rect 28825 5049 28859 5083
rect 32505 5049 32539 5083
rect 34161 5049 34195 5083
rect 9965 4981 9999 5015
rect 10609 4981 10643 5015
rect 10701 4981 10735 5015
rect 12449 4981 12483 5015
rect 17601 4981 17635 5015
rect 17969 4981 18003 5015
rect 26341 4981 26375 5015
rect 27813 4981 27847 5015
rect 30297 4981 30331 5015
rect 31033 4981 31067 5015
rect 31953 4981 31987 5015
rect 32689 4981 32723 5015
rect 36829 4981 36863 5015
rect 10609 4777 10643 4811
rect 13277 4777 13311 4811
rect 29193 4777 29227 4811
rect 34713 4777 34747 4811
rect 9781 4709 9815 4743
rect 10701 4709 10735 4743
rect 18797 4709 18831 4743
rect 26157 4709 26191 4743
rect 30021 4709 30055 4743
rect 1593 4641 1627 4675
rect 10057 4641 10091 4675
rect 12081 4641 12115 4675
rect 14657 4641 14691 4675
rect 15025 4641 15059 4675
rect 16681 4641 16715 4675
rect 26249 4641 26283 4675
rect 27905 4641 27939 4675
rect 29653 4641 29687 4675
rect 31125 4641 31159 4675
rect 32597 4641 32631 4675
rect 34069 4641 34103 4675
rect 37197 4641 37231 4675
rect 2605 4573 2639 4607
rect 13185 4573 13219 4607
rect 13829 4573 13863 4607
rect 16497 4573 16531 4607
rect 18245 4573 18279 4607
rect 26341 4573 26375 4607
rect 27629 4573 27663 4607
rect 28641 4573 28675 4607
rect 31585 4573 31619 4607
rect 33057 4573 33091 4607
rect 34437 4573 34471 4607
rect 35265 4573 35299 4607
rect 35449 4573 35483 4607
rect 36277 4573 36311 4607
rect 9413 4505 9447 4539
rect 11814 4505 11848 4539
rect 18429 4505 18463 4539
rect 25513 4505 25547 4539
rect 25789 4505 25823 4539
rect 35725 4505 35759 4539
rect 9873 4437 9907 4471
rect 12541 4437 12575 4471
rect 14105 4437 14139 4471
rect 15669 4437 15703 4471
rect 15853 4437 15887 4471
rect 17233 4437 17267 4471
rect 17693 4437 17727 4471
rect 18889 4437 18923 4471
rect 19441 4437 19475 4471
rect 26985 4437 27019 4471
rect 27077 4437 27111 4471
rect 28457 4437 28491 4471
rect 30113 4437 30147 4471
rect 13277 4233 13311 4267
rect 28917 4233 28951 4267
rect 25329 4165 25363 4199
rect 35357 4165 35391 4199
rect 2697 4097 2731 4131
rect 9321 4097 9355 4131
rect 10149 4097 10183 4131
rect 11805 4097 11839 4131
rect 12061 4097 12095 4131
rect 14390 4097 14424 4131
rect 14657 4097 14691 4131
rect 15301 4097 15335 4131
rect 17601 4097 17635 4131
rect 17785 4097 17819 4131
rect 26801 4097 26835 4131
rect 26985 4097 27019 4131
rect 27793 4097 27827 4131
rect 30481 4097 30515 4131
rect 31953 4097 31987 4131
rect 33149 4097 33183 4131
rect 33416 4097 33450 4131
rect 35909 4097 35943 4131
rect 36645 4097 36679 4131
rect 2421 4029 2455 4063
rect 10609 4029 10643 4063
rect 15577 4029 15611 4063
rect 16957 4029 16991 4063
rect 18061 4029 18095 4063
rect 19165 4029 19199 4063
rect 25605 4029 25639 4063
rect 27445 4029 27479 4063
rect 27537 4029 27571 4063
rect 29285 4029 29319 4063
rect 30757 4029 30791 4063
rect 32137 4029 32171 4063
rect 36093 4029 36127 4063
rect 25053 3961 25087 3995
rect 27353 3961 27387 3995
rect 34805 3961 34839 3995
rect 9873 3893 9907 3927
rect 13185 3893 13219 3927
rect 19809 3893 19843 3927
rect 24869 3893 24903 3927
rect 32781 3893 32815 3927
rect 34529 3893 34563 3927
rect 37013 3893 37047 3927
rect 12173 3689 12207 3723
rect 13645 3689 13679 3723
rect 16037 3689 16071 3723
rect 17509 3689 17543 3723
rect 26065 3689 26099 3723
rect 29009 3689 29043 3723
rect 30941 3689 30975 3723
rect 33885 3689 33919 3723
rect 37105 3689 37139 3723
rect 29377 3621 29411 3655
rect 33977 3621 34011 3655
rect 34161 3621 34195 3655
rect 36185 3621 36219 3655
rect 1593 3553 1627 3587
rect 10149 3553 10183 3587
rect 12265 3553 12299 3587
rect 15945 3553 15979 3587
rect 19257 3553 19291 3587
rect 26433 3553 26467 3587
rect 32505 3553 32539 3587
rect 34437 3553 34471 3587
rect 34713 3553 34747 3587
rect 36737 3553 36771 3587
rect 2605 3485 2639 3519
rect 7205 3485 7239 3519
rect 8677 3485 8711 3519
rect 10609 3485 10643 3519
rect 10793 3485 10827 3519
rect 15678 3485 15712 3519
rect 17417 3485 17451 3519
rect 18889 3485 18923 3519
rect 24685 3485 24719 3519
rect 24952 3485 24986 3519
rect 26893 3485 26927 3519
rect 27445 3485 27479 3519
rect 27629 3485 27663 3519
rect 29561 3485 29595 3519
rect 31033 3485 31067 3519
rect 32772 3485 32806 3519
rect 6653 3417 6687 3451
rect 8309 3417 8343 3451
rect 11060 3417 11094 3451
rect 12510 3417 12544 3451
rect 17172 3417 17206 3451
rect 18644 3417 18678 3451
rect 27874 3417 27908 3451
rect 29828 3417 29862 3451
rect 31300 3417 31334 3451
rect 34958 3417 34992 3451
rect 37013 3417 37047 3451
rect 14565 3349 14599 3383
rect 19901 3349 19935 3383
rect 32413 3349 32447 3383
rect 36093 3349 36127 3383
rect 12081 3145 12115 3179
rect 18797 3145 18831 3179
rect 25329 3145 25363 3179
rect 26801 3145 26835 3179
rect 26985 3145 27019 3179
rect 29561 3145 29595 3179
rect 31033 3145 31067 3179
rect 33149 3145 33183 3179
rect 35081 3145 35115 3179
rect 15301 3077 15335 3111
rect 17684 3077 17718 3111
rect 20637 3077 20671 3111
rect 26341 3077 26375 3111
rect 28098 3077 28132 3111
rect 30389 3077 30423 3111
rect 31861 3077 31895 3111
rect 36185 3077 36219 3111
rect 2605 3009 2639 3043
rect 8309 3009 8343 3043
rect 9781 3009 9815 3043
rect 11253 3009 11287 3043
rect 13461 3009 13495 3043
rect 14933 3009 14967 3043
rect 15761 3009 15795 3043
rect 17325 3009 17359 3043
rect 17417 3009 17451 3043
rect 19625 3009 19659 3043
rect 22017 3009 22051 3043
rect 23397 3009 23431 3043
rect 26065 3009 26099 3043
rect 28365 3009 28399 3043
rect 28549 3009 28583 3043
rect 30021 3009 30055 3043
rect 32229 3009 32263 3043
rect 32781 3009 32815 3043
rect 33609 3009 33643 3043
rect 35817 3009 35851 3043
rect 1593 2941 1627 2975
rect 7665 2941 7699 2975
rect 9229 2941 9263 2975
rect 10977 2941 11011 2975
rect 11621 2941 11655 2975
rect 12357 2941 12391 2975
rect 12909 2941 12943 2975
rect 14657 2941 14691 2975
rect 18889 2941 18923 2975
rect 19349 2941 19383 2975
rect 20085 2941 20119 2975
rect 22293 2941 22327 2975
rect 23949 2941 23983 2975
rect 25789 2941 25823 2975
rect 29101 2941 29135 2975
rect 31401 2941 31435 2975
rect 34069 2941 34103 2975
rect 35541 2941 35575 2975
rect 36737 2941 36771 2975
rect 11989 2873 12023 2907
rect 18981 2873 19015 2907
rect 26709 2873 26743 2907
rect 31585 2873 31619 2907
rect 35173 2873 35207 2907
rect 2881 2805 2915 2839
rect 16681 2805 16715 2839
rect 12449 2601 12483 2635
rect 15025 2601 15059 2635
rect 16681 2601 16715 2635
rect 19257 2601 19291 2635
rect 26157 2601 26191 2635
rect 28457 2601 28491 2635
rect 31033 2601 31067 2635
rect 33149 2601 33183 2635
rect 33609 2601 33643 2635
rect 36185 2601 36219 2635
rect 37289 2601 37323 2635
rect 9413 2533 9447 2567
rect 2421 2465 2455 2499
rect 5733 2465 5767 2499
rect 8309 2465 8343 2499
rect 10885 2465 10919 2499
rect 14473 2465 14507 2499
rect 17233 2465 17267 2499
rect 18153 2465 18187 2499
rect 19901 2465 19935 2499
rect 20453 2465 20487 2499
rect 22201 2465 22235 2499
rect 24869 2465 24903 2499
rect 27445 2465 27479 2499
rect 30021 2465 30055 2499
rect 31585 2465 31619 2499
rect 32505 2465 32539 2499
rect 35173 2465 35207 2499
rect 36737 2465 36771 2499
rect 2697 2397 2731 2431
rect 3341 2397 3375 2431
rect 4721 2397 4755 2431
rect 6193 2397 6227 2431
rect 8769 2397 8803 2431
rect 9229 2397 9263 2431
rect 11161 2397 11195 2431
rect 11897 2397 11931 2431
rect 12725 2397 12759 2431
rect 15209 2397 15243 2431
rect 17877 2397 17911 2431
rect 20085 2397 20119 2431
rect 21925 2397 21959 2431
rect 24409 2397 24443 2431
rect 26709 2397 26743 2431
rect 26985 2397 27019 2431
rect 29009 2397 29043 2431
rect 29561 2397 29595 2431
rect 32229 2397 32263 2431
rect 34161 2397 34195 2431
rect 34713 2397 34747 2431
rect 37473 2397 37507 2431
rect 13553 2329 13587 2363
rect 16313 2329 16347 2363
<< metal1 >>
rect 1104 36474 37812 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 37812 36474
rect 1104 36400 37812 36422
rect 29362 36252 29368 36304
rect 29420 36292 29426 36304
rect 29420 36264 32628 36292
rect 29420 36252 29426 36264
rect 2866 36184 2872 36236
rect 2924 36184 2930 36236
rect 8110 36184 8116 36236
rect 8168 36184 8174 36236
rect 13354 36184 13360 36236
rect 13412 36184 13418 36236
rect 18598 36184 18604 36236
rect 18656 36184 18662 36236
rect 20714 36184 20720 36236
rect 20772 36184 20778 36236
rect 25866 36184 25872 36236
rect 25924 36224 25930 36236
rect 32600 36233 32628 36264
rect 32858 36252 32864 36304
rect 32916 36292 32922 36304
rect 32916 36264 34928 36292
rect 32916 36252 32922 36264
rect 34900 36233 34928 36264
rect 27157 36227 27215 36233
rect 27157 36224 27169 36227
rect 25924 36196 27169 36224
rect 25924 36184 25930 36196
rect 27157 36193 27169 36196
rect 27203 36193 27215 36227
rect 29917 36227 29975 36233
rect 29917 36224 29929 36227
rect 27157 36187 27215 36193
rect 28368 36196 29929 36224
rect 2133 36159 2191 36165
rect 2133 36125 2145 36159
rect 2179 36156 2191 36159
rect 2774 36156 2780 36168
rect 2179 36128 2780 36156
rect 2179 36125 2191 36128
rect 2133 36119 2191 36125
rect 2774 36116 2780 36128
rect 2832 36116 2838 36168
rect 3602 36116 3608 36168
rect 3660 36116 3666 36168
rect 4157 36159 4215 36165
rect 4157 36125 4169 36159
rect 4203 36156 4215 36159
rect 4522 36156 4528 36168
rect 4203 36128 4528 36156
rect 4203 36125 4215 36128
rect 4157 36119 4215 36125
rect 4522 36116 4528 36128
rect 4580 36116 4586 36168
rect 6089 36159 6147 36165
rect 6089 36125 6101 36159
rect 6135 36156 6147 36159
rect 6457 36159 6515 36165
rect 6457 36156 6469 36159
rect 6135 36128 6469 36156
rect 6135 36125 6147 36128
rect 6089 36119 6147 36125
rect 6457 36125 6469 36128
rect 6503 36125 6515 36159
rect 6457 36119 6515 36125
rect 6546 36116 6552 36168
rect 6604 36156 6610 36168
rect 7009 36159 7067 36165
rect 7009 36156 7021 36159
rect 6604 36128 7021 36156
rect 6604 36116 6610 36128
rect 7009 36125 7021 36128
rect 7055 36125 7067 36159
rect 7009 36119 7067 36125
rect 8754 36116 8760 36168
rect 8812 36116 8818 36168
rect 9766 36116 9772 36168
rect 9824 36116 9830 36168
rect 11241 36159 11299 36165
rect 11241 36125 11253 36159
rect 11287 36156 11299 36159
rect 12158 36156 12164 36168
rect 11287 36128 12164 36156
rect 11287 36125 11299 36128
rect 11241 36119 11299 36125
rect 12158 36116 12164 36128
rect 12216 36116 12222 36168
rect 12434 36116 12440 36168
rect 12492 36116 12498 36168
rect 13909 36159 13967 36165
rect 13909 36125 13921 36159
rect 13955 36156 13967 36159
rect 14182 36156 14188 36168
rect 13955 36128 14188 36156
rect 13955 36125 13967 36128
rect 13909 36119 13967 36125
rect 14182 36116 14188 36128
rect 14240 36116 14246 36168
rect 14458 36116 14464 36168
rect 14516 36116 14522 36168
rect 16393 36159 16451 36165
rect 16393 36125 16405 36159
rect 16439 36156 16451 36159
rect 16945 36159 17003 36165
rect 16945 36156 16957 36159
rect 16439 36128 16957 36156
rect 16439 36125 16451 36128
rect 16393 36119 16451 36125
rect 16945 36125 16957 36128
rect 16991 36125 17003 36159
rect 16945 36119 17003 36125
rect 17586 36116 17592 36168
rect 17644 36116 17650 36168
rect 19061 36159 19119 36165
rect 19061 36125 19073 36159
rect 19107 36125 19119 36159
rect 19061 36119 19119 36125
rect 5721 36091 5779 36097
rect 5721 36057 5733 36091
rect 5767 36088 5779 36091
rect 6730 36088 6736 36100
rect 5767 36060 6736 36088
rect 5767 36057 5779 36060
rect 5721 36051 5779 36057
rect 6730 36048 6736 36060
rect 6788 36048 6794 36100
rect 10873 36091 10931 36097
rect 10873 36057 10885 36091
rect 10919 36088 10931 36091
rect 11974 36088 11980 36100
rect 10919 36060 11980 36088
rect 10919 36057 10931 36060
rect 10873 36051 10931 36057
rect 11974 36048 11980 36060
rect 12032 36048 12038 36100
rect 16025 36091 16083 36097
rect 16025 36057 16037 36091
rect 16071 36088 16083 36091
rect 17218 36088 17224 36100
rect 16071 36060 17224 36088
rect 16071 36057 16083 36060
rect 16025 36051 16083 36057
rect 17218 36048 17224 36060
rect 17276 36048 17282 36100
rect 19076 36088 19104 36119
rect 19334 36116 19340 36168
rect 19392 36156 19398 36168
rect 19797 36159 19855 36165
rect 19797 36156 19809 36159
rect 19392 36128 19809 36156
rect 19392 36116 19398 36128
rect 19797 36125 19809 36128
rect 19843 36125 19855 36159
rect 19797 36119 19855 36125
rect 20441 36159 20499 36165
rect 20441 36125 20453 36159
rect 20487 36156 20499 36159
rect 20806 36156 20812 36168
rect 20487 36128 20812 36156
rect 20487 36125 20499 36128
rect 20441 36119 20499 36125
rect 20806 36116 20812 36128
rect 20864 36116 20870 36168
rect 22278 36116 22284 36168
rect 22336 36116 22342 36168
rect 24026 36116 24032 36168
rect 24084 36156 24090 36168
rect 24489 36159 24547 36165
rect 24489 36156 24501 36159
rect 24084 36128 24501 36156
rect 24084 36116 24090 36128
rect 24489 36125 24501 36128
rect 24535 36125 24547 36159
rect 24489 36119 24547 36125
rect 25958 36116 25964 36168
rect 26016 36116 26022 36168
rect 28368 36165 28396 36196
rect 29917 36193 29929 36196
rect 29963 36193 29975 36227
rect 29917 36187 29975 36193
rect 32585 36227 32643 36233
rect 32585 36193 32597 36227
rect 32631 36193 32643 36227
rect 32585 36187 32643 36193
rect 34885 36227 34943 36233
rect 34885 36193 34897 36227
rect 34931 36193 34943 36227
rect 34885 36187 34943 36193
rect 35342 36184 35348 36236
rect 35400 36224 35406 36236
rect 36725 36227 36783 36233
rect 36725 36224 36737 36227
rect 35400 36196 36737 36224
rect 35400 36184 35406 36196
rect 36725 36193 36737 36196
rect 36771 36193 36783 36227
rect 36725 36187 36783 36193
rect 28353 36159 28411 36165
rect 28353 36125 28365 36159
rect 28399 36125 28411 36159
rect 28353 36119 28411 36125
rect 29086 36116 29092 36168
rect 29144 36116 29150 36168
rect 29641 36159 29699 36165
rect 29641 36125 29653 36159
rect 29687 36125 29699 36159
rect 29641 36119 29699 36125
rect 19076 36060 19472 36088
rect 19444 36032 19472 36060
rect 22738 36048 22744 36100
rect 22796 36048 22802 36100
rect 24854 36048 24860 36100
rect 24912 36048 24918 36100
rect 26513 36091 26571 36097
rect 26513 36057 26525 36091
rect 26559 36088 26571 36091
rect 29656 36088 29684 36119
rect 31570 36116 31576 36168
rect 31628 36116 31634 36168
rect 31662 36116 31668 36168
rect 31720 36156 31726 36168
rect 32125 36159 32183 36165
rect 32125 36156 32137 36159
rect 31720 36128 32137 36156
rect 31720 36116 31726 36128
rect 32125 36125 32137 36128
rect 32171 36125 32183 36159
rect 32125 36119 32183 36125
rect 34146 36116 34152 36168
rect 34204 36116 34210 36168
rect 35894 36116 35900 36168
rect 35952 36116 35958 36168
rect 26559 36060 29684 36088
rect 26559 36057 26571 36060
rect 26513 36051 26571 36057
rect 33686 36048 33692 36100
rect 33744 36088 33750 36100
rect 35526 36088 35532 36100
rect 33744 36060 35532 36088
rect 33744 36048 33750 36060
rect 35526 36048 35532 36060
rect 35584 36048 35590 36100
rect 1489 36023 1547 36029
rect 1489 35989 1501 36023
rect 1535 36020 1547 36023
rect 2130 36020 2136 36032
rect 1535 35992 2136 36020
rect 1535 35989 1547 35992
rect 1489 35983 1547 35989
rect 2130 35980 2136 35992
rect 2188 35980 2194 36032
rect 4706 35980 4712 36032
rect 4764 35980 4770 36032
rect 9214 35980 9220 36032
rect 9272 35980 9278 36032
rect 11790 35980 11796 36032
rect 11848 35980 11854 36032
rect 15010 35980 15016 36032
rect 15068 35980 15074 36032
rect 19242 35980 19248 36032
rect 19300 35980 19306 36032
rect 19426 35980 19432 36032
rect 19484 35980 19490 36032
rect 27062 35980 27068 36032
rect 27120 36020 27126 36032
rect 28445 36023 28503 36029
rect 28445 36020 28457 36023
rect 27120 35992 28457 36020
rect 27120 35980 27126 35992
rect 28445 35989 28457 35992
rect 28491 35989 28503 36023
rect 28445 35983 28503 35989
rect 29546 35980 29552 36032
rect 29604 36020 29610 36032
rect 31021 36023 31079 36029
rect 31021 36020 31033 36023
rect 29604 35992 31033 36020
rect 29604 35980 29610 35992
rect 31021 35989 31033 35992
rect 31067 35989 31079 36023
rect 31021 35983 31079 35989
rect 33594 35980 33600 36032
rect 33652 35980 33658 36032
rect 36170 35980 36176 36032
rect 36228 35980 36234 36032
rect 1104 35930 37812 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 37812 35930
rect 1104 35856 37812 35878
rect 22278 35776 22284 35828
rect 22336 35816 22342 35828
rect 22465 35819 22523 35825
rect 22465 35816 22477 35819
rect 22336 35788 22477 35816
rect 22336 35776 22342 35788
rect 22465 35785 22477 35788
rect 22511 35785 22523 35819
rect 22465 35779 22523 35785
rect 3602 35708 3608 35760
rect 3660 35748 3666 35760
rect 4065 35751 4123 35757
rect 4065 35748 4077 35751
rect 3660 35720 4077 35748
rect 3660 35708 3666 35720
rect 4065 35717 4077 35720
rect 4111 35717 4123 35751
rect 4065 35711 4123 35717
rect 4614 35708 4620 35760
rect 4672 35748 4678 35760
rect 4985 35751 5043 35757
rect 4985 35748 4997 35751
rect 4672 35720 4997 35748
rect 4672 35708 4678 35720
rect 4985 35717 4997 35720
rect 5031 35717 5043 35751
rect 4985 35711 5043 35717
rect 8754 35708 8760 35760
rect 8812 35748 8818 35760
rect 9309 35751 9367 35757
rect 9309 35748 9321 35751
rect 8812 35720 9321 35748
rect 8812 35708 8818 35720
rect 9309 35717 9321 35720
rect 9355 35717 9367 35751
rect 9309 35711 9367 35717
rect 14182 35708 14188 35760
rect 14240 35708 14246 35760
rect 19426 35708 19432 35760
rect 19484 35708 19490 35760
rect 20806 35708 20812 35760
rect 20864 35708 20870 35760
rect 31021 35751 31079 35757
rect 31021 35717 31033 35751
rect 31067 35748 31079 35751
rect 31662 35748 31668 35760
rect 31067 35720 31668 35748
rect 31067 35717 31079 35720
rect 31021 35711 31079 35717
rect 31662 35708 31668 35720
rect 31720 35708 31726 35760
rect 35713 35751 35771 35757
rect 35713 35717 35725 35751
rect 35759 35748 35771 35751
rect 35894 35748 35900 35760
rect 35759 35720 35900 35748
rect 35759 35717 35771 35720
rect 35713 35711 35771 35717
rect 35894 35708 35900 35720
rect 35952 35708 35958 35760
rect 2685 35683 2743 35689
rect 2685 35649 2697 35683
rect 2731 35680 2743 35683
rect 3142 35680 3148 35692
rect 2731 35652 3148 35680
rect 2731 35649 2743 35652
rect 2685 35643 2743 35649
rect 3142 35640 3148 35652
rect 3200 35640 3206 35692
rect 3694 35640 3700 35692
rect 3752 35640 3758 35692
rect 5718 35640 5724 35692
rect 5776 35680 5782 35692
rect 5997 35683 6055 35689
rect 5997 35680 6009 35683
rect 5776 35652 6009 35680
rect 5776 35640 5782 35652
rect 5997 35649 6009 35652
rect 6043 35649 6055 35683
rect 5997 35643 6055 35649
rect 6730 35640 6736 35692
rect 6788 35640 6794 35692
rect 8846 35640 8852 35692
rect 8904 35680 8910 35692
rect 8941 35683 8999 35689
rect 8941 35680 8953 35683
rect 8904 35652 8953 35680
rect 8904 35640 8910 35652
rect 8941 35649 8953 35652
rect 8987 35649 8999 35683
rect 8941 35643 8999 35649
rect 10134 35640 10140 35692
rect 10192 35640 10198 35692
rect 11974 35640 11980 35692
rect 12032 35640 12038 35692
rect 14642 35640 14648 35692
rect 14700 35680 14706 35692
rect 14737 35683 14795 35689
rect 14737 35680 14749 35683
rect 14700 35652 14749 35680
rect 14700 35640 14706 35652
rect 14737 35649 14749 35652
rect 14783 35649 14795 35683
rect 14737 35643 14795 35649
rect 15286 35640 15292 35692
rect 15344 35640 15350 35692
rect 17218 35640 17224 35692
rect 17276 35640 17282 35692
rect 19978 35640 19984 35692
rect 20036 35640 20042 35692
rect 20346 35640 20352 35692
rect 20404 35640 20410 35692
rect 22738 35640 22744 35692
rect 22796 35640 22802 35692
rect 24765 35683 24823 35689
rect 24765 35649 24777 35683
rect 24811 35680 24823 35683
rect 24854 35680 24860 35692
rect 24811 35652 24860 35680
rect 24811 35649 24823 35652
rect 24765 35643 24823 35649
rect 24854 35640 24860 35652
rect 24912 35640 24918 35692
rect 27522 35640 27528 35692
rect 27580 35640 27586 35692
rect 28077 35683 28135 35689
rect 28077 35649 28089 35683
rect 28123 35680 28135 35683
rect 28905 35683 28963 35689
rect 28905 35680 28917 35683
rect 28123 35652 28917 35680
rect 28123 35649 28135 35652
rect 28077 35643 28135 35649
rect 28905 35649 28917 35652
rect 28951 35649 28963 35683
rect 28905 35643 28963 35649
rect 30466 35640 30472 35692
rect 30524 35640 30530 35692
rect 33505 35683 33563 35689
rect 33505 35649 33517 35683
rect 33551 35649 33563 35683
rect 33505 35643 33563 35649
rect 2409 35615 2467 35621
rect 2409 35581 2421 35615
rect 2455 35612 2467 35615
rect 3786 35612 3792 35624
rect 2455 35584 3792 35612
rect 2455 35581 2467 35584
rect 2409 35575 2467 35581
rect 3786 35572 3792 35584
rect 3844 35572 3850 35624
rect 6362 35572 6368 35624
rect 6420 35612 6426 35624
rect 7193 35615 7251 35621
rect 7193 35612 7205 35615
rect 6420 35584 7205 35612
rect 6420 35572 6426 35584
rect 7193 35581 7205 35584
rect 7239 35581 7251 35615
rect 7193 35575 7251 35581
rect 9858 35572 9864 35624
rect 9916 35612 9922 35624
rect 10413 35615 10471 35621
rect 10413 35612 10425 35615
rect 9916 35584 10425 35612
rect 9916 35572 9922 35584
rect 10413 35581 10425 35584
rect 10459 35581 10471 35615
rect 10413 35575 10471 35581
rect 11606 35572 11612 35624
rect 11664 35612 11670 35624
rect 12437 35615 12495 35621
rect 12437 35612 12449 35615
rect 11664 35584 12449 35612
rect 11664 35572 11670 35584
rect 12437 35581 12449 35584
rect 12483 35581 12495 35615
rect 12437 35575 12495 35581
rect 15010 35572 15016 35624
rect 15068 35612 15074 35624
rect 15565 35615 15623 35621
rect 15565 35612 15577 35615
rect 15068 35584 15577 35612
rect 15068 35572 15074 35584
rect 15565 35581 15577 35584
rect 15611 35581 15623 35615
rect 15565 35575 15623 35581
rect 16850 35572 16856 35624
rect 16908 35612 16914 35624
rect 17681 35615 17739 35621
rect 17681 35612 17693 35615
rect 16908 35584 17693 35612
rect 16908 35572 16914 35584
rect 17681 35581 17693 35584
rect 17727 35581 17739 35615
rect 17681 35575 17739 35581
rect 21910 35572 21916 35624
rect 21968 35572 21974 35624
rect 22094 35572 22100 35624
rect 22152 35612 22158 35624
rect 23109 35615 23167 35621
rect 23109 35612 23121 35615
rect 22152 35584 23121 35612
rect 22152 35572 22158 35584
rect 23109 35581 23121 35584
rect 23155 35581 23167 35615
rect 23109 35575 23167 35581
rect 23842 35572 23848 35624
rect 23900 35612 23906 35624
rect 25041 35615 25099 35621
rect 25041 35612 25053 35615
rect 23900 35584 25053 35612
rect 23900 35572 23906 35584
rect 25041 35581 25053 35584
rect 25087 35581 25099 35615
rect 26605 35615 26663 35621
rect 26605 35612 26617 35615
rect 25041 35575 25099 35581
rect 26206 35584 26617 35612
rect 24762 35504 24768 35556
rect 24820 35544 24826 35556
rect 26206 35544 26234 35584
rect 26605 35581 26617 35584
rect 26651 35581 26663 35615
rect 26605 35575 26663 35581
rect 27338 35572 27344 35624
rect 27396 35612 27402 35624
rect 29365 35615 29423 35621
rect 29365 35612 29377 35615
rect 27396 35584 29377 35612
rect 27396 35572 27402 35584
rect 29365 35581 29377 35584
rect 29411 35581 29423 35615
rect 29365 35575 29423 35581
rect 30834 35572 30840 35624
rect 30892 35612 30898 35624
rect 32309 35615 32367 35621
rect 32309 35612 32321 35615
rect 30892 35584 32321 35612
rect 30892 35572 30898 35584
rect 32309 35581 32321 35584
rect 32355 35581 32367 35615
rect 33520 35612 33548 35643
rect 33686 35640 33692 35692
rect 33744 35640 33750 35692
rect 35161 35683 35219 35689
rect 35161 35649 35173 35683
rect 35207 35649 35219 35683
rect 35161 35643 35219 35649
rect 33965 35615 34023 35621
rect 33965 35612 33977 35615
rect 33520 35584 33977 35612
rect 32309 35575 32367 35581
rect 33965 35581 33977 35584
rect 34011 35581 34023 35615
rect 33965 35575 34023 35581
rect 24820 35516 26234 35544
rect 24820 35504 24826 35516
rect 32490 35504 32496 35556
rect 32548 35544 32554 35556
rect 35176 35544 35204 35643
rect 37001 35615 37059 35621
rect 37001 35612 37013 35615
rect 32548 35516 35204 35544
rect 36372 35584 37013 35612
rect 32548 35504 32554 35516
rect 36372 35488 36400 35584
rect 37001 35581 37013 35584
rect 37047 35581 37059 35615
rect 37001 35575 37059 35581
rect 36630 35504 36636 35556
rect 36688 35504 36694 35556
rect 23382 35436 23388 35488
rect 23440 35476 23446 35488
rect 26053 35479 26111 35485
rect 26053 35476 26065 35479
rect 23440 35448 26065 35476
rect 23440 35436 23446 35448
rect 26053 35445 26065 35448
rect 26099 35445 26111 35479
rect 26053 35439 26111 35445
rect 27249 35479 27307 35485
rect 27249 35445 27261 35479
rect 27295 35476 27307 35479
rect 28537 35479 28595 35485
rect 28537 35476 28549 35479
rect 27295 35448 28549 35476
rect 27295 35445 27307 35448
rect 27249 35439 27307 35445
rect 28537 35445 28549 35448
rect 28583 35476 28595 35479
rect 29914 35476 29920 35488
rect 28583 35448 29920 35476
rect 28583 35445 28595 35448
rect 28537 35439 28595 35445
rect 29914 35436 29920 35448
rect 29972 35476 29978 35488
rect 31389 35479 31447 35485
rect 31389 35476 31401 35479
rect 29972 35448 31401 35476
rect 29972 35436 29978 35448
rect 31389 35445 31401 35448
rect 31435 35445 31447 35479
rect 31389 35439 31447 35445
rect 36354 35436 36360 35488
rect 36412 35436 36418 35488
rect 36538 35436 36544 35488
rect 36596 35436 36602 35488
rect 1104 35386 37812 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 37812 35386
rect 1104 35312 37812 35334
rect 4433 35275 4491 35281
rect 4433 35241 4445 35275
rect 4479 35272 4491 35275
rect 4614 35272 4620 35284
rect 4479 35244 4620 35272
rect 4479 35241 4491 35244
rect 4433 35235 4491 35241
rect 4614 35232 4620 35244
rect 4672 35232 4678 35284
rect 9217 35275 9275 35281
rect 9217 35241 9229 35275
rect 9263 35272 9275 35275
rect 9766 35272 9772 35284
rect 9263 35244 9772 35272
rect 9263 35241 9275 35244
rect 9217 35235 9275 35241
rect 9766 35232 9772 35244
rect 9824 35232 9830 35284
rect 12161 35275 12219 35281
rect 12161 35241 12173 35275
rect 12207 35272 12219 35275
rect 12434 35272 12440 35284
rect 12207 35244 12440 35272
rect 12207 35241 12219 35244
rect 12161 35235 12219 35241
rect 12434 35232 12440 35244
rect 12492 35232 12498 35284
rect 14458 35232 14464 35284
rect 14516 35272 14522 35284
rect 14829 35275 14887 35281
rect 14829 35272 14841 35275
rect 14516 35244 14841 35272
rect 14516 35232 14522 35244
rect 14829 35241 14841 35244
rect 14875 35241 14887 35275
rect 17586 35272 17592 35284
rect 14829 35235 14887 35241
rect 16500 35244 17592 35272
rect 3329 35207 3387 35213
rect 3329 35173 3341 35207
rect 3375 35173 3387 35207
rect 3329 35167 3387 35173
rect 3973 35207 4031 35213
rect 3973 35173 3985 35207
rect 4019 35204 4031 35207
rect 4798 35204 4804 35216
rect 4019 35176 4804 35204
rect 4019 35173 4031 35176
rect 3973 35167 4031 35173
rect 3344 35136 3372 35167
rect 4798 35164 4804 35176
rect 4856 35164 4862 35216
rect 16500 35213 16528 35244
rect 17586 35232 17592 35244
rect 17644 35232 17650 35284
rect 19245 35275 19303 35281
rect 19245 35241 19257 35275
rect 19291 35272 19303 35275
rect 19334 35272 19340 35284
rect 19291 35244 19340 35272
rect 19291 35241 19303 35244
rect 19245 35235 19303 35241
rect 19334 35232 19340 35244
rect 19392 35232 19398 35284
rect 29365 35275 29423 35281
rect 29365 35241 29377 35275
rect 29411 35272 29423 35275
rect 31570 35272 31576 35284
rect 29411 35244 31576 35272
rect 29411 35241 29423 35244
rect 29365 35235 29423 35241
rect 31570 35232 31576 35244
rect 31628 35232 31634 35284
rect 33318 35272 33324 35284
rect 31680 35244 33324 35272
rect 9953 35207 10011 35213
rect 9953 35204 9965 35207
rect 9876 35176 9965 35204
rect 4614 35136 4620 35148
rect 3344 35108 4620 35136
rect 4614 35096 4620 35108
rect 4672 35096 4678 35148
rect 9876 35145 9904 35176
rect 9953 35173 9965 35176
rect 9999 35173 10011 35207
rect 9953 35167 10011 35173
rect 16485 35207 16543 35213
rect 16485 35173 16497 35207
rect 16531 35173 16543 35207
rect 16485 35167 16543 35173
rect 9861 35139 9919 35145
rect 9861 35105 9873 35139
rect 9907 35105 9919 35139
rect 9861 35099 9919 35105
rect 11517 35139 11575 35145
rect 11517 35105 11529 35139
rect 11563 35136 11575 35139
rect 11790 35136 11796 35148
rect 11563 35108 11796 35136
rect 11563 35105 11575 35108
rect 11517 35099 11575 35105
rect 11790 35096 11796 35108
rect 11848 35096 11854 35148
rect 14182 35096 14188 35148
rect 14240 35096 14246 35148
rect 19061 35139 19119 35145
rect 19061 35105 19073 35139
rect 19107 35136 19119 35139
rect 19242 35136 19248 35148
rect 19107 35108 19248 35136
rect 19107 35105 19119 35108
rect 19061 35099 19119 35105
rect 19242 35096 19248 35108
rect 19300 35096 19306 35148
rect 1946 35028 1952 35080
rect 2004 35028 2010 35080
rect 5813 35071 5871 35077
rect 5813 35037 5825 35071
rect 5859 35068 5871 35071
rect 7285 35071 7343 35077
rect 7285 35068 7297 35071
rect 5859 35040 7297 35068
rect 5859 35037 5871 35040
rect 5813 35031 5871 35037
rect 7285 35037 7297 35040
rect 7331 35068 7343 35071
rect 8757 35071 8815 35077
rect 8757 35068 8769 35071
rect 7331 35040 8769 35068
rect 7331 35037 7343 35040
rect 7285 35031 7343 35037
rect 8757 35037 8769 35040
rect 8803 35068 8815 35071
rect 9582 35068 9588 35080
rect 8803 35040 9588 35068
rect 8803 35037 8815 35040
rect 8757 35031 8815 35037
rect 9582 35028 9588 35040
rect 9640 35028 9646 35080
rect 11333 35071 11391 35077
rect 11333 35037 11345 35071
rect 11379 35037 11391 35071
rect 11333 35031 11391 35037
rect 13541 35071 13599 35077
rect 13541 35037 13553 35071
rect 13587 35037 13599 35071
rect 16209 35071 16267 35077
rect 16209 35068 16221 35071
rect 13541 35031 13599 35037
rect 14200 35040 16221 35068
rect 2038 34960 2044 35012
rect 2096 35000 2102 35012
rect 2194 35003 2252 35009
rect 2194 35000 2206 35003
rect 2096 34972 2206 35000
rect 2096 34960 2102 34972
rect 2194 34969 2206 34972
rect 2240 34969 2252 35003
rect 2194 34963 2252 34969
rect 2958 34960 2964 35012
rect 3016 35000 3022 35012
rect 4249 35003 4307 35009
rect 4249 35000 4261 35003
rect 3016 34972 4261 35000
rect 3016 34960 3022 34972
rect 4249 34969 4261 34972
rect 4295 35000 4307 35003
rect 4890 35000 4896 35012
rect 4295 34972 4896 35000
rect 4295 34969 4307 34972
rect 4249 34963 4307 34969
rect 4890 34960 4896 34972
rect 4948 34960 4954 35012
rect 5568 35003 5626 35009
rect 5568 34969 5580 35003
rect 5614 35000 5626 35003
rect 6362 35000 6368 35012
rect 5614 34972 6368 35000
rect 5614 34969 5626 34972
rect 5568 34963 5626 34969
rect 6362 34960 6368 34972
rect 6420 34960 6426 35012
rect 7040 35003 7098 35009
rect 7040 34969 7052 35003
rect 7086 35000 7098 35003
rect 7650 35000 7656 35012
rect 7086 34972 7656 35000
rect 7086 34969 7098 34972
rect 7040 34963 7098 34969
rect 7650 34960 7656 34972
rect 7708 34960 7714 35012
rect 8512 35003 8570 35009
rect 8512 34969 8524 35003
rect 8558 35000 8570 35003
rect 8938 35000 8944 35012
rect 8558 34972 8944 35000
rect 8558 34969 8570 34972
rect 8512 34963 8570 34969
rect 8938 34960 8944 34972
rect 8996 34960 9002 35012
rect 11088 35003 11146 35009
rect 11088 34969 11100 35003
rect 11134 35000 11146 35003
rect 11238 35000 11244 35012
rect 11134 34972 11244 35000
rect 11134 34969 11146 34972
rect 11088 34963 11146 34969
rect 11238 34960 11244 34972
rect 11296 34960 11302 35012
rect 11348 34944 11376 35031
rect 13170 34960 13176 35012
rect 13228 35000 13234 35012
rect 13274 35003 13332 35009
rect 13274 35000 13286 35003
rect 13228 34972 13286 35000
rect 13228 34960 13234 34972
rect 13274 34969 13286 34972
rect 13320 34969 13332 35003
rect 13274 34963 13332 34969
rect 13556 35000 13584 35031
rect 14200 35000 14228 35040
rect 16209 35037 16221 35040
rect 16255 35068 16267 35071
rect 18233 35071 18291 35077
rect 18233 35068 18245 35071
rect 16255 35040 18245 35068
rect 16255 35037 16267 35040
rect 16209 35031 16267 35037
rect 18233 35037 18245 35040
rect 18279 35037 18291 35071
rect 18233 35031 18291 35037
rect 20625 35071 20683 35077
rect 20625 35037 20637 35071
rect 20671 35068 20683 35071
rect 20993 35071 21051 35077
rect 20993 35068 21005 35071
rect 20671 35040 21005 35068
rect 20671 35037 20683 35040
rect 20625 35031 20683 35037
rect 20993 35037 21005 35040
rect 21039 35068 21051 35071
rect 22557 35071 22615 35077
rect 22557 35068 22569 35071
rect 21039 35040 22569 35068
rect 21039 35037 21051 35040
rect 20993 35031 21051 35037
rect 22557 35037 22569 35040
rect 22603 35068 22615 35071
rect 22833 35071 22891 35077
rect 22833 35068 22845 35071
rect 22603 35040 22845 35068
rect 22603 35037 22615 35040
rect 22557 35031 22615 35037
rect 22833 35037 22845 35040
rect 22879 35068 22891 35071
rect 22922 35068 22928 35080
rect 22879 35040 22928 35068
rect 22879 35037 22891 35040
rect 22833 35031 22891 35037
rect 22922 35028 22928 35040
rect 22980 35068 22986 35080
rect 24673 35071 24731 35077
rect 24673 35068 24685 35071
rect 22980 35040 24685 35068
rect 22980 35028 22986 35040
rect 24673 35037 24685 35040
rect 24719 35068 24731 35071
rect 26237 35071 26295 35077
rect 26237 35068 26249 35071
rect 24719 35040 26249 35068
rect 24719 35037 24731 35040
rect 24673 35031 24731 35037
rect 26237 35037 26249 35040
rect 26283 35068 26295 35071
rect 26513 35071 26571 35077
rect 26513 35068 26525 35071
rect 26283 35040 26525 35068
rect 26283 35037 26295 35040
rect 26237 35031 26295 35037
rect 26513 35037 26525 35040
rect 26559 35068 26571 35071
rect 27985 35071 28043 35077
rect 27985 35068 27997 35071
rect 26559 35040 27997 35068
rect 26559 35037 26571 35040
rect 26513 35031 26571 35037
rect 27985 35037 27997 35040
rect 28031 35068 28043 35071
rect 29825 35071 29883 35077
rect 29825 35068 29837 35071
rect 28031 35040 29837 35068
rect 28031 35037 28043 35040
rect 27985 35031 28043 35037
rect 29825 35037 29837 35040
rect 29871 35068 29883 35071
rect 29914 35068 29920 35080
rect 29871 35040 29920 35068
rect 29871 35037 29883 35040
rect 29825 35031 29883 35037
rect 29914 35028 29920 35040
rect 29972 35068 29978 35080
rect 31680 35077 31708 35244
rect 33318 35232 33324 35244
rect 33376 35232 33382 35284
rect 36538 35272 36544 35284
rect 33520 35244 36544 35272
rect 33045 35207 33103 35213
rect 33045 35173 33057 35207
rect 33091 35204 33103 35207
rect 33410 35204 33416 35216
rect 33091 35176 33416 35204
rect 33091 35173 33103 35176
rect 33045 35167 33103 35173
rect 33410 35164 33416 35176
rect 33468 35164 33474 35216
rect 31481 35071 31539 35077
rect 31481 35068 31493 35071
rect 29972 35040 31493 35068
rect 29972 35028 29978 35040
rect 31481 35037 31493 35040
rect 31527 35037 31539 35071
rect 31481 35031 31539 35037
rect 31665 35071 31723 35077
rect 31665 35037 31677 35071
rect 31711 35037 31723 35071
rect 31665 35031 31723 35037
rect 31932 35071 31990 35077
rect 31932 35037 31944 35071
rect 31978 35068 31990 35071
rect 33520 35068 33548 35244
rect 36538 35232 36544 35244
rect 36596 35232 36602 35284
rect 34514 35164 34520 35216
rect 34572 35164 34578 35216
rect 36446 35164 36452 35216
rect 36504 35204 36510 35216
rect 37001 35207 37059 35213
rect 37001 35204 37013 35207
rect 36504 35176 37013 35204
rect 36504 35164 36510 35176
rect 37001 35173 37013 35176
rect 37047 35173 37059 35207
rect 37001 35167 37059 35173
rect 34532 35136 34560 35164
rect 36173 35139 36231 35145
rect 36173 35136 36185 35139
rect 34440 35108 34560 35136
rect 35866 35108 36185 35136
rect 34440 35068 34468 35108
rect 31978 35040 33548 35068
rect 34164 35040 34468 35068
rect 31978 35037 31990 35040
rect 31932 35031 31990 35037
rect 13556 34972 14228 35000
rect 15964 35003 16022 35009
rect 13556 34944 13584 34972
rect 15964 34969 15976 35003
rect 16010 35000 16022 35003
rect 16010 34972 16344 35000
rect 16010 34969 16022 34972
rect 15964 34963 16022 34969
rect 1118 34892 1124 34944
rect 1176 34932 1182 34944
rect 3050 34932 3056 34944
rect 1176 34904 3056 34932
rect 1176 34892 1182 34904
rect 3050 34892 3056 34904
rect 3108 34892 3114 34944
rect 3789 34935 3847 34941
rect 3789 34901 3801 34935
rect 3835 34932 3847 34935
rect 3878 34932 3884 34944
rect 3835 34904 3884 34932
rect 3835 34901 3847 34904
rect 3789 34895 3847 34901
rect 3878 34892 3884 34904
rect 3936 34892 3942 34944
rect 5902 34892 5908 34944
rect 5960 34892 5966 34944
rect 7374 34892 7380 34944
rect 7432 34892 7438 34944
rect 11330 34892 11336 34944
rect 11388 34892 11394 34944
rect 12066 34892 12072 34944
rect 12124 34892 12130 34944
rect 13538 34892 13544 34944
rect 13596 34892 13602 34944
rect 14734 34892 14740 34944
rect 14792 34892 14798 34944
rect 16316 34941 16344 34972
rect 16758 34960 16764 35012
rect 16816 34960 16822 35012
rect 17988 35003 18046 35009
rect 17988 34969 18000 35003
rect 18034 35000 18046 35003
rect 18966 35000 18972 35012
rect 18034 34972 18972 35000
rect 18034 34969 18046 34972
rect 17988 34963 18046 34969
rect 18966 34960 18972 34972
rect 19024 34960 19030 35012
rect 20162 34960 20168 35012
rect 20220 35000 20226 35012
rect 20358 35003 20416 35009
rect 20358 35000 20370 35003
rect 20220 34972 20370 35000
rect 20220 34960 20226 34972
rect 20358 34969 20370 34972
rect 20404 34969 20416 35003
rect 20358 34963 20416 34969
rect 22094 34960 22100 35012
rect 22152 35000 22158 35012
rect 22290 35003 22348 35009
rect 22290 35000 22302 35003
rect 22152 34972 22302 35000
rect 22152 34960 22158 34972
rect 22290 34969 22302 34972
rect 22336 34969 22348 35003
rect 22290 34963 22348 34969
rect 23100 35003 23158 35009
rect 23100 34969 23112 35003
rect 23146 35000 23158 35003
rect 23934 35000 23940 35012
rect 23146 34972 23940 35000
rect 23146 34969 23158 34972
rect 23100 34963 23158 34969
rect 23934 34960 23940 34972
rect 23992 34960 23998 35012
rect 25992 35003 26050 35009
rect 25992 34969 26004 35003
rect 26038 35000 26050 35003
rect 26142 35000 26148 35012
rect 26038 34972 26148 35000
rect 26038 34969 26050 34972
rect 25992 34963 26050 34969
rect 26142 34960 26148 34972
rect 26200 34960 26206 35012
rect 26780 35003 26838 35009
rect 26780 34969 26792 35003
rect 26826 35000 26838 35003
rect 27430 35000 27436 35012
rect 26826 34972 27436 35000
rect 26826 34969 26838 34972
rect 26780 34963 26838 34969
rect 27430 34960 27436 34972
rect 27488 34960 27494 35012
rect 28252 35003 28310 35009
rect 28252 34969 28264 35003
rect 28298 35000 28310 35003
rect 28534 35000 28540 35012
rect 28298 34972 28540 35000
rect 28298 34969 28310 34972
rect 28252 34963 28310 34969
rect 28534 34960 28540 34972
rect 28592 34960 28598 35012
rect 30098 35009 30104 35012
rect 30092 34963 30104 35009
rect 30098 34960 30104 34963
rect 30156 34960 30162 35012
rect 31386 34960 31392 35012
rect 31444 35000 31450 35012
rect 34164 35000 34192 35040
rect 34514 35028 34520 35080
rect 34572 35028 34578 35080
rect 34790 35028 34796 35080
rect 34848 35028 34854 35080
rect 31444 34972 34192 35000
rect 34272 35003 34330 35009
rect 31444 34960 31450 34972
rect 34272 34969 34284 35003
rect 34318 35000 34330 35003
rect 34698 35000 34704 35012
rect 34318 34972 34704 35000
rect 34318 34969 34330 34972
rect 34272 34963 34330 34969
rect 34698 34960 34704 34972
rect 34756 34960 34762 35012
rect 35345 35003 35403 35009
rect 35345 34969 35357 35003
rect 35391 35000 35403 35003
rect 35618 35000 35624 35012
rect 35391 34972 35624 35000
rect 35391 34969 35403 34972
rect 35345 34963 35403 34969
rect 35618 34960 35624 34972
rect 35676 34960 35682 35012
rect 16301 34935 16359 34941
rect 16301 34901 16313 34935
rect 16347 34901 16359 34935
rect 16301 34895 16359 34901
rect 16850 34892 16856 34944
rect 16908 34892 16914 34944
rect 18414 34892 18420 34944
rect 18472 34892 18478 34944
rect 21174 34892 21180 34944
rect 21232 34892 21238 34944
rect 24210 34892 24216 34944
rect 24268 34892 24274 34944
rect 24854 34892 24860 34944
rect 24912 34892 24918 34944
rect 27890 34892 27896 34944
rect 27948 34892 27954 34944
rect 31202 34892 31208 34944
rect 31260 34892 31266 34944
rect 32122 34892 32128 34944
rect 32180 34932 32186 34944
rect 33137 34935 33195 34941
rect 33137 34932 33149 34935
rect 32180 34904 33149 34932
rect 32180 34892 32186 34904
rect 33137 34901 33149 34904
rect 33183 34901 33195 34935
rect 33137 34895 33195 34901
rect 34146 34892 34152 34944
rect 34204 34932 34210 34944
rect 35866 34932 35894 35108
rect 36173 35105 36185 35108
rect 36219 35105 36231 35139
rect 36173 35099 36231 35105
rect 36262 35028 36268 35080
rect 36320 35068 36326 35080
rect 36725 35071 36783 35077
rect 36725 35068 36737 35071
rect 36320 35040 36737 35068
rect 36320 35028 36326 35040
rect 36725 35037 36737 35040
rect 36771 35037 36783 35071
rect 36725 35031 36783 35037
rect 36078 34960 36084 35012
rect 36136 35000 36142 35012
rect 37369 35003 37427 35009
rect 37369 35000 37381 35003
rect 36136 34972 37381 35000
rect 36136 34960 36142 34972
rect 37369 34969 37381 34972
rect 37415 34969 37427 35003
rect 37369 34963 37427 34969
rect 34204 34904 35894 34932
rect 34204 34892 34210 34904
rect 36906 34892 36912 34944
rect 36964 34892 36970 34944
rect 1104 34842 37812 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 37812 34842
rect 1104 34768 37812 34790
rect 1949 34731 2007 34737
rect 1949 34697 1961 34731
rect 1995 34728 2007 34731
rect 2038 34728 2044 34740
rect 1995 34700 2044 34728
rect 1995 34697 2007 34700
rect 1949 34691 2007 34697
rect 2038 34688 2044 34700
rect 2096 34688 2102 34740
rect 2774 34688 2780 34740
rect 2832 34688 2838 34740
rect 5718 34728 5724 34740
rect 5644 34700 5724 34728
rect 2682 34660 2688 34672
rect 1964 34632 2688 34660
rect 1964 34604 1992 34632
rect 2682 34620 2688 34632
rect 2740 34660 2746 34672
rect 5644 34669 5672 34700
rect 5718 34688 5724 34700
rect 5776 34688 5782 34740
rect 5902 34688 5908 34740
rect 5960 34728 5966 34740
rect 5960 34700 6408 34728
rect 5960 34688 5966 34700
rect 5629 34663 5687 34669
rect 2740 34632 4200 34660
rect 2740 34620 2746 34632
rect 1946 34552 1952 34604
rect 2004 34552 2010 34604
rect 2130 34552 2136 34604
rect 2188 34552 2194 34604
rect 3878 34552 3884 34604
rect 3936 34601 3942 34604
rect 4172 34601 4200 34632
rect 5629 34629 5641 34663
rect 5675 34629 5687 34663
rect 5629 34623 5687 34629
rect 3936 34592 3948 34601
rect 4157 34595 4215 34601
rect 3936 34564 3981 34592
rect 3936 34555 3948 34564
rect 4157 34561 4169 34595
rect 4203 34561 4215 34595
rect 4157 34555 4215 34561
rect 3936 34552 3942 34555
rect 5994 34552 6000 34604
rect 6052 34552 6058 34604
rect 6380 34601 6408 34700
rect 7374 34688 7380 34740
rect 7432 34688 7438 34740
rect 8757 34731 8815 34737
rect 8757 34697 8769 34731
rect 8803 34728 8815 34731
rect 8846 34728 8852 34740
rect 8803 34700 8852 34728
rect 8803 34697 8815 34700
rect 8757 34691 8815 34697
rect 8846 34688 8852 34700
rect 8904 34688 8910 34740
rect 8938 34688 8944 34740
rect 8996 34688 9002 34740
rect 9677 34731 9735 34737
rect 9677 34728 9689 34731
rect 9416 34700 9689 34728
rect 7392 34601 7420 34688
rect 9416 34669 9444 34700
rect 9677 34697 9689 34700
rect 9723 34728 9735 34731
rect 11054 34728 11060 34740
rect 9723 34700 11060 34728
rect 9723 34697 9735 34700
rect 9677 34691 9735 34697
rect 11054 34688 11060 34700
rect 11112 34688 11118 34740
rect 11238 34688 11244 34740
rect 11296 34728 11302 34740
rect 11517 34731 11575 34737
rect 11517 34728 11529 34731
rect 11296 34700 11529 34728
rect 11296 34688 11302 34700
rect 11517 34697 11529 34700
rect 11563 34697 11575 34731
rect 11517 34691 11575 34697
rect 12158 34688 12164 34740
rect 12216 34688 12222 34740
rect 14734 34688 14740 34740
rect 14792 34688 14798 34740
rect 15286 34688 15292 34740
rect 15344 34728 15350 34740
rect 15344 34700 15608 34728
rect 15344 34688 15350 34700
rect 9401 34663 9459 34669
rect 9401 34629 9413 34663
rect 9447 34629 9459 34663
rect 11330 34660 11336 34672
rect 9401 34623 9459 34629
rect 9600 34632 11336 34660
rect 6365 34595 6423 34601
rect 6365 34561 6377 34595
rect 6411 34561 6423 34595
rect 6365 34555 6423 34561
rect 7377 34595 7435 34601
rect 7377 34561 7389 34595
rect 7423 34561 7435 34595
rect 7377 34555 7435 34561
rect 9600 34536 9628 34632
rect 11330 34620 11336 34632
rect 11388 34660 11394 34672
rect 13538 34660 13544 34672
rect 11388 34632 13544 34660
rect 11388 34620 11394 34632
rect 13538 34620 13544 34632
rect 13596 34660 13602 34672
rect 13596 34632 14688 34660
rect 13596 34620 13602 34632
rect 10134 34552 10140 34604
rect 10192 34552 10198 34604
rect 10594 34552 10600 34604
rect 10652 34552 10658 34604
rect 12066 34592 12072 34604
rect 11716 34564 12072 34592
rect 1489 34527 1547 34533
rect 1489 34493 1501 34527
rect 1535 34524 1547 34527
rect 2958 34524 2964 34536
rect 1535 34496 2964 34524
rect 1535 34493 1547 34496
rect 1489 34487 1547 34493
rect 2958 34484 2964 34496
rect 3016 34484 3022 34536
rect 8202 34484 8208 34536
rect 8260 34484 8266 34536
rect 9582 34484 9588 34536
rect 9640 34484 9646 34536
rect 1857 34459 1915 34465
rect 1857 34425 1869 34459
rect 1903 34456 1915 34459
rect 2590 34456 2596 34468
rect 1903 34428 2596 34456
rect 1903 34425 1915 34428
rect 1857 34419 1915 34425
rect 2590 34416 2596 34428
rect 2648 34456 2654 34468
rect 2685 34459 2743 34465
rect 2685 34456 2697 34459
rect 2648 34428 2697 34456
rect 2648 34416 2654 34428
rect 2685 34425 2697 34428
rect 2731 34425 2743 34459
rect 2685 34419 2743 34425
rect 9125 34459 9183 34465
rect 9125 34425 9137 34459
rect 9171 34456 9183 34459
rect 9214 34456 9220 34468
rect 9171 34428 9220 34456
rect 9171 34425 9183 34428
rect 9125 34419 9183 34425
rect 9214 34416 9220 34428
rect 9272 34416 9278 34468
rect 11054 34416 11060 34468
rect 11112 34416 11118 34468
rect 11716 34465 11744 34564
rect 12066 34552 12072 34564
rect 12124 34592 12130 34604
rect 12713 34595 12771 34601
rect 12713 34592 12725 34595
rect 12124 34564 12725 34592
rect 12124 34552 12130 34564
rect 12713 34561 12725 34564
rect 12759 34561 12771 34595
rect 12713 34555 12771 34561
rect 14389 34595 14447 34601
rect 14389 34561 14401 34595
rect 14435 34592 14447 34595
rect 14550 34592 14556 34604
rect 14435 34564 14556 34592
rect 14435 34561 14447 34564
rect 14389 34555 14447 34561
rect 14550 34552 14556 34564
rect 14608 34552 14614 34604
rect 14660 34601 14688 34632
rect 14645 34595 14703 34601
rect 14645 34561 14657 34595
rect 14691 34561 14703 34595
rect 14752 34592 14780 34688
rect 15580 34669 15608 34700
rect 16850 34688 16856 34740
rect 16908 34688 16914 34740
rect 17770 34688 17776 34740
rect 17828 34688 17834 34740
rect 18966 34688 18972 34740
rect 19024 34688 19030 34740
rect 19889 34731 19947 34737
rect 19889 34697 19901 34731
rect 19935 34728 19947 34731
rect 19978 34728 19984 34740
rect 19935 34700 19984 34728
rect 19935 34697 19947 34700
rect 19889 34691 19947 34697
rect 19978 34688 19984 34700
rect 20036 34688 20042 34740
rect 20162 34688 20168 34740
rect 20220 34688 20226 34740
rect 23934 34688 23940 34740
rect 23992 34688 23998 34740
rect 24026 34688 24032 34740
rect 24084 34688 24090 34740
rect 24210 34688 24216 34740
rect 24268 34688 24274 34740
rect 24762 34688 24768 34740
rect 24820 34688 24826 34740
rect 24854 34688 24860 34740
rect 24912 34728 24918 34740
rect 24912 34700 25544 34728
rect 24912 34688 24918 34700
rect 15565 34663 15623 34669
rect 15565 34629 15577 34663
rect 15611 34629 15623 34663
rect 15565 34623 15623 34629
rect 15197 34595 15255 34601
rect 15197 34592 15209 34595
rect 14752 34564 15209 34592
rect 14645 34555 14703 34561
rect 15197 34561 15209 34564
rect 15243 34561 15255 34595
rect 16868 34592 16896 34688
rect 17037 34595 17095 34601
rect 17037 34592 17049 34595
rect 16868 34564 17049 34592
rect 15197 34555 15255 34561
rect 17037 34561 17049 34564
rect 17083 34561 17095 34595
rect 17037 34555 17095 34561
rect 11977 34527 12035 34533
rect 11977 34493 11989 34527
rect 12023 34493 12035 34527
rect 11977 34487 12035 34493
rect 11701 34459 11759 34465
rect 11701 34425 11713 34459
rect 11747 34425 11759 34459
rect 11701 34419 11759 34425
rect 7006 34348 7012 34400
rect 7064 34348 7070 34400
rect 8018 34348 8024 34400
rect 8076 34348 8082 34400
rect 11072 34388 11100 34416
rect 11992 34388 12020 34487
rect 16850 34484 16856 34536
rect 16908 34484 16914 34536
rect 17681 34527 17739 34533
rect 17681 34493 17693 34527
rect 17727 34524 17739 34527
rect 18325 34527 18383 34533
rect 18325 34524 18337 34527
rect 17727 34496 18337 34524
rect 17727 34493 17739 34496
rect 17681 34487 17739 34493
rect 18325 34493 18337 34496
rect 18371 34493 18383 34527
rect 18325 34487 18383 34493
rect 18506 34484 18512 34536
rect 18564 34484 18570 34536
rect 19245 34527 19303 34533
rect 19245 34524 19257 34527
rect 18800 34496 19257 34524
rect 18414 34416 18420 34468
rect 18472 34456 18478 34468
rect 18800 34465 18828 34496
rect 19245 34493 19257 34496
rect 19291 34493 19303 34527
rect 19245 34487 19303 34493
rect 19981 34527 20039 34533
rect 19981 34493 19993 34527
rect 20027 34524 20039 34527
rect 20180 34524 20208 34688
rect 20441 34663 20499 34669
rect 20441 34629 20453 34663
rect 20487 34660 20499 34663
rect 20809 34663 20867 34669
rect 20809 34660 20821 34663
rect 20487 34632 20821 34660
rect 20487 34629 20499 34632
rect 20441 34623 20499 34629
rect 20809 34629 20821 34632
rect 20855 34660 20867 34663
rect 22370 34660 22376 34672
rect 20855 34632 22376 34660
rect 20855 34629 20867 34632
rect 20809 34623 20867 34629
rect 22370 34620 22376 34632
rect 22428 34620 22434 34672
rect 21174 34552 21180 34604
rect 21232 34592 21238 34604
rect 21821 34595 21879 34601
rect 21821 34592 21833 34595
rect 21232 34564 21833 34592
rect 21232 34552 21238 34564
rect 21821 34561 21833 34564
rect 21867 34561 21879 34595
rect 21821 34555 21879 34561
rect 21910 34552 21916 34604
rect 21968 34592 21974 34604
rect 22557 34595 22615 34601
rect 22557 34592 22569 34595
rect 21968 34564 22569 34592
rect 21968 34552 21974 34564
rect 22557 34561 22569 34564
rect 22603 34561 22615 34595
rect 22557 34555 22615 34561
rect 23382 34552 23388 34604
rect 23440 34552 23446 34604
rect 21928 34524 21956 34552
rect 20027 34496 20208 34524
rect 21744 34496 21956 34524
rect 22465 34527 22523 34533
rect 20027 34493 20039 34496
rect 19981 34487 20039 34493
rect 18785 34459 18843 34465
rect 18785 34456 18797 34459
rect 18472 34428 18797 34456
rect 18472 34416 18478 34428
rect 18785 34425 18797 34428
rect 18831 34425 18843 34459
rect 18785 34419 18843 34425
rect 20165 34459 20223 34465
rect 20165 34425 20177 34459
rect 20211 34456 20223 34459
rect 21744 34456 21772 34496
rect 22465 34493 22477 34527
rect 22511 34524 22523 34527
rect 23109 34527 23167 34533
rect 23109 34524 23121 34527
rect 22511 34496 23121 34524
rect 22511 34493 22523 34496
rect 22465 34487 22523 34493
rect 23109 34493 23121 34496
rect 23155 34493 23167 34527
rect 23952 34524 23980 34688
rect 24228 34601 24256 34688
rect 25516 34601 25544 34700
rect 26142 34688 26148 34740
rect 26200 34728 26206 34740
rect 26237 34731 26295 34737
rect 26237 34728 26249 34731
rect 26200 34700 26249 34728
rect 26200 34688 26206 34700
rect 26237 34697 26249 34700
rect 26283 34697 26295 34731
rect 26237 34691 26295 34697
rect 27522 34688 27528 34740
rect 27580 34728 27586 34740
rect 27617 34731 27675 34737
rect 27617 34728 27629 34731
rect 27580 34700 27629 34728
rect 27580 34688 27586 34700
rect 27617 34697 27629 34700
rect 27663 34697 27675 34731
rect 27617 34691 27675 34697
rect 27890 34688 27896 34740
rect 27948 34688 27954 34740
rect 28534 34688 28540 34740
rect 28592 34688 28598 34740
rect 29086 34688 29092 34740
rect 29144 34688 29150 34740
rect 34606 34728 34612 34740
rect 32416 34700 34612 34728
rect 24213 34595 24271 34601
rect 24213 34561 24225 34595
rect 24259 34561 24271 34595
rect 24213 34555 24271 34561
rect 25501 34595 25559 34601
rect 25501 34561 25513 34595
rect 25547 34561 25559 34595
rect 25501 34555 25559 34561
rect 25608 34564 26740 34592
rect 24857 34527 24915 34533
rect 24857 34524 24869 34527
rect 23952 34496 24869 34524
rect 23109 34487 23167 34493
rect 24857 34493 24869 34496
rect 24903 34493 24915 34527
rect 24857 34487 24915 34493
rect 25317 34527 25375 34533
rect 25317 34493 25329 34527
rect 25363 34524 25375 34527
rect 25406 34524 25412 34536
rect 25363 34496 25412 34524
rect 25363 34493 25375 34496
rect 25317 34487 25375 34493
rect 25406 34484 25412 34496
rect 25464 34524 25470 34536
rect 25608 34524 25636 34564
rect 26712 34536 26740 34564
rect 27062 34552 27068 34604
rect 27120 34552 27126 34604
rect 27801 34595 27859 34601
rect 27801 34561 27813 34595
rect 27847 34592 27859 34595
rect 27908 34592 27936 34688
rect 28353 34663 28411 34669
rect 28353 34629 28365 34663
rect 28399 34660 28411 34663
rect 29104 34660 29132 34688
rect 28399 34632 29132 34660
rect 28399 34629 28411 34632
rect 28353 34623 28411 34629
rect 27847 34564 27936 34592
rect 30469 34595 30527 34601
rect 27847 34561 27859 34564
rect 27801 34555 27859 34561
rect 30469 34561 30481 34595
rect 30515 34592 30527 34595
rect 31662 34592 31668 34604
rect 30515 34564 31668 34592
rect 30515 34561 30527 34564
rect 30469 34555 30527 34561
rect 31662 34552 31668 34564
rect 31720 34552 31726 34604
rect 31938 34552 31944 34604
rect 31996 34552 32002 34604
rect 25464 34496 25636 34524
rect 26145 34527 26203 34533
rect 25464 34484 25470 34496
rect 26145 34493 26157 34527
rect 26191 34524 26203 34527
rect 26602 34524 26608 34536
rect 26191 34496 26608 34524
rect 26191 34493 26203 34496
rect 26145 34487 26203 34493
rect 26602 34484 26608 34496
rect 26660 34484 26666 34536
rect 26694 34484 26700 34536
rect 26752 34484 26758 34536
rect 20211 34428 21772 34456
rect 25041 34459 25099 34465
rect 20211 34425 20223 34428
rect 20165 34419 20223 34425
rect 25041 34425 25053 34459
rect 25087 34456 25099 34459
rect 25958 34456 25964 34468
rect 25087 34428 25964 34456
rect 25087 34425 25099 34428
rect 25041 34419 25099 34425
rect 25958 34416 25964 34428
rect 26016 34416 26022 34468
rect 26421 34459 26479 34465
rect 26421 34425 26433 34459
rect 26467 34456 26479 34459
rect 27080 34456 27108 34552
rect 28997 34527 29055 34533
rect 28997 34493 29009 34527
rect 29043 34524 29055 34527
rect 29638 34524 29644 34536
rect 29043 34496 29644 34524
rect 29043 34493 29055 34496
rect 28997 34487 29055 34493
rect 29638 34484 29644 34496
rect 29696 34484 29702 34536
rect 30009 34527 30067 34533
rect 30009 34493 30021 34527
rect 30055 34524 30067 34527
rect 31386 34524 31392 34536
rect 30055 34496 31392 34524
rect 30055 34493 30067 34496
rect 30009 34487 30067 34493
rect 31386 34484 31392 34496
rect 31444 34484 31450 34536
rect 31481 34527 31539 34533
rect 31481 34493 31493 34527
rect 31527 34524 31539 34527
rect 32416 34524 32444 34700
rect 34606 34688 34612 34700
rect 34664 34688 34670 34740
rect 33318 34620 33324 34672
rect 33376 34660 33382 34672
rect 34514 34660 34520 34672
rect 33376 34632 34520 34660
rect 33376 34620 33382 34632
rect 34514 34620 34520 34632
rect 34572 34660 34578 34672
rect 35342 34660 35348 34672
rect 34572 34632 35348 34660
rect 34572 34620 34578 34632
rect 35342 34620 35348 34632
rect 35400 34660 35406 34672
rect 35400 34632 36860 34660
rect 35400 34620 35406 34632
rect 32950 34552 32956 34604
rect 33008 34592 33014 34604
rect 33238 34595 33296 34601
rect 33238 34592 33250 34595
rect 33008 34564 33250 34592
rect 33008 34552 33014 34564
rect 33238 34561 33250 34564
rect 33284 34561 33296 34595
rect 33336 34592 33364 34620
rect 33505 34595 33563 34601
rect 33505 34592 33517 34595
rect 33336 34564 33517 34592
rect 33238 34555 33296 34561
rect 33505 34561 33517 34564
rect 33551 34561 33563 34595
rect 33505 34555 33563 34561
rect 34054 34552 34060 34604
rect 34112 34552 34118 34604
rect 36561 34595 36619 34601
rect 36561 34561 36573 34595
rect 36607 34592 36619 34595
rect 36722 34592 36728 34604
rect 36607 34564 36728 34592
rect 36607 34561 36619 34564
rect 36561 34555 36619 34561
rect 36722 34552 36728 34564
rect 36780 34552 36786 34604
rect 36832 34601 36860 34632
rect 36817 34595 36875 34601
rect 36817 34561 36829 34595
rect 36863 34561 36875 34595
rect 36817 34555 36875 34561
rect 31527 34496 32444 34524
rect 31527 34493 31539 34496
rect 31481 34487 31539 34493
rect 34330 34484 34336 34536
rect 34388 34484 34394 34536
rect 34514 34484 34520 34536
rect 34572 34524 34578 34536
rect 34572 34496 35480 34524
rect 34572 34484 34578 34496
rect 35452 34465 35480 34496
rect 26467 34428 27108 34456
rect 28721 34459 28779 34465
rect 26467 34425 26479 34428
rect 26421 34419 26479 34425
rect 28721 34425 28733 34459
rect 28767 34456 28779 34459
rect 35437 34459 35495 34465
rect 28767 34428 32628 34456
rect 28767 34425 28779 34428
rect 28721 34419 28779 34425
rect 12066 34388 12072 34400
rect 11072 34360 12072 34388
rect 12066 34348 12072 34360
rect 12124 34348 12130 34400
rect 13262 34348 13268 34400
rect 13320 34348 13326 34400
rect 30926 34348 30932 34400
rect 30984 34388 30990 34400
rect 32125 34391 32183 34397
rect 32125 34388 32137 34391
rect 30984 34360 32137 34388
rect 30984 34348 30990 34360
rect 32125 34357 32137 34360
rect 32171 34357 32183 34391
rect 32600 34388 32628 34428
rect 35437 34425 35449 34459
rect 35483 34425 35495 34459
rect 35437 34419 35495 34425
rect 34146 34388 34152 34400
rect 32600 34360 34152 34388
rect 32125 34351 32183 34357
rect 34146 34348 34152 34360
rect 34204 34348 34210 34400
rect 1104 34298 37812 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 37812 34298
rect 1104 34224 37812 34246
rect 3605 34187 3663 34193
rect 3605 34153 3617 34187
rect 3651 34184 3663 34187
rect 3694 34184 3700 34196
rect 3651 34156 3700 34184
rect 3651 34153 3663 34156
rect 3605 34147 3663 34153
rect 3694 34144 3700 34156
rect 3752 34144 3758 34196
rect 5905 34187 5963 34193
rect 5905 34153 5917 34187
rect 5951 34184 5963 34187
rect 5994 34184 6000 34196
rect 5951 34156 6000 34184
rect 5951 34153 5963 34156
rect 5905 34147 5963 34153
rect 5994 34144 6000 34156
rect 6052 34144 6058 34196
rect 6273 34187 6331 34193
rect 6273 34153 6285 34187
rect 6319 34184 6331 34187
rect 6546 34184 6552 34196
rect 6319 34156 6552 34184
rect 6319 34153 6331 34156
rect 6273 34147 6331 34153
rect 6546 34144 6552 34156
rect 6604 34144 6610 34196
rect 7650 34144 7656 34196
rect 7708 34144 7714 34196
rect 8202 34144 8208 34196
rect 8260 34184 8266 34196
rect 8573 34187 8631 34193
rect 8573 34184 8585 34187
rect 8260 34156 8585 34184
rect 8260 34144 8266 34156
rect 8573 34153 8585 34156
rect 8619 34153 8631 34187
rect 8573 34147 8631 34153
rect 10594 34144 10600 34196
rect 10652 34144 10658 34196
rect 12066 34144 12072 34196
rect 12124 34184 12130 34196
rect 12124 34156 12756 34184
rect 12124 34144 12130 34156
rect 7561 34119 7619 34125
rect 7561 34085 7573 34119
rect 7607 34116 7619 34119
rect 8220 34116 8248 34144
rect 7607 34088 8248 34116
rect 7607 34085 7619 34088
rect 7561 34079 7619 34085
rect 2590 34008 2596 34060
rect 2648 34048 2654 34060
rect 2961 34051 3019 34057
rect 2961 34048 2973 34051
rect 2648 34020 2973 34048
rect 2648 34008 2654 34020
rect 2961 34017 2973 34020
rect 3007 34017 3019 34051
rect 2961 34011 3019 34017
rect 4246 34008 4252 34060
rect 4304 34008 4310 34060
rect 4798 34008 4804 34060
rect 4856 34048 4862 34060
rect 5258 34048 5264 34060
rect 4856 34020 5264 34048
rect 4856 34008 4862 34020
rect 5258 34008 5264 34020
rect 5316 34008 5322 34060
rect 6917 34051 6975 34057
rect 6917 34017 6929 34051
rect 6963 34048 6975 34051
rect 7006 34048 7012 34060
rect 6963 34020 7012 34048
rect 6963 34017 6975 34020
rect 6917 34011 6975 34017
rect 7006 34008 7012 34020
rect 7064 34008 7070 34060
rect 8018 34008 8024 34060
rect 8076 34008 8082 34060
rect 9214 34008 9220 34060
rect 9272 34048 9278 34060
rect 12728 34057 12756 34156
rect 13170 34144 13176 34196
rect 13228 34144 13234 34196
rect 14182 34144 14188 34196
rect 14240 34184 14246 34196
rect 14734 34184 14740 34196
rect 14240 34156 14740 34184
rect 14240 34144 14246 34156
rect 14734 34144 14740 34156
rect 14792 34184 14798 34196
rect 15105 34187 15163 34193
rect 15105 34184 15117 34187
rect 14792 34156 15117 34184
rect 14792 34144 14798 34156
rect 15105 34153 15117 34156
rect 15151 34153 15163 34187
rect 15105 34147 15163 34153
rect 21913 34187 21971 34193
rect 21913 34153 21925 34187
rect 21959 34184 21971 34187
rect 22094 34184 22100 34196
rect 21959 34156 22100 34184
rect 21959 34153 21971 34156
rect 21913 34147 21971 34153
rect 22094 34144 22100 34156
rect 22152 34144 22158 34196
rect 22922 34144 22928 34196
rect 22980 34184 22986 34196
rect 23017 34187 23075 34193
rect 23017 34184 23029 34187
rect 22980 34156 23029 34184
rect 22980 34144 22986 34156
rect 23017 34153 23029 34156
rect 23063 34153 23075 34187
rect 23017 34147 23075 34153
rect 25406 34144 25412 34196
rect 25464 34144 25470 34196
rect 25958 34144 25964 34196
rect 26016 34184 26022 34196
rect 26053 34187 26111 34193
rect 26053 34184 26065 34187
rect 26016 34156 26065 34184
rect 26016 34144 26022 34156
rect 26053 34153 26065 34156
rect 26099 34153 26111 34187
rect 26053 34147 26111 34153
rect 27430 34144 27436 34196
rect 27488 34144 27494 34196
rect 30098 34144 30104 34196
rect 30156 34144 30162 34196
rect 32398 34184 32404 34196
rect 30208 34156 32404 34184
rect 13081 34119 13139 34125
rect 13081 34085 13093 34119
rect 13127 34116 13139 34119
rect 13906 34116 13912 34128
rect 13127 34088 13912 34116
rect 13127 34085 13139 34088
rect 13081 34079 13139 34085
rect 13906 34076 13912 34088
rect 13964 34116 13970 34128
rect 14093 34119 14151 34125
rect 14093 34116 14105 34119
rect 13964 34088 14105 34116
rect 13964 34076 13970 34088
rect 14093 34085 14105 34088
rect 14139 34085 14151 34119
rect 14093 34079 14151 34085
rect 22005 34119 22063 34125
rect 22005 34085 22017 34119
rect 22051 34116 22063 34119
rect 23382 34116 23388 34128
rect 22051 34088 23388 34116
rect 22051 34085 22063 34088
rect 22005 34079 22063 34085
rect 23382 34076 23388 34088
rect 23440 34076 23446 34128
rect 9953 34051 10011 34057
rect 9953 34048 9965 34051
rect 9272 34020 9965 34048
rect 9272 34008 9278 34020
rect 9953 34017 9965 34020
rect 9999 34017 10011 34051
rect 9953 34011 10011 34017
rect 12713 34051 12771 34057
rect 12713 34017 12725 34051
rect 12759 34017 12771 34051
rect 12713 34011 12771 34017
rect 13262 34008 13268 34060
rect 13320 34008 13326 34060
rect 15010 34008 15016 34060
rect 15068 34048 15074 34060
rect 15657 34051 15715 34057
rect 15657 34048 15669 34051
rect 15068 34020 15669 34048
rect 15068 34008 15074 34020
rect 15657 34017 15669 34020
rect 15703 34017 15715 34051
rect 15657 34011 15715 34017
rect 22370 34008 22376 34060
rect 22428 34048 22434 34060
rect 22741 34051 22799 34057
rect 22741 34048 22753 34051
rect 22428 34020 22753 34048
rect 22428 34008 22434 34020
rect 22741 34017 22753 34020
rect 22787 34048 22799 34051
rect 25424 34048 25452 34144
rect 27617 34119 27675 34125
rect 27617 34085 27629 34119
rect 27663 34085 27675 34119
rect 27617 34079 27675 34085
rect 22787 34020 25452 34048
rect 22787 34017 22799 34020
rect 22741 34011 22799 34017
rect 26602 34008 26608 34060
rect 26660 34008 26666 34060
rect 27632 34048 27660 34079
rect 30006 34076 30012 34128
rect 30064 34076 30070 34128
rect 28718 34048 28724 34060
rect 27632 34020 28724 34048
rect 28718 34008 28724 34020
rect 28776 34008 28782 34060
rect 29638 34008 29644 34060
rect 29696 34048 29702 34060
rect 30208 34048 30236 34156
rect 32398 34144 32404 34156
rect 32456 34184 32462 34196
rect 32769 34187 32827 34193
rect 32769 34184 32781 34187
rect 32456 34156 32781 34184
rect 32456 34144 32462 34156
rect 32769 34153 32781 34156
rect 32815 34184 32827 34187
rect 35250 34184 35256 34196
rect 32815 34156 35256 34184
rect 32815 34153 32827 34156
rect 32769 34147 32827 34153
rect 35250 34144 35256 34156
rect 35308 34144 35314 34196
rect 35345 34187 35403 34193
rect 35345 34153 35357 34187
rect 35391 34184 35403 34187
rect 35434 34184 35440 34196
rect 35391 34156 35440 34184
rect 35391 34153 35403 34156
rect 35345 34147 35403 34153
rect 35434 34144 35440 34156
rect 35492 34144 35498 34196
rect 35621 34119 35679 34125
rect 31128 34088 35480 34116
rect 31128 34057 31156 34088
rect 29696 34020 30236 34048
rect 31113 34051 31171 34057
rect 29696 34008 29702 34020
rect 31113 34017 31125 34051
rect 31159 34017 31171 34051
rect 32033 34051 32091 34057
rect 32033 34048 32045 34051
rect 31113 34011 31171 34017
rect 31588 34020 32045 34048
rect 2685 33983 2743 33989
rect 2685 33949 2697 33983
rect 2731 33980 2743 33983
rect 3234 33980 3240 33992
rect 2731 33952 3240 33980
rect 2731 33949 2743 33952
rect 2685 33943 2743 33949
rect 3234 33940 3240 33952
rect 3292 33940 3298 33992
rect 3786 33940 3792 33992
rect 3844 33940 3850 33992
rect 4890 33940 4896 33992
rect 4948 33980 4954 33992
rect 6822 33980 6828 33992
rect 4948 33952 6828 33980
rect 4948 33940 4954 33952
rect 6822 33940 6828 33952
rect 6880 33980 6886 33992
rect 7193 33983 7251 33989
rect 7193 33980 7205 33983
rect 6880 33952 7205 33980
rect 6880 33940 6886 33952
rect 7193 33949 7205 33952
rect 7239 33949 7251 33983
rect 7193 33943 7251 33949
rect 13909 33983 13967 33989
rect 13909 33949 13921 33983
rect 13955 33980 13967 33983
rect 14645 33983 14703 33989
rect 14645 33980 14657 33983
rect 13955 33952 14657 33980
rect 13955 33949 13967 33952
rect 13909 33943 13967 33949
rect 14645 33949 14657 33952
rect 14691 33949 14703 33983
rect 14645 33943 14703 33949
rect 28074 33940 28080 33992
rect 28132 33940 28138 33992
rect 29365 33983 29423 33989
rect 29365 33949 29377 33983
rect 29411 33980 29423 33983
rect 30466 33980 30472 33992
rect 29411 33952 30472 33980
rect 29411 33949 29423 33952
rect 29365 33943 29423 33949
rect 30466 33940 30472 33952
rect 30524 33940 30530 33992
rect 31588 33989 31616 34020
rect 32033 34017 32045 34020
rect 32079 34017 32091 34051
rect 32033 34011 32091 34017
rect 33410 34008 33416 34060
rect 33468 34048 33474 34060
rect 34701 34051 34759 34057
rect 34701 34048 34713 34051
rect 33468 34020 34713 34048
rect 33468 34008 33474 34020
rect 34701 34017 34713 34020
rect 34747 34017 34759 34051
rect 35452 34048 35480 34088
rect 35621 34085 35633 34119
rect 35667 34116 35679 34119
rect 35710 34116 35716 34128
rect 35667 34088 35716 34116
rect 35667 34085 35679 34088
rect 35621 34079 35679 34085
rect 35710 34076 35716 34088
rect 35768 34076 35774 34128
rect 36170 34116 36176 34128
rect 35912 34088 36176 34116
rect 35802 34048 35808 34060
rect 35452 34020 35808 34048
rect 34701 34011 34759 34017
rect 35802 34008 35808 34020
rect 35860 34008 35866 34060
rect 35912 34057 35940 34088
rect 36170 34076 36176 34088
rect 36228 34116 36234 34128
rect 36354 34116 36360 34128
rect 36228 34088 36360 34116
rect 36228 34076 36234 34088
rect 36354 34076 36360 34088
rect 36412 34116 36418 34128
rect 37093 34119 37151 34125
rect 37093 34116 37105 34119
rect 36412 34088 37105 34116
rect 36412 34076 36418 34088
rect 37093 34085 37105 34088
rect 37139 34085 37151 34119
rect 37093 34079 37151 34085
rect 35897 34051 35955 34057
rect 35897 34017 35909 34051
rect 35943 34017 35955 34051
rect 35897 34011 35955 34017
rect 31573 33983 31631 33989
rect 31573 33949 31585 33983
rect 31619 33949 31631 33983
rect 31573 33943 31631 33949
rect 31754 33940 31760 33992
rect 31812 33940 31818 33992
rect 33226 33940 33232 33992
rect 33284 33940 33290 33992
rect 34606 33940 34612 33992
rect 34664 33980 34670 33992
rect 36173 33983 36231 33989
rect 36173 33980 36185 33983
rect 34664 33952 36185 33980
rect 34664 33940 34670 33952
rect 36173 33949 36185 33952
rect 36219 33949 36231 33983
rect 36173 33943 36231 33949
rect 2317 33915 2375 33921
rect 2317 33881 2329 33915
rect 2363 33912 2375 33915
rect 27893 33915 27951 33921
rect 2363 33884 2912 33912
rect 2363 33881 2375 33884
rect 2317 33875 2375 33881
rect 2884 33856 2912 33884
rect 27893 33881 27905 33915
rect 27939 33881 27951 33915
rect 27893 33875 27951 33881
rect 30668 33884 33548 33912
rect 2866 33804 2872 33856
rect 2924 33804 2930 33856
rect 17310 33804 17316 33856
rect 17368 33844 17374 33856
rect 18325 33847 18383 33853
rect 18325 33844 18337 33847
rect 17368 33816 18337 33844
rect 17368 33804 17374 33816
rect 18325 33813 18337 33816
rect 18371 33844 18383 33847
rect 18506 33844 18512 33856
rect 18371 33816 18512 33844
rect 18371 33813 18383 33816
rect 18325 33807 18383 33813
rect 18506 33804 18512 33816
rect 18564 33804 18570 33856
rect 26694 33804 26700 33856
rect 26752 33844 26758 33856
rect 27065 33847 27123 33853
rect 27065 33844 27077 33847
rect 26752 33816 27077 33844
rect 26752 33804 26758 33816
rect 27065 33813 27077 33816
rect 27111 33844 27123 33847
rect 27908 33844 27936 33875
rect 30668 33856 30696 33884
rect 27982 33844 27988 33856
rect 27111 33816 27988 33844
rect 27111 33813 27123 33816
rect 27065 33807 27123 33813
rect 27982 33804 27988 33816
rect 28040 33804 28046 33856
rect 28629 33847 28687 33853
rect 28629 33813 28641 33847
rect 28675 33844 28687 33847
rect 29178 33844 29184 33856
rect 28675 33816 29184 33844
rect 28675 33813 28687 33816
rect 28629 33807 28687 33813
rect 29178 33804 29184 33816
rect 29236 33804 29242 33856
rect 30650 33804 30656 33856
rect 30708 33804 30714 33856
rect 33520 33844 33548 33884
rect 33594 33872 33600 33924
rect 33652 33872 33658 33924
rect 35710 33912 35716 33924
rect 34624 33884 35716 33912
rect 34422 33844 34428 33856
rect 33520 33816 34428 33844
rect 34422 33804 34428 33816
rect 34480 33844 34486 33856
rect 34624 33844 34652 33884
rect 35710 33872 35716 33884
rect 35768 33872 35774 33924
rect 36538 33872 36544 33924
rect 36596 33872 36602 33924
rect 34480 33816 34652 33844
rect 34480 33804 34486 33816
rect 34698 33804 34704 33856
rect 34756 33844 34762 33856
rect 35437 33847 35495 33853
rect 35437 33844 35449 33847
rect 34756 33816 35449 33844
rect 34756 33804 34762 33816
rect 35437 33813 35449 33816
rect 35483 33813 35495 33847
rect 35437 33807 35495 33813
rect 35526 33804 35532 33856
rect 35584 33844 35590 33856
rect 36262 33844 36268 33856
rect 35584 33816 36268 33844
rect 35584 33804 35590 33816
rect 36262 33804 36268 33816
rect 36320 33804 36326 33856
rect 1104 33754 37812 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 37812 33754
rect 1104 33680 37812 33702
rect 5258 33600 5264 33652
rect 5316 33640 5322 33652
rect 5353 33643 5411 33649
rect 5353 33640 5365 33643
rect 5316 33612 5365 33640
rect 5316 33600 5322 33612
rect 5353 33609 5365 33612
rect 5399 33609 5411 33643
rect 5353 33603 5411 33609
rect 6362 33600 6368 33652
rect 6420 33600 6426 33652
rect 6822 33600 6828 33652
rect 6880 33600 6886 33652
rect 12066 33600 12072 33652
rect 12124 33640 12130 33652
rect 13265 33643 13323 33649
rect 13265 33640 13277 33643
rect 12124 33612 13277 33640
rect 12124 33600 12130 33612
rect 13265 33609 13277 33612
rect 13311 33609 13323 33643
rect 13265 33603 13323 33609
rect 2498 33464 2504 33516
rect 2556 33504 2562 33516
rect 2685 33507 2743 33513
rect 2685 33504 2697 33507
rect 2556 33476 2697 33504
rect 2556 33464 2562 33476
rect 2685 33473 2697 33476
rect 2731 33473 2743 33507
rect 2685 33467 2743 33473
rect 2866 33464 2872 33516
rect 2924 33464 2930 33516
rect 4706 33464 4712 33516
rect 4764 33464 4770 33516
rect 6840 33513 6868 33600
rect 6825 33507 6883 33513
rect 6825 33473 6837 33507
rect 6871 33473 6883 33507
rect 6825 33467 6883 33473
rect 2409 33439 2467 33445
rect 2409 33405 2421 33439
rect 2455 33436 2467 33439
rect 2590 33436 2596 33448
rect 2455 33408 2596 33436
rect 2455 33405 2467 33408
rect 2409 33399 2467 33405
rect 2590 33396 2596 33408
rect 2648 33396 2654 33448
rect 3326 33396 3332 33448
rect 3384 33396 3390 33448
rect 5994 33396 6000 33448
rect 6052 33396 6058 33448
rect 13280 33436 13308 33603
rect 13906 33600 13912 33652
rect 13964 33600 13970 33652
rect 14550 33600 14556 33652
rect 14608 33640 14614 33652
rect 14645 33643 14703 33649
rect 14645 33640 14657 33643
rect 14608 33612 14657 33640
rect 14608 33600 14614 33612
rect 14645 33609 14657 33612
rect 14691 33609 14703 33643
rect 16850 33640 16856 33652
rect 14645 33603 14703 33609
rect 15396 33612 16856 33640
rect 13924 33513 13952 33600
rect 13909 33507 13967 33513
rect 13909 33473 13921 33507
rect 13955 33473 13967 33507
rect 13909 33467 13967 33473
rect 14553 33507 14611 33513
rect 14553 33473 14565 33507
rect 14599 33504 14611 33507
rect 14642 33504 14648 33516
rect 14599 33476 14648 33504
rect 14599 33473 14611 33476
rect 14553 33467 14611 33473
rect 14642 33464 14648 33476
rect 14700 33464 14706 33516
rect 15396 33445 15424 33612
rect 16850 33600 16856 33612
rect 16908 33640 16914 33652
rect 17310 33640 17316 33652
rect 16908 33612 17316 33640
rect 16908 33600 16914 33612
rect 17310 33600 17316 33612
rect 17368 33600 17374 33652
rect 28718 33600 28724 33652
rect 28776 33640 28782 33652
rect 28905 33643 28963 33649
rect 28905 33640 28917 33643
rect 28776 33612 28917 33640
rect 28776 33600 28782 33612
rect 28905 33609 28917 33612
rect 28951 33609 28963 33643
rect 28905 33603 28963 33609
rect 29638 33600 29644 33652
rect 29696 33600 29702 33652
rect 31205 33643 31263 33649
rect 31205 33609 31217 33643
rect 31251 33640 31263 33643
rect 31754 33640 31760 33652
rect 31251 33612 31760 33640
rect 31251 33609 31263 33612
rect 31205 33603 31263 33609
rect 31754 33600 31760 33612
rect 31812 33600 31818 33652
rect 33134 33640 33140 33652
rect 31864 33612 33140 33640
rect 27982 33532 27988 33584
rect 28040 33572 28046 33584
rect 28813 33575 28871 33581
rect 28813 33572 28825 33575
rect 28040 33544 28825 33572
rect 28040 33532 28046 33544
rect 28813 33541 28825 33544
rect 28859 33572 28871 33575
rect 29656 33572 29684 33600
rect 28859 33544 29684 33572
rect 30469 33575 30527 33581
rect 28859 33541 28871 33544
rect 28813 33535 28871 33541
rect 30469 33541 30481 33575
rect 30515 33572 30527 33575
rect 31864 33572 31892 33612
rect 33134 33600 33140 33612
rect 33192 33600 33198 33652
rect 35526 33640 35532 33652
rect 33888 33612 35532 33640
rect 30515 33544 31892 33572
rect 30515 33541 30527 33544
rect 30469 33535 30527 33541
rect 31938 33532 31944 33584
rect 31996 33572 32002 33584
rect 32953 33575 33011 33581
rect 32953 33572 32965 33575
rect 31996 33544 32965 33572
rect 31996 33532 32002 33544
rect 32953 33541 32965 33544
rect 32999 33541 33011 33575
rect 32953 33535 33011 33541
rect 28074 33464 28080 33516
rect 28132 33464 28138 33516
rect 29546 33464 29552 33516
rect 29604 33464 29610 33516
rect 29917 33507 29975 33513
rect 29917 33473 29929 33507
rect 29963 33504 29975 33507
rect 30926 33504 30932 33516
rect 29963 33476 30932 33504
rect 29963 33473 29975 33476
rect 29917 33467 29975 33473
rect 30926 33464 30932 33476
rect 30984 33464 30990 33516
rect 31202 33464 31208 33516
rect 31260 33504 31266 33516
rect 31297 33507 31355 33513
rect 31297 33504 31309 33507
rect 31260 33476 31309 33504
rect 31260 33464 31266 33476
rect 31297 33473 31309 33476
rect 31343 33473 31355 33507
rect 31297 33467 31355 33473
rect 32398 33464 32404 33516
rect 32456 33464 32462 33516
rect 32582 33464 32588 33516
rect 32640 33464 32646 33516
rect 15105 33439 15163 33445
rect 15105 33436 15117 33439
rect 13280 33408 15117 33436
rect 15105 33405 15117 33408
rect 15151 33436 15163 33439
rect 15381 33439 15439 33445
rect 15381 33436 15393 33439
rect 15151 33408 15393 33436
rect 15151 33405 15163 33408
rect 15105 33399 15163 33405
rect 15381 33405 15393 33408
rect 15427 33405 15439 33439
rect 15381 33399 15439 33405
rect 6546 33328 6552 33380
rect 6604 33328 6610 33380
rect 14734 33328 14740 33380
rect 14792 33328 14798 33380
rect 28092 33368 28120 33464
rect 30650 33396 30656 33448
rect 30708 33396 30714 33448
rect 31941 33439 31999 33445
rect 31941 33405 31953 33439
rect 31987 33436 31999 33439
rect 33888 33436 33916 33612
rect 35526 33600 35532 33612
rect 35584 33600 35590 33652
rect 35710 33600 35716 33652
rect 35768 33640 35774 33652
rect 35894 33640 35900 33652
rect 35768 33612 35900 33640
rect 35768 33600 35774 33612
rect 35894 33600 35900 33612
rect 35952 33640 35958 33652
rect 36170 33640 36176 33652
rect 35952 33612 36176 33640
rect 35952 33600 35958 33612
rect 36170 33600 36176 33612
rect 36228 33600 36234 33652
rect 35100 33575 35158 33581
rect 35100 33541 35112 33575
rect 35146 33572 35158 33575
rect 36906 33572 36912 33584
rect 35146 33544 36912 33572
rect 35146 33541 35158 33544
rect 35100 33535 35158 33541
rect 36906 33532 36912 33544
rect 36964 33532 36970 33584
rect 33962 33464 33968 33516
rect 34020 33504 34026 33516
rect 34020 33476 35296 33504
rect 34020 33464 34026 33476
rect 31987 33408 33916 33436
rect 35268 33436 35296 33476
rect 35342 33464 35348 33516
rect 35400 33504 35406 33516
rect 35437 33507 35495 33513
rect 35437 33504 35449 33507
rect 35400 33476 35449 33504
rect 35400 33464 35406 33476
rect 35437 33473 35449 33476
rect 35483 33473 35495 33507
rect 35693 33507 35751 33513
rect 35693 33504 35705 33507
rect 35437 33467 35495 33473
rect 35544 33476 35705 33504
rect 35544 33436 35572 33476
rect 35693 33473 35705 33476
rect 35739 33473 35751 33507
rect 35693 33467 35751 33473
rect 35268 33408 35572 33436
rect 31987 33405 31999 33408
rect 31941 33399 31999 33405
rect 33965 33371 34023 33377
rect 33965 33368 33977 33371
rect 28092 33340 33977 33368
rect 33965 33337 33977 33340
rect 34011 33337 34023 33371
rect 33965 33331 34023 33337
rect 4706 33260 4712 33312
rect 4764 33300 4770 33312
rect 5445 33303 5503 33309
rect 5445 33300 5457 33303
rect 4764 33272 5457 33300
rect 4764 33260 4770 33272
rect 5445 33269 5457 33272
rect 5491 33269 5503 33303
rect 5445 33263 5503 33269
rect 33597 33303 33655 33309
rect 33597 33269 33609 33303
rect 33643 33300 33655 33303
rect 34146 33300 34152 33312
rect 33643 33272 34152 33300
rect 33643 33269 33655 33272
rect 33597 33263 33655 33269
rect 34146 33260 34152 33272
rect 34204 33260 34210 33312
rect 34698 33260 34704 33312
rect 34756 33300 34762 33312
rect 36817 33303 36875 33309
rect 36817 33300 36829 33303
rect 34756 33272 36829 33300
rect 34756 33260 34762 33272
rect 36817 33269 36829 33272
rect 36863 33269 36875 33303
rect 36817 33263 36875 33269
rect 1104 33210 37812 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 37812 33210
rect 1104 33136 37812 33158
rect 32490 33056 32496 33108
rect 32548 33056 32554 33108
rect 32950 33056 32956 33108
rect 33008 33096 33014 33108
rect 33045 33099 33103 33105
rect 33045 33096 33057 33099
rect 33008 33068 33057 33096
rect 33008 33056 33014 33068
rect 33045 33065 33057 33068
rect 33091 33065 33103 33099
rect 36078 33096 36084 33108
rect 33045 33059 33103 33065
rect 35866 33068 36084 33096
rect 32398 33028 32404 33040
rect 31220 33000 32404 33028
rect 1578 32920 1584 32972
rect 1636 32920 1642 32972
rect 29178 32920 29184 32972
rect 29236 32960 29242 32972
rect 31220 32969 31248 33000
rect 32398 32988 32404 33000
rect 32456 32988 32462 33040
rect 32766 32988 32772 33040
rect 32824 33028 32830 33040
rect 32861 33031 32919 33037
rect 32861 33028 32873 33031
rect 32824 33000 32873 33028
rect 32824 32988 32830 33000
rect 32861 32997 32873 33000
rect 32907 32997 32919 33031
rect 32861 32991 32919 32997
rect 33318 32988 33324 33040
rect 33376 33028 33382 33040
rect 35069 33031 35127 33037
rect 35069 33028 35081 33031
rect 33376 33000 35081 33028
rect 33376 32988 33382 33000
rect 35069 32997 35081 33000
rect 35115 32997 35127 33031
rect 35069 32991 35127 32997
rect 29641 32963 29699 32969
rect 29641 32960 29653 32963
rect 29236 32932 29653 32960
rect 29236 32920 29242 32932
rect 29641 32929 29653 32932
rect 29687 32929 29699 32963
rect 29641 32923 29699 32929
rect 31205 32963 31263 32969
rect 31205 32929 31217 32963
rect 31251 32929 31263 32963
rect 31205 32923 31263 32929
rect 31757 32963 31815 32969
rect 31757 32929 31769 32963
rect 31803 32960 31815 32963
rect 33336 32960 33364 32988
rect 31803 32932 33364 32960
rect 31803 32929 31815 32932
rect 31757 32923 31815 32929
rect 34238 32920 34244 32972
rect 34296 32920 34302 32972
rect 2590 32852 2596 32904
rect 2648 32852 2654 32904
rect 2961 32895 3019 32901
rect 2961 32861 2973 32895
rect 3007 32892 3019 32895
rect 3786 32892 3792 32904
rect 3007 32864 3792 32892
rect 3007 32861 3019 32864
rect 2961 32855 3019 32861
rect 3786 32852 3792 32864
rect 3844 32852 3850 32904
rect 5077 32895 5135 32901
rect 5077 32861 5089 32895
rect 5123 32892 5135 32895
rect 6270 32892 6276 32904
rect 5123 32864 6276 32892
rect 5123 32861 5135 32864
rect 5077 32855 5135 32861
rect 6270 32852 6276 32864
rect 6328 32852 6334 32904
rect 30469 32895 30527 32901
rect 30469 32861 30481 32895
rect 30515 32861 30527 32895
rect 30469 32855 30527 32861
rect 31849 32895 31907 32901
rect 31849 32861 31861 32895
rect 31895 32892 31907 32895
rect 32030 32892 32036 32904
rect 31895 32864 32036 32892
rect 31895 32861 31907 32864
rect 31849 32855 31907 32861
rect 4522 32784 4528 32836
rect 4580 32784 4586 32836
rect 3510 32716 3516 32768
rect 3568 32716 3574 32768
rect 30282 32716 30288 32768
rect 30340 32716 30346 32768
rect 30484 32756 30512 32855
rect 32030 32852 32036 32864
rect 32088 32852 32094 32904
rect 32306 32852 32312 32904
rect 32364 32892 32370 32904
rect 32585 32895 32643 32901
rect 32585 32892 32597 32895
rect 32364 32864 32597 32892
rect 32364 32852 32370 32864
rect 32585 32861 32597 32864
rect 32631 32861 32643 32895
rect 32585 32855 32643 32861
rect 33321 32895 33379 32901
rect 33321 32861 33333 32895
rect 33367 32892 33379 32895
rect 33594 32892 33600 32904
rect 33367 32864 33600 32892
rect 33367 32861 33379 32864
rect 33321 32855 33379 32861
rect 33594 32852 33600 32864
rect 33652 32852 33658 32904
rect 35866 32892 35894 33068
rect 36078 33056 36084 33068
rect 36136 33096 36142 33108
rect 36354 33096 36360 33108
rect 36136 33068 36360 33096
rect 36136 33056 36142 33068
rect 36354 33056 36360 33068
rect 36412 33056 36418 33108
rect 34808 32864 35894 32892
rect 35989 32895 36047 32901
rect 31021 32827 31079 32833
rect 31021 32793 31033 32827
rect 31067 32824 31079 32827
rect 31938 32824 31944 32836
rect 31067 32796 31944 32824
rect 31067 32793 31079 32796
rect 31021 32787 31079 32793
rect 31938 32784 31944 32796
rect 31996 32784 32002 32836
rect 34238 32784 34244 32836
rect 34296 32824 34302 32836
rect 34808 32833 34836 32864
rect 35989 32861 36001 32895
rect 36035 32892 36047 32895
rect 36170 32892 36176 32904
rect 36035 32864 36176 32892
rect 36035 32861 36047 32864
rect 35989 32855 36047 32861
rect 36170 32852 36176 32864
rect 36228 32852 36234 32904
rect 36262 32852 36268 32904
rect 36320 32852 36326 32904
rect 34793 32827 34851 32833
rect 34793 32824 34805 32827
rect 34296 32796 34805 32824
rect 34296 32784 34302 32796
rect 34793 32793 34805 32796
rect 34839 32793 34851 32827
rect 35526 32824 35532 32836
rect 34793 32787 34851 32793
rect 35268 32796 35532 32824
rect 34514 32756 34520 32768
rect 30484 32728 34520 32756
rect 34514 32716 34520 32728
rect 34572 32716 34578 32768
rect 35268 32765 35296 32796
rect 35526 32784 35532 32796
rect 35584 32784 35590 32836
rect 37182 32784 37188 32836
rect 37240 32784 37246 32836
rect 35253 32759 35311 32765
rect 35253 32725 35265 32759
rect 35299 32725 35311 32759
rect 35253 32719 35311 32725
rect 35345 32759 35403 32765
rect 35345 32725 35357 32759
rect 35391 32756 35403 32759
rect 35434 32756 35440 32768
rect 35391 32728 35440 32756
rect 35391 32725 35403 32728
rect 35345 32719 35403 32725
rect 35434 32716 35440 32728
rect 35492 32716 35498 32768
rect 1104 32666 37812 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 37812 32666
rect 1104 32592 37812 32614
rect 4522 32512 4528 32564
rect 4580 32512 4586 32564
rect 4985 32555 5043 32561
rect 4985 32521 4997 32555
rect 5031 32552 5043 32555
rect 5994 32552 6000 32564
rect 5031 32524 6000 32552
rect 5031 32521 5043 32524
rect 4985 32515 5043 32521
rect 5994 32512 6000 32524
rect 6052 32512 6058 32564
rect 31941 32555 31999 32561
rect 31941 32521 31953 32555
rect 31987 32552 31999 32555
rect 33226 32552 33232 32564
rect 31987 32524 33232 32552
rect 31987 32521 31999 32524
rect 31941 32515 31999 32521
rect 33226 32512 33232 32524
rect 33284 32512 33290 32564
rect 36538 32552 36544 32564
rect 35866 32524 36544 32552
rect 3050 32444 3056 32496
rect 3108 32444 3114 32496
rect 2590 32376 2596 32428
rect 2648 32376 2654 32428
rect 4249 32419 4307 32425
rect 4249 32385 4261 32419
rect 4295 32416 4307 32419
rect 4540 32416 4568 32512
rect 32677 32487 32735 32493
rect 32677 32453 32689 32487
rect 32723 32484 32735 32487
rect 34238 32484 34244 32496
rect 32723 32456 34244 32484
rect 32723 32453 32735 32456
rect 32677 32447 32735 32453
rect 34238 32444 34244 32456
rect 34296 32444 34302 32496
rect 35866 32484 35894 32524
rect 36538 32512 36544 32524
rect 36596 32512 36602 32564
rect 35636 32456 35894 32484
rect 4295 32388 4568 32416
rect 4295 32385 4307 32388
rect 4249 32379 4307 32385
rect 4614 32376 4620 32428
rect 4672 32376 4678 32428
rect 34149 32419 34207 32425
rect 34149 32385 34161 32419
rect 34195 32416 34207 32419
rect 34330 32416 34336 32428
rect 34195 32388 34336 32416
rect 34195 32385 34207 32388
rect 34149 32379 34207 32385
rect 34330 32376 34336 32388
rect 34388 32376 34394 32428
rect 35636 32425 35664 32456
rect 36078 32444 36084 32496
rect 36136 32484 36142 32496
rect 36173 32487 36231 32493
rect 36173 32484 36185 32487
rect 36136 32456 36185 32484
rect 36136 32444 36142 32456
rect 36173 32453 36185 32456
rect 36219 32453 36231 32487
rect 36173 32447 36231 32453
rect 36354 32444 36360 32496
rect 36412 32484 36418 32496
rect 36725 32487 36783 32493
rect 36725 32484 36737 32487
rect 36412 32456 36737 32484
rect 36412 32444 36418 32456
rect 36725 32453 36737 32456
rect 36771 32484 36783 32487
rect 36814 32484 36820 32496
rect 36771 32456 36820 32484
rect 36771 32453 36783 32456
rect 36725 32447 36783 32453
rect 36814 32444 36820 32456
rect 36872 32444 36878 32496
rect 35621 32419 35679 32425
rect 35621 32385 35633 32419
rect 35667 32385 35679 32419
rect 35621 32379 35679 32385
rect 35802 32376 35808 32428
rect 35860 32376 35866 32428
rect 1578 32308 1584 32360
rect 1636 32308 1642 32360
rect 4433 32351 4491 32357
rect 4433 32317 4445 32351
rect 4479 32348 4491 32351
rect 4632 32348 4660 32376
rect 4479 32320 4660 32348
rect 4479 32317 4491 32320
rect 4433 32311 4491 32317
rect 30650 32308 30656 32360
rect 30708 32308 30714 32360
rect 31205 32351 31263 32357
rect 31205 32317 31217 32351
rect 31251 32348 31263 32351
rect 31389 32351 31447 32357
rect 31389 32348 31401 32351
rect 31251 32320 31401 32348
rect 31251 32317 31263 32320
rect 31205 32311 31263 32317
rect 31389 32317 31401 32320
rect 31435 32348 31447 32351
rect 31435 32320 32628 32348
rect 31435 32317 31447 32320
rect 31389 32311 31447 32317
rect 30282 32240 30288 32292
rect 30340 32280 30346 32292
rect 32309 32283 32367 32289
rect 32309 32280 32321 32283
rect 30340 32252 32321 32280
rect 30340 32240 30346 32252
rect 32309 32249 32321 32252
rect 32355 32249 32367 32283
rect 32600 32280 32628 32320
rect 33686 32308 33692 32360
rect 33744 32308 33750 32360
rect 35161 32351 35219 32357
rect 35161 32317 35173 32351
rect 35207 32348 35219 32351
rect 35710 32348 35716 32360
rect 35207 32320 35716 32348
rect 35207 32317 35219 32320
rect 35161 32311 35219 32317
rect 35710 32308 35716 32320
rect 35768 32308 35774 32360
rect 36630 32280 36636 32292
rect 32600 32252 36636 32280
rect 32309 32243 32367 32249
rect 36630 32240 36636 32252
rect 36688 32240 36694 32292
rect 32217 32215 32275 32221
rect 32217 32181 32229 32215
rect 32263 32212 32275 32215
rect 33962 32212 33968 32224
rect 32263 32184 33968 32212
rect 32263 32181 32275 32184
rect 32217 32175 32275 32181
rect 33962 32172 33968 32184
rect 34020 32172 34026 32224
rect 1104 32122 37812 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 37812 32122
rect 1104 32048 37812 32070
rect 2590 31968 2596 32020
rect 2648 31968 2654 32020
rect 30282 31968 30288 32020
rect 30340 31968 30346 32020
rect 30650 31968 30656 32020
rect 30708 32008 30714 32020
rect 31481 32011 31539 32017
rect 31481 32008 31493 32011
rect 30708 31980 31493 32008
rect 30708 31968 30714 31980
rect 31481 31977 31493 31980
rect 31527 31977 31539 32011
rect 31481 31971 31539 31977
rect 32582 31968 32588 32020
rect 32640 31968 32646 32020
rect 33318 31968 33324 32020
rect 33376 31968 33382 32020
rect 34790 32008 34796 32020
rect 33796 31980 34796 32008
rect 2409 31875 2467 31881
rect 2409 31841 2421 31875
rect 2455 31872 2467 31875
rect 2608 31872 2636 31968
rect 2455 31844 2636 31872
rect 30300 31872 30328 31968
rect 31389 31943 31447 31949
rect 31389 31909 31401 31943
rect 31435 31940 31447 31943
rect 32600 31940 32628 31968
rect 31435 31912 32628 31940
rect 31435 31909 31447 31912
rect 31389 31903 31447 31909
rect 30745 31875 30803 31881
rect 30745 31872 30757 31875
rect 30300 31844 30757 31872
rect 2455 31841 2467 31844
rect 2409 31835 2467 31841
rect 30745 31841 30757 31844
rect 30791 31841 30803 31875
rect 30745 31835 30803 31841
rect 32122 31832 32128 31884
rect 32180 31832 32186 31884
rect 33229 31875 33287 31881
rect 33229 31841 33241 31875
rect 33275 31872 33287 31875
rect 33336 31872 33364 31968
rect 33275 31844 33364 31872
rect 33275 31841 33287 31844
rect 33229 31835 33287 31841
rect 2685 31807 2743 31813
rect 2685 31773 2697 31807
rect 2731 31804 2743 31807
rect 2774 31804 2780 31816
rect 2731 31776 2780 31804
rect 2731 31773 2743 31776
rect 2685 31767 2743 31773
rect 2774 31764 2780 31776
rect 2832 31764 2838 31816
rect 2958 31764 2964 31816
rect 3016 31764 3022 31816
rect 3513 31807 3571 31813
rect 3513 31773 3525 31807
rect 3559 31804 3571 31807
rect 3789 31807 3847 31813
rect 3789 31804 3801 31807
rect 3559 31776 3801 31804
rect 3559 31773 3571 31776
rect 3513 31767 3571 31773
rect 3789 31773 3801 31776
rect 3835 31773 3847 31807
rect 3789 31767 3847 31773
rect 8110 31764 8116 31816
rect 8168 31764 8174 31816
rect 8757 31807 8815 31813
rect 8757 31773 8769 31807
rect 8803 31804 8815 31807
rect 10870 31804 10876 31816
rect 8803 31776 10876 31804
rect 8803 31773 8815 31776
rect 8757 31767 8815 31773
rect 10870 31764 10876 31776
rect 10928 31764 10934 31816
rect 32309 31807 32367 31813
rect 32309 31773 32321 31807
rect 32355 31804 32367 31807
rect 32766 31804 32772 31816
rect 32355 31776 32772 31804
rect 32355 31773 32367 31776
rect 32309 31767 32367 31773
rect 32766 31764 32772 31776
rect 32824 31764 32830 31816
rect 32861 31807 32919 31813
rect 32861 31773 32873 31807
rect 32907 31804 32919 31807
rect 33796 31804 33824 31980
rect 34790 31968 34796 31980
rect 34848 31968 34854 32020
rect 35434 31968 35440 32020
rect 35492 31968 35498 32020
rect 36170 31968 36176 32020
rect 36228 32008 36234 32020
rect 36817 32011 36875 32017
rect 36817 32008 36829 32011
rect 36228 31980 36829 32008
rect 36228 31968 36234 31980
rect 36817 31977 36829 31980
rect 36863 31977 36875 32011
rect 36817 31971 36875 31977
rect 35452 31940 35480 31968
rect 33980 31912 35480 31940
rect 33980 31881 34008 31912
rect 36722 31900 36728 31952
rect 36780 31940 36786 31952
rect 36909 31943 36967 31949
rect 36909 31940 36921 31943
rect 36780 31912 36921 31940
rect 36780 31900 36786 31912
rect 36909 31909 36921 31912
rect 36955 31909 36967 31943
rect 36909 31903 36967 31909
rect 36998 31900 37004 31952
rect 37056 31900 37062 31952
rect 33965 31875 34023 31881
rect 33965 31841 33977 31875
rect 34011 31841 34023 31875
rect 34606 31872 34612 31884
rect 33965 31835 34023 31841
rect 34440 31844 34612 31872
rect 34440 31804 34468 31844
rect 34606 31832 34612 31844
rect 34664 31832 34670 31884
rect 35342 31832 35348 31884
rect 35400 31872 35406 31884
rect 35437 31875 35495 31881
rect 35437 31872 35449 31875
rect 35400 31844 35449 31872
rect 35400 31832 35406 31844
rect 35437 31841 35449 31844
rect 35483 31841 35495 31875
rect 35437 31835 35495 31841
rect 36814 31832 36820 31884
rect 36872 31872 36878 31884
rect 37369 31875 37427 31881
rect 37369 31872 37381 31875
rect 36872 31844 37381 31872
rect 36872 31832 36878 31844
rect 37369 31841 37381 31844
rect 37415 31841 37427 31875
rect 37369 31835 37427 31841
rect 32907 31776 33824 31804
rect 33888 31776 34468 31804
rect 34517 31807 34575 31813
rect 32907 31773 32919 31776
rect 32861 31767 32919 31773
rect 33781 31739 33839 31745
rect 33781 31705 33793 31739
rect 33827 31736 33839 31739
rect 33888 31736 33916 31776
rect 34517 31773 34529 31807
rect 34563 31804 34575 31807
rect 34790 31804 34796 31816
rect 34563 31776 34796 31804
rect 34563 31773 34575 31776
rect 34517 31767 34575 31773
rect 34790 31764 34796 31776
rect 34848 31764 34854 31816
rect 35526 31764 35532 31816
rect 35584 31804 35590 31816
rect 35693 31807 35751 31813
rect 35693 31804 35705 31807
rect 35584 31776 35705 31804
rect 35584 31764 35590 31776
rect 35693 31773 35705 31776
rect 35739 31773 35751 31807
rect 35693 31767 35751 31773
rect 33827 31708 33916 31736
rect 33827 31705 33839 31708
rect 33781 31699 33839 31705
rect 4430 31628 4436 31680
rect 4488 31628 4494 31680
rect 34238 31628 34244 31680
rect 34296 31668 34302 31680
rect 34606 31668 34612 31680
rect 34296 31640 34612 31668
rect 34296 31628 34302 31640
rect 34606 31628 34612 31640
rect 34664 31628 34670 31680
rect 35345 31671 35403 31677
rect 35345 31637 35357 31671
rect 35391 31668 35403 31671
rect 35526 31668 35532 31680
rect 35391 31640 35532 31668
rect 35391 31637 35403 31640
rect 35345 31631 35403 31637
rect 35526 31628 35532 31640
rect 35584 31628 35590 31680
rect 1104 31578 37812 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 37812 31578
rect 1104 31504 37812 31526
rect 2774 31424 2780 31476
rect 2832 31464 2838 31476
rect 3605 31467 3663 31473
rect 3605 31464 3617 31467
rect 2832 31436 3617 31464
rect 2832 31424 2838 31436
rect 3605 31433 3617 31436
rect 3651 31433 3663 31467
rect 3605 31427 3663 31433
rect 34149 31467 34207 31473
rect 34149 31433 34161 31467
rect 34195 31464 34207 31467
rect 35802 31464 35808 31476
rect 34195 31436 35808 31464
rect 34195 31433 34207 31436
rect 34149 31427 34207 31433
rect 35802 31424 35808 31436
rect 35860 31424 35866 31476
rect 36814 31424 36820 31476
rect 36872 31424 36878 31476
rect 33520 31368 35894 31396
rect 2590 31288 2596 31340
rect 2648 31288 2654 31340
rect 4249 31331 4307 31337
rect 4249 31297 4261 31331
rect 4295 31328 4307 31331
rect 4430 31328 4436 31340
rect 4295 31300 4436 31328
rect 4295 31297 4307 31300
rect 4249 31291 4307 31297
rect 4430 31288 4436 31300
rect 4488 31328 4494 31340
rect 4614 31328 4620 31340
rect 4488 31300 4620 31328
rect 4488 31288 4494 31300
rect 4614 31288 4620 31300
rect 4672 31288 4678 31340
rect 31938 31288 31944 31340
rect 31996 31328 32002 31340
rect 32769 31331 32827 31337
rect 32769 31328 32781 31331
rect 31996 31300 32781 31328
rect 31996 31288 32002 31300
rect 32769 31297 32781 31300
rect 32815 31297 32827 31331
rect 32769 31291 32827 31297
rect 33520 31272 33548 31368
rect 35434 31288 35440 31340
rect 35492 31288 35498 31340
rect 35526 31288 35532 31340
rect 35584 31328 35590 31340
rect 35759 31331 35817 31337
rect 35759 31328 35771 31331
rect 35584 31300 35771 31328
rect 35584 31288 35590 31300
rect 35759 31297 35771 31300
rect 35805 31297 35817 31331
rect 35759 31291 35817 31297
rect 1578 31220 1584 31272
rect 1636 31220 1642 31272
rect 2866 31220 2872 31272
rect 2924 31220 2930 31272
rect 33502 31220 33508 31272
rect 33560 31220 33566 31272
rect 35161 31263 35219 31269
rect 35161 31229 35173 31263
rect 35207 31229 35219 31263
rect 35866 31260 35894 31368
rect 36262 31356 36268 31408
rect 36320 31356 36326 31408
rect 36998 31260 37004 31272
rect 35866 31232 37004 31260
rect 35161 31223 35219 31229
rect 33410 31152 33416 31204
rect 33468 31192 33474 31204
rect 35176 31192 35204 31223
rect 36998 31220 37004 31232
rect 37056 31220 37062 31272
rect 37826 31192 37832 31204
rect 33468 31164 34284 31192
rect 35176 31164 37832 31192
rect 33468 31152 33474 31164
rect 3513 31127 3571 31133
rect 3513 31093 3525 31127
rect 3559 31124 3571 31127
rect 4062 31124 4068 31136
rect 3559 31096 4068 31124
rect 3559 31093 3571 31096
rect 3513 31087 3571 31093
rect 4062 31084 4068 31096
rect 4120 31084 4126 31136
rect 34256 31124 34284 31164
rect 37826 31152 37832 31164
rect 37884 31152 37890 31204
rect 36446 31124 36452 31136
rect 34256 31096 36452 31124
rect 36446 31084 36452 31096
rect 36504 31084 36510 31136
rect 1104 31034 37812 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 37812 31034
rect 1104 30960 37812 30982
rect 2590 30920 2596 30932
rect 2424 30892 2596 30920
rect 2424 30793 2452 30892
rect 2590 30880 2596 30892
rect 2648 30880 2654 30932
rect 2866 30880 2872 30932
rect 2924 30880 2930 30932
rect 3234 30880 3240 30932
rect 3292 30920 3298 30932
rect 3789 30923 3847 30929
rect 3789 30920 3801 30923
rect 3292 30892 3801 30920
rect 3292 30880 3298 30892
rect 3789 30889 3801 30892
rect 3835 30889 3847 30923
rect 3789 30883 3847 30889
rect 33410 30880 33416 30932
rect 33468 30880 33474 30932
rect 33781 30923 33839 30929
rect 33781 30889 33793 30923
rect 33827 30920 33839 30923
rect 34054 30920 34060 30932
rect 33827 30892 34060 30920
rect 33827 30889 33839 30892
rect 33781 30883 33839 30889
rect 34054 30880 34060 30892
rect 34112 30880 34118 30932
rect 4614 30812 4620 30864
rect 4672 30812 4678 30864
rect 2409 30787 2467 30793
rect 2409 30753 2421 30787
rect 2455 30753 2467 30787
rect 2409 30747 2467 30753
rect 4890 30744 4896 30796
rect 4948 30784 4954 30796
rect 4985 30787 5043 30793
rect 4985 30784 4997 30787
rect 4948 30756 4997 30784
rect 4948 30744 4954 30756
rect 4985 30753 4997 30756
rect 5031 30753 5043 30787
rect 4985 30747 5043 30753
rect 32398 30744 32404 30796
rect 32456 30744 32462 30796
rect 33229 30787 33287 30793
rect 33229 30753 33241 30787
rect 33275 30784 33287 30787
rect 33428 30784 33456 30880
rect 34790 30812 34796 30864
rect 34848 30852 34854 30864
rect 35069 30855 35127 30861
rect 35069 30852 35081 30855
rect 34848 30824 35081 30852
rect 34848 30812 34854 30824
rect 35069 30821 35081 30824
rect 35115 30821 35127 30855
rect 35069 30815 35127 30821
rect 33275 30756 33456 30784
rect 34517 30787 34575 30793
rect 33275 30753 33287 30756
rect 33229 30747 33287 30753
rect 34517 30753 34529 30787
rect 34563 30784 34575 30787
rect 34698 30784 34704 30796
rect 34563 30756 34704 30784
rect 34563 30753 34575 30756
rect 34517 30747 34575 30753
rect 34698 30744 34704 30756
rect 34756 30744 34762 30796
rect 2685 30719 2743 30725
rect 2685 30685 2697 30719
rect 2731 30716 2743 30719
rect 3050 30716 3056 30728
rect 2731 30688 3056 30716
rect 2731 30685 2743 30688
rect 2685 30679 2743 30685
rect 3050 30676 3056 30688
rect 3108 30676 3114 30728
rect 3418 30676 3424 30728
rect 3476 30676 3482 30728
rect 4433 30719 4491 30725
rect 4433 30685 4445 30719
rect 4479 30716 4491 30719
rect 4706 30716 4712 30728
rect 4479 30688 4712 30716
rect 4479 30685 4491 30688
rect 4433 30679 4491 30685
rect 4706 30676 4712 30688
rect 4764 30676 4770 30728
rect 32416 30716 32444 30744
rect 33873 30719 33931 30725
rect 33873 30716 33885 30719
rect 32416 30688 33885 30716
rect 33873 30685 33885 30688
rect 33919 30685 33931 30719
rect 33873 30679 33931 30685
rect 35250 30676 35256 30728
rect 35308 30716 35314 30728
rect 35345 30719 35403 30725
rect 35345 30716 35357 30719
rect 35308 30688 35357 30716
rect 35308 30676 35314 30688
rect 35345 30685 35357 30688
rect 35391 30685 35403 30719
rect 35345 30679 35403 30685
rect 35986 30676 35992 30728
rect 36044 30676 36050 30728
rect 36262 30676 36268 30728
rect 36320 30676 36326 30728
rect 34790 30608 34796 30660
rect 34848 30608 34854 30660
rect 37182 30608 37188 30660
rect 37240 30608 37246 30660
rect 4525 30583 4583 30589
rect 4525 30549 4537 30583
rect 4571 30580 4583 30583
rect 4614 30580 4620 30592
rect 4571 30552 4620 30580
rect 4571 30549 4583 30552
rect 4525 30543 4583 30549
rect 4614 30540 4620 30552
rect 4672 30540 4678 30592
rect 35253 30583 35311 30589
rect 35253 30549 35265 30583
rect 35299 30580 35311 30583
rect 35526 30580 35532 30592
rect 35299 30552 35532 30580
rect 35299 30549 35311 30552
rect 35253 30543 35311 30549
rect 35526 30540 35532 30552
rect 35584 30540 35590 30592
rect 1104 30490 37812 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 37812 30490
rect 1104 30416 37812 30438
rect 3050 30336 3056 30388
rect 3108 30376 3114 30388
rect 3108 30348 3464 30376
rect 3108 30336 3114 30348
rect 3436 30317 3464 30348
rect 35986 30336 35992 30388
rect 36044 30376 36050 30388
rect 36817 30379 36875 30385
rect 36817 30376 36829 30379
rect 36044 30348 36829 30376
rect 36044 30336 36050 30348
rect 36817 30345 36829 30348
rect 36863 30345 36875 30379
rect 36817 30339 36875 30345
rect 3421 30311 3479 30317
rect 2700 30280 3372 30308
rect 2700 30252 2728 30280
rect 2682 30200 2688 30252
rect 2740 30200 2746 30252
rect 3073 30243 3131 30249
rect 3073 30209 3085 30243
rect 3119 30240 3131 30243
rect 3234 30240 3240 30252
rect 3119 30212 3240 30240
rect 3119 30209 3131 30212
rect 3073 30203 3131 30209
rect 3234 30200 3240 30212
rect 3292 30200 3298 30252
rect 3344 30249 3372 30280
rect 3421 30277 3433 30311
rect 3467 30277 3479 30311
rect 3421 30271 3479 30277
rect 34514 30268 34520 30320
rect 34572 30308 34578 30320
rect 34609 30311 34667 30317
rect 34609 30308 34621 30311
rect 34572 30280 34621 30308
rect 34572 30268 34578 30280
rect 34609 30277 34621 30280
rect 34655 30277 34667 30311
rect 34609 30271 34667 30277
rect 35526 30268 35532 30320
rect 35584 30308 35590 30320
rect 35682 30311 35740 30317
rect 35682 30308 35694 30311
rect 35584 30280 35694 30308
rect 35584 30268 35590 30280
rect 35682 30277 35694 30280
rect 35728 30277 35740 30311
rect 35682 30271 35740 30277
rect 3329 30243 3387 30249
rect 3329 30209 3341 30243
rect 3375 30209 3387 30243
rect 3329 30203 3387 30209
rect 33134 30200 33140 30252
rect 33192 30240 33198 30252
rect 33965 30243 34023 30249
rect 33965 30240 33977 30243
rect 33192 30212 33977 30240
rect 33192 30200 33198 30212
rect 33965 30209 33977 30212
rect 34011 30209 34023 30243
rect 33965 30203 34023 30209
rect 35250 30200 35256 30252
rect 35308 30200 35314 30252
rect 35342 30200 35348 30252
rect 35400 30240 35406 30252
rect 35437 30243 35495 30249
rect 35437 30240 35449 30243
rect 35400 30212 35449 30240
rect 35400 30200 35406 30212
rect 35437 30209 35449 30212
rect 35483 30209 35495 30243
rect 35437 30203 35495 30209
rect 4062 30132 4068 30184
rect 4120 30132 4126 30184
rect 1949 30039 2007 30045
rect 1949 30005 1961 30039
rect 1995 30036 2007 30039
rect 2958 30036 2964 30048
rect 1995 30008 2964 30036
rect 1995 30005 2007 30008
rect 1949 29999 2007 30005
rect 2958 29996 2964 30008
rect 3016 29996 3022 30048
rect 34698 29996 34704 30048
rect 34756 29996 34762 30048
rect 1104 29946 37812 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 37812 29946
rect 1104 29872 37812 29894
rect 1949 29835 2007 29841
rect 1949 29801 1961 29835
rect 1995 29832 2007 29835
rect 3418 29832 3424 29844
rect 1995 29804 3424 29832
rect 1995 29801 2007 29804
rect 1949 29795 2007 29801
rect 3418 29792 3424 29804
rect 3476 29792 3482 29844
rect 3786 29792 3792 29844
rect 3844 29792 3850 29844
rect 6270 29792 6276 29844
rect 6328 29792 6334 29844
rect 10870 29792 10876 29844
rect 10928 29792 10934 29844
rect 34698 29792 34704 29844
rect 34756 29792 34762 29844
rect 34790 29792 34796 29844
rect 34848 29832 34854 29844
rect 35069 29835 35127 29841
rect 35069 29832 35081 29835
rect 34848 29804 35081 29832
rect 34848 29792 34854 29804
rect 35069 29801 35081 29804
rect 35115 29832 35127 29835
rect 35710 29832 35716 29844
rect 35115 29804 35716 29832
rect 35115 29801 35127 29804
rect 35069 29795 35127 29801
rect 35710 29792 35716 29804
rect 35768 29832 35774 29844
rect 37369 29835 37427 29841
rect 37369 29832 37381 29835
rect 35768 29804 37381 29832
rect 35768 29792 35774 29804
rect 37369 29801 37381 29804
rect 37415 29801 37427 29835
rect 37369 29795 37427 29801
rect 6914 29656 6920 29708
rect 6972 29696 6978 29708
rect 8110 29696 8116 29708
rect 6972 29668 8116 29696
rect 6972 29656 6978 29668
rect 8110 29656 8116 29668
rect 8168 29656 8174 29708
rect 34716 29696 34744 29792
rect 35345 29699 35403 29705
rect 35345 29696 35357 29699
rect 34716 29668 35357 29696
rect 35345 29665 35357 29668
rect 35391 29665 35403 29699
rect 35345 29659 35403 29665
rect 36262 29656 36268 29708
rect 36320 29696 36326 29708
rect 36449 29699 36507 29705
rect 36449 29696 36461 29699
rect 36320 29668 36461 29696
rect 36320 29656 36326 29668
rect 36449 29665 36461 29668
rect 36495 29665 36507 29699
rect 36449 29659 36507 29665
rect 2682 29588 2688 29640
rect 2740 29628 2746 29640
rect 3329 29631 3387 29637
rect 3329 29628 3341 29631
rect 2740 29600 3341 29628
rect 2740 29588 2746 29600
rect 3329 29597 3341 29600
rect 3375 29597 3387 29631
rect 3329 29591 3387 29597
rect 3786 29588 3792 29640
rect 3844 29628 3850 29640
rect 4341 29631 4399 29637
rect 4341 29628 4353 29631
rect 3844 29600 4353 29628
rect 3844 29588 3850 29600
rect 4341 29597 4353 29600
rect 4387 29597 4399 29631
rect 4341 29591 4399 29597
rect 4614 29588 4620 29640
rect 4672 29588 4678 29640
rect 11517 29631 11575 29637
rect 11517 29597 11529 29631
rect 11563 29628 11575 29631
rect 13446 29628 13452 29640
rect 11563 29600 13452 29628
rect 11563 29597 11575 29600
rect 11517 29591 11575 29597
rect 13446 29588 13452 29600
rect 13504 29588 13510 29640
rect 35989 29631 36047 29637
rect 35989 29597 36001 29631
rect 36035 29628 36047 29631
rect 36173 29631 36231 29637
rect 36173 29628 36185 29631
rect 36035 29600 36185 29628
rect 36035 29597 36047 29600
rect 35989 29591 36047 29597
rect 36173 29597 36185 29600
rect 36219 29597 36231 29631
rect 36173 29591 36231 29597
rect 3084 29563 3142 29569
rect 3084 29529 3096 29563
rect 3130 29560 3142 29563
rect 4632 29560 4660 29588
rect 3130 29532 4660 29560
rect 3130 29529 3142 29532
rect 3084 29523 3142 29529
rect 1104 29402 37812 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 37812 29402
rect 1104 29328 37812 29350
rect 3234 29248 3240 29300
rect 3292 29288 3298 29300
rect 4341 29291 4399 29297
rect 4341 29288 4353 29291
rect 3292 29260 4353 29288
rect 3292 29248 3298 29260
rect 4341 29257 4353 29260
rect 4387 29257 4399 29291
rect 4341 29251 4399 29257
rect 32766 29248 32772 29300
rect 32824 29248 32830 29300
rect 34698 29248 34704 29300
rect 34756 29248 34762 29300
rect 4801 29223 4859 29229
rect 4801 29189 4813 29223
rect 4847 29220 4859 29223
rect 4890 29220 4896 29232
rect 4847 29192 4896 29220
rect 4847 29189 4859 29192
rect 4801 29183 4859 29189
rect 4890 29180 4896 29192
rect 4948 29220 4954 29232
rect 5353 29223 5411 29229
rect 5353 29220 5365 29223
rect 4948 29192 5365 29220
rect 4948 29180 4954 29192
rect 5353 29189 5365 29192
rect 5399 29189 5411 29223
rect 5353 29183 5411 29189
rect 2685 29155 2743 29161
rect 2685 29121 2697 29155
rect 2731 29152 2743 29155
rect 2774 29152 2780 29164
rect 2731 29124 2780 29152
rect 2731 29121 2743 29124
rect 2685 29115 2743 29121
rect 2774 29112 2780 29124
rect 2832 29112 2838 29164
rect 4062 29112 4068 29164
rect 4120 29152 4126 29164
rect 30374 29152 30380 29164
rect 4120 29124 5028 29152
rect 4120 29112 4126 29124
rect 1578 29044 1584 29096
rect 1636 29044 1642 29096
rect 2961 29087 3019 29093
rect 2961 29053 2973 29087
rect 3007 29084 3019 29087
rect 3605 29087 3663 29093
rect 3605 29084 3617 29087
rect 3007 29056 3617 29084
rect 3007 29053 3019 29056
rect 2961 29047 3019 29053
rect 3605 29053 3617 29056
rect 3651 29053 3663 29087
rect 3605 29047 3663 29053
rect 4154 29044 4160 29096
rect 4212 29044 4218 29096
rect 4525 29019 4583 29025
rect 4525 28985 4537 29019
rect 4571 29016 4583 29019
rect 4614 29016 4620 29028
rect 4571 28988 4620 29016
rect 4571 28985 4583 28988
rect 4525 28979 4583 28985
rect 4614 28976 4620 28988
rect 4672 28976 4678 29028
rect 5000 29025 5028 29124
rect 28460 29124 30380 29152
rect 20438 29044 20444 29096
rect 20496 29044 20502 29096
rect 28460 29028 28488 29124
rect 30374 29112 30380 29124
rect 30432 29112 30438 29164
rect 34425 29155 34483 29161
rect 34425 29121 34437 29155
rect 34471 29152 34483 29155
rect 34606 29152 34612 29164
rect 34471 29124 34612 29152
rect 34471 29121 34483 29124
rect 34425 29115 34483 29121
rect 34606 29112 34612 29124
rect 34664 29112 34670 29164
rect 32122 29044 32128 29096
rect 32180 29044 32186 29096
rect 4985 29019 5043 29025
rect 4985 28985 4997 29019
rect 5031 28985 5043 29019
rect 19889 29019 19947 29025
rect 19889 29016 19901 29019
rect 4985 28979 5043 28985
rect 19260 28988 19901 29016
rect 19260 28960 19288 28988
rect 19889 28985 19901 28988
rect 19935 28985 19947 29019
rect 19889 28979 19947 28985
rect 28442 28976 28448 29028
rect 28500 28976 28506 29028
rect 29089 29019 29147 29025
rect 29089 28985 29101 29019
rect 29135 29016 29147 29019
rect 29914 29016 29920 29028
rect 29135 28988 29920 29016
rect 29135 28985 29147 28988
rect 29089 28979 29147 28985
rect 29914 28976 29920 28988
rect 29972 28976 29978 29028
rect 34716 29025 34744 29248
rect 35805 29155 35863 29161
rect 35805 29121 35817 29155
rect 35851 29152 35863 29155
rect 36078 29152 36084 29164
rect 35851 29124 36084 29152
rect 35851 29121 35863 29124
rect 35805 29115 35863 29121
rect 36078 29112 36084 29124
rect 36136 29112 36142 29164
rect 35621 29087 35679 29093
rect 35621 29053 35633 29087
rect 35667 29084 35679 29087
rect 35667 29056 35894 29084
rect 35667 29053 35679 29056
rect 35621 29047 35679 29053
rect 34701 29019 34759 29025
rect 34701 28985 34713 29019
rect 34747 28985 34759 29019
rect 34701 28979 34759 28985
rect 34790 28976 34796 29028
rect 34848 29016 34854 29028
rect 34977 29019 35035 29025
rect 34977 29016 34989 29019
rect 34848 28988 34989 29016
rect 34848 28976 34854 28988
rect 34977 28985 34989 28988
rect 35023 28985 35035 29019
rect 35866 29016 35894 29056
rect 36906 29044 36912 29096
rect 36964 29044 36970 29096
rect 36814 29016 36820 29028
rect 35866 28988 36820 29016
rect 34977 28979 35035 28985
rect 36814 28976 36820 28988
rect 36872 28976 36878 29028
rect 3513 28951 3571 28957
rect 3513 28917 3525 28951
rect 3559 28948 3571 28951
rect 3878 28948 3884 28960
rect 3559 28920 3884 28948
rect 3559 28917 3571 28920
rect 3513 28911 3571 28917
rect 3878 28908 3884 28920
rect 3936 28908 3942 28960
rect 4890 28908 4896 28960
rect 4948 28908 4954 28960
rect 19242 28908 19248 28960
rect 19300 28908 19306 28960
rect 34885 28951 34943 28957
rect 34885 28917 34897 28951
rect 34931 28948 34943 28951
rect 35526 28948 35532 28960
rect 34931 28920 35532 28948
rect 34931 28917 34943 28920
rect 34885 28911 34943 28917
rect 35526 28908 35532 28920
rect 35584 28908 35590 28960
rect 1104 28858 37812 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 37812 28858
rect 1104 28784 37812 28806
rect 3329 28747 3387 28753
rect 3329 28713 3341 28747
rect 3375 28744 3387 28747
rect 4062 28744 4068 28756
rect 3375 28716 4068 28744
rect 3375 28713 3387 28716
rect 3329 28707 3387 28713
rect 4062 28704 4068 28716
rect 4120 28704 4126 28756
rect 19889 28747 19947 28753
rect 19889 28713 19901 28747
rect 19935 28744 19947 28747
rect 20346 28744 20352 28756
rect 19935 28716 20352 28744
rect 19935 28713 19947 28716
rect 19889 28707 19947 28713
rect 20346 28704 20352 28716
rect 20404 28704 20410 28756
rect 30374 28704 30380 28756
rect 30432 28744 30438 28756
rect 31021 28747 31079 28753
rect 31021 28744 31033 28747
rect 30432 28716 31033 28744
rect 30432 28704 30438 28716
rect 31021 28713 31033 28716
rect 31067 28713 31079 28747
rect 31021 28707 31079 28713
rect 32677 28747 32735 28753
rect 32677 28713 32689 28747
rect 32723 28744 32735 28747
rect 35342 28744 35348 28756
rect 32723 28716 35348 28744
rect 32723 28713 32735 28716
rect 32677 28707 32735 28713
rect 1946 28500 1952 28552
rect 2004 28540 2010 28552
rect 2682 28540 2688 28552
rect 2004 28512 2688 28540
rect 2004 28500 2010 28512
rect 2682 28500 2688 28512
rect 2740 28500 2746 28552
rect 3878 28500 3884 28552
rect 3936 28500 3942 28552
rect 4890 28500 4896 28552
rect 4948 28500 4954 28552
rect 19242 28500 19248 28552
rect 19300 28500 19306 28552
rect 31036 28540 31064 28707
rect 35342 28704 35348 28716
rect 35400 28704 35406 28756
rect 36814 28704 36820 28756
rect 36872 28704 36878 28756
rect 35360 28608 35388 28704
rect 35437 28611 35495 28617
rect 35437 28608 35449 28611
rect 35360 28580 35449 28608
rect 35437 28577 35449 28580
rect 35483 28577 35495 28611
rect 35437 28571 35495 28577
rect 31205 28543 31263 28549
rect 31205 28540 31217 28543
rect 31036 28512 31217 28540
rect 31205 28509 31217 28512
rect 31251 28509 31263 28543
rect 31205 28503 31263 28509
rect 34793 28543 34851 28549
rect 34793 28509 34805 28543
rect 34839 28540 34851 28543
rect 35158 28540 35164 28552
rect 34839 28512 35164 28540
rect 34839 28509 34851 28512
rect 34793 28503 34851 28509
rect 35158 28500 35164 28512
rect 35216 28500 35222 28552
rect 35526 28500 35532 28552
rect 35584 28540 35590 28552
rect 35693 28543 35751 28549
rect 35693 28540 35705 28543
rect 35584 28512 35705 28540
rect 35584 28500 35590 28512
rect 35693 28509 35705 28512
rect 35739 28509 35751 28543
rect 35693 28503 35751 28509
rect 2216 28475 2274 28481
rect 2216 28441 2228 28475
rect 2262 28472 2274 28475
rect 4908 28472 4936 28500
rect 2262 28444 4936 28472
rect 2262 28441 2274 28444
rect 2216 28435 2274 28441
rect 4430 28364 4436 28416
rect 4488 28364 4494 28416
rect 35345 28407 35403 28413
rect 35345 28373 35357 28407
rect 35391 28404 35403 28407
rect 35526 28404 35532 28416
rect 35391 28376 35532 28404
rect 35391 28373 35403 28376
rect 35345 28367 35403 28373
rect 35526 28364 35532 28376
rect 35584 28364 35590 28416
rect 1104 28314 37812 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 37812 28314
rect 1104 28240 37812 28262
rect 4430 28160 4436 28212
rect 4488 28160 4494 28212
rect 35526 28160 35532 28212
rect 35584 28160 35590 28212
rect 2774 28092 2780 28144
rect 2832 28132 2838 28144
rect 3605 28135 3663 28141
rect 3605 28132 3617 28135
rect 2832 28104 3617 28132
rect 2832 28092 2838 28104
rect 3605 28101 3617 28104
rect 3651 28101 3663 28135
rect 3605 28095 3663 28101
rect 2590 28024 2596 28076
rect 2648 28024 2654 28076
rect 4157 28067 4215 28073
rect 4157 28033 4169 28067
rect 4203 28064 4215 28067
rect 4448 28064 4476 28160
rect 4203 28036 4476 28064
rect 4203 28033 4215 28036
rect 4157 28027 4215 28033
rect 34790 28024 34796 28076
rect 34848 28064 34854 28076
rect 34977 28067 35035 28073
rect 34977 28064 34989 28067
rect 34848 28036 34989 28064
rect 34848 28024 34854 28036
rect 34977 28033 34989 28036
rect 35023 28033 35035 28067
rect 35544 28064 35572 28160
rect 36078 28092 36084 28144
rect 36136 28132 36142 28144
rect 36173 28135 36231 28141
rect 36173 28132 36185 28135
rect 36136 28104 36185 28132
rect 36136 28092 36142 28104
rect 36173 28101 36185 28104
rect 36219 28101 36231 28135
rect 36173 28095 36231 28101
rect 35805 28067 35863 28073
rect 35805 28064 35817 28067
rect 35544 28036 35817 28064
rect 34977 28027 35035 28033
rect 35805 28033 35817 28036
rect 35851 28033 35863 28067
rect 35805 28027 35863 28033
rect 1578 27956 1584 28008
rect 1636 27956 1642 28008
rect 35158 27956 35164 28008
rect 35216 27996 35222 28008
rect 35434 27996 35440 28008
rect 35216 27968 35440 27996
rect 35216 27956 35222 27968
rect 35434 27956 35440 27968
rect 35492 27996 35498 28008
rect 35621 27999 35679 28005
rect 35621 27996 35633 27999
rect 35492 27968 35633 27996
rect 35492 27956 35498 27968
rect 35621 27965 35633 27968
rect 35667 27965 35679 27999
rect 35621 27959 35679 27965
rect 1104 27770 37812 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 37812 27770
rect 1104 27696 37812 27718
rect 2498 27548 2504 27600
rect 2556 27588 2562 27600
rect 3789 27591 3847 27597
rect 3789 27588 3801 27591
rect 2556 27560 3801 27588
rect 2556 27548 2562 27560
rect 3789 27557 3801 27560
rect 3835 27557 3847 27591
rect 3789 27551 3847 27557
rect 3878 27548 3884 27600
rect 3936 27588 3942 27600
rect 4617 27591 4675 27597
rect 4617 27588 4629 27591
rect 3936 27560 4629 27588
rect 3936 27548 3942 27560
rect 4617 27557 4629 27560
rect 4663 27557 4675 27591
rect 4617 27551 4675 27557
rect 35161 27591 35219 27597
rect 35161 27557 35173 27591
rect 35207 27588 35219 27591
rect 35434 27588 35440 27600
rect 35207 27560 35440 27588
rect 35207 27557 35219 27560
rect 35161 27551 35219 27557
rect 35434 27548 35440 27560
rect 35492 27548 35498 27600
rect 2409 27523 2467 27529
rect 2409 27489 2421 27523
rect 2455 27520 2467 27523
rect 2590 27520 2596 27532
rect 2455 27492 2596 27520
rect 2455 27489 2467 27492
rect 2409 27483 2467 27489
rect 2590 27480 2596 27492
rect 2648 27480 2654 27532
rect 4982 27480 4988 27532
rect 5040 27480 5046 27532
rect 34514 27480 34520 27532
rect 34572 27520 34578 27532
rect 34793 27523 34851 27529
rect 34793 27520 34805 27523
rect 34572 27492 34805 27520
rect 34572 27480 34578 27492
rect 34793 27489 34805 27492
rect 34839 27520 34851 27523
rect 35802 27520 35808 27532
rect 34839 27492 35808 27520
rect 34839 27489 34851 27492
rect 34793 27483 34851 27489
rect 35802 27480 35808 27492
rect 35860 27480 35866 27532
rect 2685 27455 2743 27461
rect 2685 27421 2697 27455
rect 2731 27452 2743 27455
rect 2869 27455 2927 27461
rect 2869 27452 2881 27455
rect 2731 27424 2881 27452
rect 2731 27421 2743 27424
rect 2685 27415 2743 27421
rect 2869 27421 2881 27424
rect 2915 27421 2927 27455
rect 2869 27415 2927 27421
rect 3513 27455 3571 27461
rect 3513 27421 3525 27455
rect 3559 27452 3571 27455
rect 4338 27452 4344 27464
rect 3559 27424 4344 27452
rect 3559 27421 3571 27424
rect 3513 27415 3571 27421
rect 4338 27412 4344 27424
rect 4396 27412 4402 27464
rect 4433 27455 4491 27461
rect 4433 27421 4445 27455
rect 4479 27452 4491 27455
rect 4614 27452 4620 27464
rect 4479 27424 4620 27452
rect 4479 27421 4491 27424
rect 4433 27415 4491 27421
rect 4614 27412 4620 27424
rect 4672 27412 4678 27464
rect 35986 27412 35992 27464
rect 36044 27412 36050 27464
rect 36262 27412 36268 27464
rect 36320 27412 36326 27464
rect 3234 27344 3240 27396
rect 3292 27384 3298 27396
rect 35526 27384 35532 27396
rect 3292 27356 4568 27384
rect 3292 27344 3298 27356
rect 4540 27325 4568 27356
rect 35268 27356 35532 27384
rect 35268 27325 35296 27356
rect 35526 27344 35532 27356
rect 35584 27344 35590 27396
rect 37274 27344 37280 27396
rect 37332 27344 37338 27396
rect 4525 27319 4583 27325
rect 4525 27285 4537 27319
rect 4571 27285 4583 27319
rect 4525 27279 4583 27285
rect 35253 27319 35311 27325
rect 35253 27285 35265 27319
rect 35299 27285 35311 27319
rect 35253 27279 35311 27285
rect 35345 27319 35403 27325
rect 35345 27285 35357 27319
rect 35391 27316 35403 27319
rect 35434 27316 35440 27328
rect 35391 27288 35440 27316
rect 35391 27285 35403 27288
rect 35345 27279 35403 27285
rect 35434 27276 35440 27288
rect 35492 27276 35498 27328
rect 1104 27226 37812 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 37812 27226
rect 1104 27152 37812 27174
rect 3142 27072 3148 27124
rect 3200 27072 3206 27124
rect 3329 27115 3387 27121
rect 3329 27081 3341 27115
rect 3375 27112 3387 27115
rect 3786 27112 3792 27124
rect 3375 27084 3792 27112
rect 3375 27081 3387 27084
rect 3329 27075 3387 27081
rect 3786 27072 3792 27084
rect 3844 27072 3850 27124
rect 4338 27072 4344 27124
rect 4396 27072 4402 27124
rect 4614 27072 4620 27124
rect 4672 27112 4678 27124
rect 4801 27115 4859 27121
rect 4801 27112 4813 27115
rect 4672 27084 4813 27112
rect 4672 27072 4678 27084
rect 4801 27081 4813 27084
rect 4847 27081 4859 27115
rect 4801 27075 4859 27081
rect 13446 27072 13452 27124
rect 13504 27072 13510 27124
rect 16761 27115 16819 27121
rect 16761 27112 16773 27115
rect 16546 27084 16773 27112
rect 3160 27044 3188 27072
rect 3421 27047 3479 27053
rect 3421 27044 3433 27047
rect 3160 27016 3433 27044
rect 3421 27013 3433 27016
rect 3467 27013 3479 27047
rect 4356 27044 4384 27072
rect 4982 27044 4988 27056
rect 4356 27016 4988 27044
rect 3421 27007 3479 27013
rect 4982 27004 4988 27016
rect 5040 27044 5046 27056
rect 5537 27047 5595 27053
rect 5537 27044 5549 27047
rect 5040 27016 5549 27044
rect 5040 27004 5046 27016
rect 5537 27013 5549 27016
rect 5583 27013 5595 27047
rect 9582 27044 9588 27056
rect 5537 27007 5595 27013
rect 8312 27016 9588 27044
rect 1946 26936 1952 26988
rect 2004 26936 2010 26988
rect 2216 26979 2274 26985
rect 2216 26945 2228 26979
rect 2262 26976 2274 26979
rect 3326 26976 3332 26988
rect 2262 26948 3332 26976
rect 2262 26945 2274 26948
rect 2216 26939 2274 26945
rect 3326 26936 3332 26948
rect 3384 26936 3390 26988
rect 3510 26936 3516 26988
rect 3568 26976 3574 26988
rect 3970 26976 3976 26988
rect 3568 26948 3976 26976
rect 3568 26936 3574 26948
rect 3970 26936 3976 26948
rect 4028 26936 4034 26988
rect 8312 26920 8340 27016
rect 9582 27004 9588 27016
rect 9640 27044 9646 27056
rect 9640 27016 14872 27044
rect 9640 27004 9646 27016
rect 14844 26985 14872 27016
rect 14573 26979 14631 26985
rect 14573 26945 14585 26979
rect 14619 26976 14631 26979
rect 14829 26979 14887 26985
rect 14619 26948 14780 26976
rect 14619 26945 14631 26948
rect 14573 26939 14631 26945
rect 4062 26868 4068 26920
rect 4120 26908 4126 26920
rect 4157 26911 4215 26917
rect 4157 26908 4169 26911
rect 4120 26880 4169 26908
rect 4120 26868 4126 26880
rect 4157 26877 4169 26880
rect 4203 26877 4215 26911
rect 4157 26871 4215 26877
rect 4890 26868 4896 26920
rect 4948 26868 4954 26920
rect 8294 26868 8300 26920
rect 8352 26868 8358 26920
rect 14752 26908 14780 26948
rect 14829 26945 14841 26979
rect 14875 26945 14887 26979
rect 14829 26939 14887 26945
rect 16546 26908 16574 27084
rect 16761 27081 16773 27084
rect 16807 27081 16819 27115
rect 16761 27075 16819 27081
rect 35434 27072 35440 27124
rect 35492 27072 35498 27124
rect 35526 27072 35532 27124
rect 35584 27072 35590 27124
rect 35986 27072 35992 27124
rect 36044 27112 36050 27124
rect 36817 27115 36875 27121
rect 36817 27112 36829 27115
rect 36044 27084 36829 27112
rect 36044 27072 36050 27084
rect 36817 27081 36829 27084
rect 36863 27081 36875 27115
rect 36817 27075 36875 27081
rect 19242 27044 19248 27056
rect 14752 26880 16574 26908
rect 16960 27016 19248 27044
rect 16960 26849 16988 27016
rect 19242 27004 19248 27016
rect 19300 27004 19306 27056
rect 35452 27044 35480 27072
rect 35268 27016 35480 27044
rect 35544 27044 35572 27072
rect 35682 27047 35740 27053
rect 35682 27044 35694 27047
rect 35544 27016 35694 27044
rect 35268 26985 35296 27016
rect 35682 27013 35694 27016
rect 35728 27013 35740 27047
rect 35682 27007 35740 27013
rect 17589 26979 17647 26985
rect 17589 26945 17601 26979
rect 17635 26976 17647 26979
rect 35253 26979 35311 26985
rect 17635 26948 17908 26976
rect 17635 26945 17647 26948
rect 17589 26939 17647 26945
rect 17221 26911 17279 26917
rect 17221 26877 17233 26911
rect 17267 26908 17279 26911
rect 17267 26880 17356 26908
rect 17267 26877 17279 26880
rect 17221 26871 17279 26877
rect 16945 26843 17003 26849
rect 16945 26809 16957 26843
rect 16991 26809 17003 26843
rect 16945 26803 17003 26809
rect 17328 26784 17356 26880
rect 17880 26784 17908 26948
rect 35253 26945 35265 26979
rect 35299 26945 35311 26979
rect 35253 26939 35311 26945
rect 35342 26936 35348 26988
rect 35400 26976 35406 26988
rect 35437 26979 35495 26985
rect 35437 26976 35449 26979
rect 35400 26948 35449 26976
rect 35400 26936 35406 26948
rect 35437 26945 35449 26948
rect 35483 26945 35495 26979
rect 35437 26939 35495 26945
rect 17310 26732 17316 26784
rect 17368 26772 17374 26784
rect 17405 26775 17463 26781
rect 17405 26772 17417 26775
rect 17368 26744 17417 26772
rect 17368 26732 17374 26744
rect 17405 26741 17417 26744
rect 17451 26741 17463 26775
rect 17405 26735 17463 26741
rect 17862 26732 17868 26784
rect 17920 26732 17926 26784
rect 34698 26732 34704 26784
rect 34756 26732 34762 26784
rect 1104 26682 37812 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 37812 26682
rect 1104 26608 37812 26630
rect 3326 26528 3332 26580
rect 3384 26528 3390 26580
rect 4433 26571 4491 26577
rect 4433 26537 4445 26571
rect 4479 26568 4491 26571
rect 4890 26568 4896 26580
rect 4479 26540 4896 26568
rect 4479 26537 4491 26540
rect 4433 26531 4491 26537
rect 4890 26528 4896 26540
rect 4948 26528 4954 26580
rect 31481 26571 31539 26577
rect 31481 26537 31493 26571
rect 31527 26568 31539 26571
rect 33502 26568 33508 26580
rect 31527 26540 33508 26568
rect 31527 26537 31539 26540
rect 31481 26531 31539 26537
rect 33502 26528 33508 26540
rect 33560 26528 33566 26580
rect 36262 26528 36268 26580
rect 36320 26528 36326 26580
rect 3344 26500 3372 26528
rect 4525 26503 4583 26509
rect 4525 26500 4537 26503
rect 3344 26472 4537 26500
rect 4525 26469 4537 26472
rect 4571 26469 4583 26503
rect 4525 26463 4583 26469
rect 1946 26392 1952 26444
rect 2004 26392 2010 26444
rect 5261 26435 5319 26441
rect 5261 26432 5273 26435
rect 2976 26404 5273 26432
rect 1964 26364 1992 26392
rect 2976 26364 3004 26404
rect 5261 26401 5273 26404
rect 5307 26401 5319 26435
rect 5261 26395 5319 26401
rect 34698 26392 34704 26444
rect 34756 26432 34762 26444
rect 35345 26435 35403 26441
rect 35345 26432 35357 26435
rect 34756 26404 35357 26432
rect 34756 26392 34762 26404
rect 35345 26401 35357 26404
rect 35391 26401 35403 26435
rect 36280 26432 36308 26528
rect 36449 26435 36507 26441
rect 36449 26432 36461 26435
rect 36280 26404 36461 26432
rect 35345 26395 35403 26401
rect 36449 26401 36461 26404
rect 36495 26401 36507 26435
rect 36449 26395 36507 26401
rect 1964 26336 3004 26364
rect 3234 26324 3240 26376
rect 3292 26324 3298 26376
rect 3789 26367 3847 26373
rect 3789 26364 3801 26367
rect 3344 26336 3801 26364
rect 2216 26299 2274 26305
rect 2216 26265 2228 26299
rect 2262 26296 2274 26299
rect 3252 26296 3280 26324
rect 2262 26268 3280 26296
rect 2262 26265 2274 26268
rect 2216 26259 2274 26265
rect 3344 26237 3372 26336
rect 3789 26333 3801 26336
rect 3835 26333 3847 26367
rect 3789 26327 3847 26333
rect 4709 26367 4767 26373
rect 4709 26333 4721 26367
rect 4755 26364 4767 26367
rect 4798 26364 4804 26376
rect 4755 26336 4804 26364
rect 4755 26333 4767 26336
rect 4709 26327 4767 26333
rect 4798 26324 4804 26336
rect 4856 26324 4862 26376
rect 4893 26367 4951 26373
rect 4893 26333 4905 26367
rect 4939 26364 4951 26367
rect 6914 26364 6920 26376
rect 4939 26336 6920 26364
rect 4939 26333 4951 26336
rect 4893 26327 4951 26333
rect 6914 26324 6920 26336
rect 6972 26324 6978 26376
rect 28994 26324 29000 26376
rect 29052 26364 29058 26376
rect 30837 26367 30895 26373
rect 30837 26364 30849 26367
rect 29052 26336 30849 26364
rect 29052 26324 29058 26336
rect 30837 26333 30849 26336
rect 30883 26333 30895 26367
rect 30837 26327 30895 26333
rect 35989 26367 36047 26373
rect 35989 26333 36001 26367
rect 36035 26364 36047 26367
rect 36173 26367 36231 26373
rect 36173 26364 36185 26367
rect 36035 26336 36185 26364
rect 36035 26333 36047 26336
rect 35989 26327 36047 26333
rect 36173 26333 36185 26336
rect 36219 26333 36231 26367
rect 36173 26327 36231 26333
rect 7009 26299 7067 26305
rect 7009 26265 7021 26299
rect 7055 26296 7067 26299
rect 7377 26299 7435 26305
rect 7377 26296 7389 26299
rect 7055 26268 7389 26296
rect 7055 26265 7067 26268
rect 7009 26259 7067 26265
rect 7377 26265 7389 26268
rect 7423 26296 7435 26299
rect 8386 26296 8392 26308
rect 7423 26268 8392 26296
rect 7423 26265 7435 26268
rect 7377 26259 7435 26265
rect 8386 26256 8392 26268
rect 8444 26256 8450 26308
rect 17310 26256 17316 26308
rect 17368 26256 17374 26308
rect 34977 26299 35035 26305
rect 34977 26265 34989 26299
rect 35023 26296 35035 26299
rect 35023 26268 35057 26296
rect 35023 26265 35035 26268
rect 34977 26259 35035 26265
rect 3329 26231 3387 26237
rect 3329 26197 3341 26231
rect 3375 26197 3387 26231
rect 3329 26191 3387 26197
rect 34514 26188 34520 26240
rect 34572 26228 34578 26240
rect 34992 26228 35020 26259
rect 34572 26200 35020 26228
rect 34572 26188 34578 26200
rect 1104 26138 37812 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 37812 26138
rect 1104 26064 37812 26086
rect 8294 25984 8300 26036
rect 8352 25984 8358 26036
rect 20346 25984 20352 26036
rect 20404 25984 20410 26036
rect 2685 25891 2743 25897
rect 2685 25857 2697 25891
rect 2731 25888 2743 25891
rect 2774 25888 2780 25900
rect 2731 25860 2780 25888
rect 2731 25857 2743 25860
rect 2685 25851 2743 25857
rect 2774 25848 2780 25860
rect 2832 25848 2838 25900
rect 8386 25848 8392 25900
rect 8444 25888 8450 25900
rect 9585 25891 9643 25897
rect 9585 25888 9597 25891
rect 8444 25860 9597 25888
rect 8444 25848 8450 25860
rect 9585 25857 9597 25860
rect 9631 25888 9643 25891
rect 9631 25860 9996 25888
rect 9631 25857 9643 25860
rect 9585 25851 9643 25857
rect 934 25780 940 25832
rect 992 25820 998 25832
rect 1581 25823 1639 25829
rect 1581 25820 1593 25823
rect 992 25792 1593 25820
rect 992 25780 998 25792
rect 1581 25789 1593 25792
rect 1627 25789 1639 25823
rect 1581 25783 1639 25789
rect 2961 25823 3019 25829
rect 2961 25789 2973 25823
rect 3007 25820 3019 25823
rect 3605 25823 3663 25829
rect 3605 25820 3617 25823
rect 3007 25792 3617 25820
rect 3007 25789 3019 25792
rect 2961 25783 3019 25789
rect 3605 25789 3617 25792
rect 3651 25789 3663 25823
rect 3605 25783 3663 25789
rect 3694 25780 3700 25832
rect 3752 25820 3758 25832
rect 4157 25823 4215 25829
rect 4157 25820 4169 25823
rect 3752 25792 4169 25820
rect 3752 25780 3758 25792
rect 4157 25789 4169 25792
rect 4203 25789 4215 25823
rect 4157 25783 4215 25789
rect 4798 25780 4804 25832
rect 4856 25820 4862 25832
rect 5353 25823 5411 25829
rect 5353 25820 5365 25823
rect 4856 25792 5365 25820
rect 4856 25780 4862 25792
rect 5353 25789 5365 25792
rect 5399 25789 5411 25823
rect 5353 25783 5411 25789
rect 4525 25755 4583 25761
rect 4525 25721 4537 25755
rect 4571 25752 4583 25755
rect 4614 25752 4620 25764
rect 4571 25724 4620 25752
rect 4571 25721 4583 25724
rect 4525 25715 4583 25721
rect 4614 25712 4620 25724
rect 4672 25712 4678 25764
rect 4982 25712 4988 25764
rect 5040 25712 5046 25764
rect 9968 25761 9996 25860
rect 35894 25848 35900 25900
rect 35952 25848 35958 25900
rect 19426 25780 19432 25832
rect 19484 25820 19490 25832
rect 19705 25823 19763 25829
rect 19705 25820 19717 25823
rect 19484 25792 19717 25820
rect 19484 25780 19490 25792
rect 19705 25789 19717 25792
rect 19751 25789 19763 25823
rect 19705 25783 19763 25789
rect 34425 25823 34483 25829
rect 34425 25789 34437 25823
rect 34471 25820 34483 25823
rect 34514 25820 34520 25832
rect 34471 25792 34520 25820
rect 34471 25789 34483 25792
rect 34425 25783 34483 25789
rect 34514 25780 34520 25792
rect 34572 25780 34578 25832
rect 35618 25780 35624 25832
rect 35676 25780 35682 25832
rect 36909 25823 36967 25829
rect 36909 25789 36921 25823
rect 36955 25820 36967 25823
rect 37458 25820 37464 25832
rect 36955 25792 37464 25820
rect 36955 25789 36967 25792
rect 36909 25783 36967 25789
rect 37458 25780 37464 25792
rect 37516 25780 37522 25832
rect 9953 25755 10011 25761
rect 9953 25721 9965 25755
rect 9999 25752 10011 25755
rect 20254 25752 20260 25764
rect 9999 25724 20260 25752
rect 9999 25721 10011 25724
rect 9953 25715 10011 25721
rect 20254 25712 20260 25724
rect 20312 25752 20318 25764
rect 28442 25752 28448 25764
rect 20312 25724 28448 25752
rect 20312 25712 20318 25724
rect 28442 25712 28448 25724
rect 28500 25712 28506 25764
rect 34698 25712 34704 25764
rect 34756 25712 34762 25764
rect 34790 25712 34796 25764
rect 34848 25752 34854 25764
rect 34977 25755 35035 25761
rect 34977 25752 34989 25755
rect 34848 25724 34989 25752
rect 34848 25712 34854 25724
rect 34977 25721 34989 25724
rect 35023 25721 35035 25755
rect 34977 25715 35035 25721
rect 3513 25687 3571 25693
rect 3513 25653 3525 25687
rect 3559 25684 3571 25687
rect 3786 25684 3792 25696
rect 3559 25656 3792 25684
rect 3559 25653 3571 25656
rect 3513 25647 3571 25653
rect 3786 25644 3792 25656
rect 3844 25644 3850 25696
rect 4341 25687 4399 25693
rect 4341 25653 4353 25687
rect 4387 25684 4399 25687
rect 4706 25684 4712 25696
rect 4387 25656 4712 25684
rect 4387 25653 4399 25656
rect 4341 25647 4399 25653
rect 4706 25644 4712 25656
rect 4764 25644 4770 25696
rect 4890 25644 4896 25696
rect 4948 25644 4954 25696
rect 34885 25687 34943 25693
rect 34885 25653 34897 25687
rect 34931 25684 34943 25687
rect 35342 25684 35348 25696
rect 34931 25656 35348 25684
rect 34931 25653 34943 25656
rect 34885 25647 34943 25653
rect 35342 25644 35348 25656
rect 35400 25644 35406 25696
rect 1104 25594 37812 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 37812 25594
rect 1104 25520 37812 25542
rect 3329 25483 3387 25489
rect 3329 25449 3341 25483
rect 3375 25480 3387 25483
rect 3694 25480 3700 25492
rect 3375 25452 3700 25480
rect 3375 25449 3387 25452
rect 3329 25443 3387 25449
rect 3694 25440 3700 25452
rect 3752 25440 3758 25492
rect 4890 25440 4896 25492
rect 4948 25440 4954 25492
rect 31573 25483 31631 25489
rect 31573 25449 31585 25483
rect 31619 25480 31631 25483
rect 32122 25480 32128 25492
rect 31619 25452 32128 25480
rect 31619 25449 31631 25452
rect 31573 25443 31631 25449
rect 32122 25440 32128 25452
rect 32180 25440 32186 25492
rect 35342 25440 35348 25492
rect 35400 25440 35406 25492
rect 35618 25440 35624 25492
rect 35676 25480 35682 25492
rect 36817 25483 36875 25489
rect 36817 25480 36829 25483
rect 35676 25452 36829 25480
rect 35676 25440 35682 25452
rect 36817 25449 36829 25452
rect 36863 25449 36875 25483
rect 36817 25443 36875 25449
rect 4908 25344 4936 25440
rect 3528 25316 4936 25344
rect 35360 25344 35388 25440
rect 35360 25316 35572 25344
rect 1946 25236 1952 25288
rect 2004 25236 2010 25288
rect 2216 25279 2274 25285
rect 2216 25245 2228 25279
rect 2262 25276 2274 25279
rect 3528 25276 3556 25316
rect 2262 25248 3556 25276
rect 2262 25245 2274 25248
rect 2216 25239 2274 25245
rect 3786 25236 3792 25288
rect 3844 25276 3850 25288
rect 4154 25276 4160 25288
rect 3844 25248 4160 25276
rect 3844 25236 3850 25248
rect 4154 25236 4160 25248
rect 4212 25236 4218 25288
rect 29638 25236 29644 25288
rect 29696 25276 29702 25288
rect 30929 25279 30987 25285
rect 30929 25276 30941 25279
rect 29696 25248 30941 25276
rect 29696 25236 29702 25248
rect 30929 25245 30941 25248
rect 30975 25245 30987 25279
rect 30929 25239 30987 25245
rect 34793 25279 34851 25285
rect 34793 25245 34805 25279
rect 34839 25276 34851 25279
rect 35158 25276 35164 25288
rect 34839 25248 35164 25276
rect 34839 25245 34851 25248
rect 34793 25239 34851 25245
rect 35158 25236 35164 25248
rect 35216 25236 35222 25288
rect 35434 25236 35440 25288
rect 35492 25236 35498 25288
rect 35544 25276 35572 25316
rect 35693 25279 35751 25285
rect 35693 25276 35705 25279
rect 35544 25248 35705 25276
rect 35693 25245 35705 25248
rect 35739 25245 35751 25279
rect 35693 25239 35751 25245
rect 4430 25100 4436 25152
rect 4488 25100 4494 25152
rect 35342 25100 35348 25152
rect 35400 25100 35406 25152
rect 1104 25050 37812 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 37812 25050
rect 1104 24976 37812 24998
rect 35158 24896 35164 24948
rect 35216 24936 35222 24948
rect 35526 24936 35532 24948
rect 35216 24908 35532 24936
rect 35216 24896 35222 24908
rect 35526 24896 35532 24908
rect 35584 24936 35590 24948
rect 35621 24939 35679 24945
rect 35621 24936 35633 24939
rect 35584 24908 35633 24936
rect 35584 24896 35590 24908
rect 35621 24905 35633 24908
rect 35667 24905 35679 24939
rect 35621 24899 35679 24905
rect 2774 24828 2780 24880
rect 2832 24868 2838 24880
rect 3605 24871 3663 24877
rect 3605 24868 3617 24871
rect 2832 24840 3617 24868
rect 2832 24828 2838 24840
rect 3605 24837 3617 24840
rect 3651 24837 3663 24871
rect 3605 24831 3663 24837
rect 35894 24828 35900 24880
rect 35952 24868 35958 24880
rect 35952 24840 36216 24868
rect 35952 24828 35958 24840
rect 2590 24760 2596 24812
rect 2648 24760 2654 24812
rect 4157 24803 4215 24809
rect 4157 24769 4169 24803
rect 4203 24800 4215 24803
rect 4430 24800 4436 24812
rect 4203 24772 4436 24800
rect 4203 24769 4215 24772
rect 4157 24763 4215 24769
rect 4430 24760 4436 24772
rect 4488 24760 4494 24812
rect 34790 24760 34796 24812
rect 34848 24800 34854 24812
rect 34977 24803 35035 24809
rect 34977 24800 34989 24803
rect 34848 24772 34989 24800
rect 34848 24760 34854 24772
rect 34977 24769 34989 24772
rect 35023 24769 35035 24803
rect 34977 24763 35035 24769
rect 35342 24760 35348 24812
rect 35400 24800 35406 24812
rect 36188 24809 36216 24840
rect 35805 24803 35863 24809
rect 35805 24800 35817 24803
rect 35400 24772 35817 24800
rect 35400 24760 35406 24772
rect 35805 24769 35817 24772
rect 35851 24769 35863 24803
rect 35805 24763 35863 24769
rect 36173 24803 36231 24809
rect 36173 24769 36185 24803
rect 36219 24769 36231 24803
rect 36173 24763 36231 24769
rect 934 24692 940 24744
rect 992 24732 998 24744
rect 1581 24735 1639 24741
rect 1581 24732 1593 24735
rect 992 24704 1593 24732
rect 992 24692 998 24704
rect 1581 24701 1593 24704
rect 1627 24701 1639 24735
rect 1581 24695 1639 24701
rect 4614 24692 4620 24744
rect 4672 24732 4678 24744
rect 4798 24732 4804 24744
rect 4672 24704 4804 24732
rect 4672 24692 4678 24704
rect 4798 24692 4804 24704
rect 4856 24692 4862 24744
rect 4154 24624 4160 24676
rect 4212 24664 4218 24676
rect 4433 24667 4491 24673
rect 4433 24664 4445 24667
rect 4212 24636 4445 24664
rect 4212 24624 4218 24636
rect 4433 24633 4445 24636
rect 4479 24633 4491 24667
rect 4433 24627 4491 24633
rect 3234 24556 3240 24608
rect 3292 24596 3298 24608
rect 4341 24599 4399 24605
rect 4341 24596 4353 24599
rect 3292 24568 4353 24596
rect 3292 24556 3298 24568
rect 4341 24565 4353 24568
rect 4387 24565 4399 24599
rect 4341 24559 4399 24565
rect 1104 24506 37812 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 37812 24506
rect 1104 24432 37812 24454
rect 35161 24327 35219 24333
rect 35161 24293 35173 24327
rect 35207 24324 35219 24327
rect 35526 24324 35532 24336
rect 35207 24296 35532 24324
rect 35207 24293 35219 24296
rect 35161 24287 35219 24293
rect 35526 24284 35532 24296
rect 35584 24284 35590 24336
rect 2774 24148 2780 24200
rect 2832 24188 2838 24200
rect 3329 24191 3387 24197
rect 3329 24188 3341 24191
rect 2832 24160 3341 24188
rect 2832 24148 2838 24160
rect 3329 24157 3341 24160
rect 3375 24157 3387 24191
rect 3329 24151 3387 24157
rect 3786 24148 3792 24200
rect 3844 24148 3850 24200
rect 4706 24148 4712 24200
rect 4764 24148 4770 24200
rect 35986 24148 35992 24200
rect 36044 24148 36050 24200
rect 36262 24148 36268 24200
rect 36320 24148 36326 24200
rect 3084 24123 3142 24129
rect 3084 24089 3096 24123
rect 3130 24120 3142 24123
rect 4724 24120 4752 24148
rect 3130 24092 4752 24120
rect 3130 24089 3142 24092
rect 3084 24083 3142 24089
rect 34514 24080 34520 24132
rect 34572 24120 34578 24132
rect 34793 24123 34851 24129
rect 34793 24120 34805 24123
rect 34572 24092 34805 24120
rect 34572 24080 34578 24092
rect 34793 24089 34805 24092
rect 34839 24120 34851 24123
rect 36078 24120 36084 24132
rect 34839 24092 36084 24120
rect 34839 24089 34851 24092
rect 34793 24083 34851 24089
rect 36078 24080 36084 24092
rect 36136 24080 36142 24132
rect 37274 24080 37280 24132
rect 37332 24080 37338 24132
rect 1949 24055 2007 24061
rect 1949 24021 1961 24055
rect 1995 24052 2007 24055
rect 2958 24052 2964 24064
rect 1995 24024 2964 24052
rect 1995 24021 2007 24024
rect 1949 24015 2007 24021
rect 2958 24012 2964 24024
rect 3016 24012 3022 24064
rect 4430 24012 4436 24064
rect 4488 24012 4494 24064
rect 35250 24012 35256 24064
rect 35308 24012 35314 24064
rect 35342 24012 35348 24064
rect 35400 24012 35406 24064
rect 1104 23962 37812 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 37812 23962
rect 1104 23888 37812 23910
rect 3234 23848 3240 23860
rect 2231 23820 3240 23848
rect 2231 23789 2259 23820
rect 3234 23808 3240 23820
rect 3292 23808 3298 23860
rect 3329 23851 3387 23857
rect 3329 23817 3341 23851
rect 3375 23848 3387 23851
rect 3786 23848 3792 23860
rect 3375 23820 3792 23848
rect 3375 23817 3387 23820
rect 3329 23811 3387 23817
rect 3786 23808 3792 23820
rect 3844 23808 3850 23860
rect 4062 23808 4068 23860
rect 4120 23808 4126 23860
rect 4430 23808 4436 23860
rect 4488 23808 4494 23860
rect 35250 23808 35256 23860
rect 35308 23848 35314 23860
rect 35308 23820 35725 23848
rect 35308 23808 35314 23820
rect 2216 23783 2274 23789
rect 2216 23749 2228 23783
rect 2262 23749 2274 23783
rect 2216 23743 2274 23749
rect 4448 23712 4476 23808
rect 35342 23740 35348 23792
rect 35400 23740 35406 23792
rect 35697 23789 35725 23820
rect 35986 23808 35992 23860
rect 36044 23848 36050 23860
rect 36817 23851 36875 23857
rect 36817 23848 36829 23851
rect 36044 23820 36829 23848
rect 36044 23808 36050 23820
rect 36817 23817 36829 23820
rect 36863 23817 36875 23851
rect 36817 23811 36875 23817
rect 35682 23783 35740 23789
rect 35682 23749 35694 23783
rect 35728 23749 35740 23783
rect 35682 23743 35740 23749
rect 4709 23715 4767 23721
rect 4709 23712 4721 23715
rect 4448 23684 4721 23712
rect 4709 23681 4721 23684
rect 4755 23681 4767 23715
rect 4709 23675 4767 23681
rect 34793 23715 34851 23721
rect 34793 23681 34805 23715
rect 34839 23712 34851 23715
rect 35360 23712 35388 23740
rect 34839 23684 35388 23712
rect 34839 23681 34851 23684
rect 34793 23675 34851 23681
rect 1946 23604 1952 23656
rect 2004 23604 2010 23656
rect 3418 23604 3424 23656
rect 3476 23604 3482 23656
rect 35434 23604 35440 23656
rect 35492 23604 35498 23656
rect 1964 23508 1992 23604
rect 2682 23508 2688 23520
rect 1964 23480 2688 23508
rect 2682 23468 2688 23480
rect 2740 23468 2746 23520
rect 4062 23468 4068 23520
rect 4120 23508 4126 23520
rect 4157 23511 4215 23517
rect 4157 23508 4169 23511
rect 4120 23480 4169 23508
rect 4120 23468 4126 23480
rect 4157 23477 4169 23480
rect 4203 23477 4215 23511
rect 4157 23471 4215 23477
rect 35345 23511 35403 23517
rect 35345 23477 35357 23511
rect 35391 23508 35403 23511
rect 35618 23508 35624 23520
rect 35391 23480 35624 23508
rect 35391 23477 35403 23480
rect 35345 23471 35403 23477
rect 35618 23468 35624 23480
rect 35676 23468 35682 23520
rect 1104 23418 37812 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 37812 23418
rect 1104 23344 37812 23366
rect 4062 23304 4068 23316
rect 3528 23276 4068 23304
rect 2409 23171 2467 23177
rect 2409 23137 2421 23171
rect 2455 23168 2467 23171
rect 2590 23168 2596 23180
rect 2455 23140 2596 23168
rect 2455 23137 2467 23140
rect 2409 23131 2467 23137
rect 2590 23128 2596 23140
rect 2648 23128 2654 23180
rect 3528 23177 3556 23276
rect 4062 23264 4068 23276
rect 4120 23264 4126 23316
rect 28994 23264 29000 23316
rect 29052 23264 29058 23316
rect 3513 23171 3571 23177
rect 3513 23137 3525 23171
rect 3559 23137 3571 23171
rect 3513 23131 3571 23137
rect 36262 23128 36268 23180
rect 36320 23168 36326 23180
rect 36449 23171 36507 23177
rect 36449 23168 36461 23171
rect 36320 23140 36461 23168
rect 36320 23128 36326 23140
rect 36449 23137 36461 23140
rect 36495 23137 36507 23171
rect 36449 23131 36507 23137
rect 2685 23103 2743 23109
rect 2685 23069 2697 23103
rect 2731 23100 2743 23103
rect 2869 23103 2927 23109
rect 2869 23100 2881 23103
rect 2731 23072 2881 23100
rect 2731 23069 2743 23072
rect 2685 23063 2743 23069
rect 2869 23069 2881 23072
rect 2915 23069 2927 23103
rect 2869 23063 2927 23069
rect 28350 23060 28356 23112
rect 28408 23060 28414 23112
rect 35437 23103 35495 23109
rect 35437 23069 35449 23103
rect 35483 23100 35495 23103
rect 35618 23100 35624 23112
rect 35483 23072 35624 23100
rect 35483 23069 35495 23072
rect 35437 23063 35495 23069
rect 35618 23060 35624 23072
rect 35676 23060 35682 23112
rect 35989 23103 36047 23109
rect 35989 23069 36001 23103
rect 36035 23100 36047 23103
rect 36173 23103 36231 23109
rect 36173 23100 36185 23103
rect 36035 23072 36185 23100
rect 36035 23069 36047 23072
rect 35989 23063 36047 23069
rect 36173 23069 36185 23072
rect 36219 23069 36231 23103
rect 36173 23063 36231 23069
rect 1104 22874 37812 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 37812 22874
rect 1104 22800 37812 22822
rect 36078 22720 36084 22772
rect 36136 22720 36142 22772
rect 2590 22584 2596 22636
rect 2648 22584 2654 22636
rect 1578 22516 1584 22568
rect 1636 22516 1642 22568
rect 2958 22516 2964 22568
rect 3016 22556 3022 22568
rect 3421 22559 3479 22565
rect 3421 22556 3433 22559
rect 3016 22528 3433 22556
rect 3016 22516 3022 22528
rect 3421 22525 3433 22528
rect 3467 22525 3479 22559
rect 3421 22519 3479 22525
rect 4062 22516 4068 22568
rect 4120 22556 4126 22568
rect 4614 22556 4620 22568
rect 4120 22528 4620 22556
rect 4120 22516 4126 22528
rect 4614 22516 4620 22528
rect 4672 22516 4678 22568
rect 36446 22516 36452 22568
rect 36504 22516 36510 22568
rect 3789 22491 3847 22497
rect 3789 22457 3801 22491
rect 3835 22488 3847 22491
rect 4154 22488 4160 22500
rect 3835 22460 4160 22488
rect 3835 22457 3847 22460
rect 3789 22451 3847 22457
rect 4154 22448 4160 22460
rect 4212 22448 4218 22500
rect 2866 22380 2872 22432
rect 2924 22380 2930 22432
rect 3602 22380 3608 22432
rect 3660 22380 3666 22432
rect 37090 22380 37096 22432
rect 37148 22380 37154 22432
rect 1104 22330 37812 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 37812 22330
rect 1104 22256 37812 22278
rect 35618 22108 35624 22160
rect 35676 22108 35682 22160
rect 35989 22083 36047 22089
rect 35989 22049 36001 22083
rect 36035 22080 36047 22083
rect 36078 22080 36084 22092
rect 36035 22052 36084 22080
rect 36035 22049 36047 22052
rect 35989 22043 36047 22049
rect 36078 22040 36084 22052
rect 36136 22040 36142 22092
rect 2774 21972 2780 22024
rect 2832 22012 2838 22024
rect 3329 22015 3387 22021
rect 3329 22012 3341 22015
rect 2832 21984 3341 22012
rect 2832 21972 2838 21984
rect 3329 21981 3341 21984
rect 3375 21981 3387 22015
rect 3329 21975 3387 21981
rect 3602 21972 3608 22024
rect 3660 21972 3666 22024
rect 4433 22015 4491 22021
rect 4433 21981 4445 22015
rect 4479 22012 4491 22015
rect 4479 21984 4660 22012
rect 4479 21981 4491 21984
rect 4433 21975 4491 21981
rect 2958 21904 2964 21956
rect 3016 21904 3022 21956
rect 3084 21947 3142 21953
rect 3084 21913 3096 21947
rect 3130 21944 3142 21947
rect 3620 21944 3648 21972
rect 3130 21916 3648 21944
rect 3130 21913 3142 21916
rect 3084 21907 3142 21913
rect 1949 21879 2007 21885
rect 1949 21845 1961 21879
rect 1995 21876 2007 21879
rect 2976 21876 3004 21904
rect 4632 21888 4660 21984
rect 19426 21972 19432 22024
rect 19484 21972 19490 22024
rect 20717 22015 20775 22021
rect 20717 21981 20729 22015
rect 20763 22012 20775 22015
rect 20763 21984 21128 22012
rect 20763 21981 20775 21984
rect 20717 21975 20775 21981
rect 1995 21848 3004 21876
rect 1995 21845 2007 21848
rect 1949 21839 2007 21845
rect 3786 21836 3792 21888
rect 3844 21836 3850 21888
rect 4614 21836 4620 21888
rect 4672 21836 4678 21888
rect 19337 21879 19395 21885
rect 19337 21845 19349 21879
rect 19383 21876 19395 21879
rect 19444 21876 19472 21972
rect 20346 21904 20352 21956
rect 20404 21944 20410 21956
rect 20450 21947 20508 21953
rect 20450 21944 20462 21947
rect 20404 21916 20462 21944
rect 20404 21904 20410 21916
rect 20450 21913 20462 21916
rect 20496 21913 20508 21947
rect 20450 21907 20508 21913
rect 21100 21885 21128 21984
rect 24118 21972 24124 22024
rect 24176 22012 24182 22024
rect 36173 22015 36231 22021
rect 36173 22012 36185 22015
rect 24176 21984 36185 22012
rect 24176 21972 24182 21984
rect 36173 21981 36185 21984
rect 36219 21981 36231 22015
rect 36173 21975 36231 21981
rect 36538 21904 36544 21956
rect 36596 21904 36602 21956
rect 19383 21848 19472 21876
rect 21085 21879 21143 21885
rect 19383 21845 19395 21848
rect 19337 21839 19395 21845
rect 21085 21845 21097 21879
rect 21131 21876 21143 21879
rect 28166 21876 28172 21888
rect 21131 21848 28172 21876
rect 21131 21845 21143 21848
rect 21085 21839 21143 21845
rect 28166 21836 28172 21848
rect 28224 21836 28230 21888
rect 35526 21836 35532 21888
rect 35584 21836 35590 21888
rect 1104 21786 37812 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 37812 21786
rect 1104 21712 37812 21734
rect 3786 21632 3792 21684
rect 3844 21632 3850 21684
rect 29638 21632 29644 21684
rect 29696 21632 29702 21684
rect 29914 21632 29920 21684
rect 29972 21632 29978 21684
rect 36538 21672 36544 21684
rect 35912 21644 36544 21672
rect 2317 21607 2375 21613
rect 2317 21573 2329 21607
rect 2363 21604 2375 21607
rect 2590 21604 2596 21616
rect 2363 21576 2596 21604
rect 2363 21573 2375 21576
rect 2317 21567 2375 21573
rect 2590 21564 2596 21576
rect 2648 21564 2654 21616
rect 3804 21604 3832 21632
rect 2700 21576 3832 21604
rect 2700 21545 2728 21576
rect 28166 21564 28172 21616
rect 28224 21604 28230 21616
rect 29932 21604 29960 21632
rect 28224 21576 29960 21604
rect 28224 21564 28230 21576
rect 2685 21539 2743 21545
rect 2685 21505 2697 21539
rect 2731 21505 2743 21539
rect 2685 21499 2743 21505
rect 2866 21496 2872 21548
rect 2924 21496 2930 21548
rect 3513 21539 3571 21545
rect 3513 21505 3525 21539
rect 3559 21536 3571 21539
rect 28184 21536 28212 21564
rect 35912 21545 35940 21644
rect 36538 21632 36544 21644
rect 36596 21632 36602 21684
rect 36909 21607 36967 21613
rect 36909 21573 36921 21607
rect 36955 21604 36967 21607
rect 37458 21604 37464 21616
rect 36955 21576 37464 21604
rect 36955 21573 36967 21576
rect 36909 21567 36967 21573
rect 37458 21564 37464 21576
rect 37516 21564 37522 21616
rect 28261 21539 28319 21545
rect 28261 21536 28273 21539
rect 3559 21508 4660 21536
rect 28184 21508 28273 21536
rect 3559 21505 3571 21508
rect 3513 21499 3571 21505
rect 4632 21480 4660 21508
rect 28261 21505 28273 21508
rect 28307 21505 28319 21539
rect 28517 21539 28575 21545
rect 28517 21536 28529 21539
rect 28261 21499 28319 21505
rect 28368 21508 28529 21536
rect 4062 21428 4068 21480
rect 4120 21428 4126 21480
rect 4614 21428 4620 21480
rect 4672 21428 4678 21480
rect 27522 21428 27528 21480
rect 27580 21468 27586 21480
rect 28368 21468 28396 21508
rect 28517 21505 28529 21508
rect 28563 21505 28575 21539
rect 28517 21499 28575 21505
rect 35897 21539 35955 21545
rect 35897 21505 35909 21539
rect 35943 21505 35955 21539
rect 35897 21499 35955 21505
rect 27580 21440 28396 21468
rect 27580 21428 27586 21440
rect 3789 21403 3847 21409
rect 3789 21369 3801 21403
rect 3835 21400 3847 21403
rect 3970 21400 3976 21412
rect 3835 21372 3976 21400
rect 3835 21369 3847 21372
rect 3789 21363 3847 21369
rect 3970 21360 3976 21372
rect 4028 21360 4034 21412
rect 3602 21292 3608 21344
rect 3660 21292 3666 21344
rect 1104 21242 37812 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 37812 21242
rect 1104 21168 37812 21190
rect 36817 21131 36875 21137
rect 36817 21128 36829 21131
rect 35268 21100 36829 21128
rect 4614 21020 4620 21072
rect 4672 21020 4678 21072
rect 4062 20952 4068 21004
rect 4120 20992 4126 21004
rect 4985 20995 5043 21001
rect 4985 20992 4997 20995
rect 4120 20964 4997 20992
rect 4120 20952 4126 20964
rect 4985 20961 4997 20964
rect 5031 20961 5043 20995
rect 4985 20955 5043 20961
rect 34793 20995 34851 21001
rect 34793 20961 34805 20995
rect 34839 20992 34851 20995
rect 35268 20992 35296 21100
rect 36817 21097 36829 21100
rect 36863 21097 36875 21131
rect 36817 21091 36875 21097
rect 34839 20964 35296 20992
rect 34839 20961 34851 20964
rect 34793 20955 34851 20961
rect 35434 20952 35440 21004
rect 35492 20952 35498 21004
rect 2685 20927 2743 20933
rect 2685 20893 2697 20927
rect 2731 20924 2743 20927
rect 2866 20924 2872 20936
rect 2731 20896 2872 20924
rect 2731 20893 2743 20896
rect 2685 20887 2743 20893
rect 2866 20884 2872 20896
rect 2924 20884 2930 20936
rect 2961 20927 3019 20933
rect 2961 20893 2973 20927
rect 3007 20924 3019 20927
rect 3789 20927 3847 20933
rect 3789 20924 3801 20927
rect 3007 20896 3801 20924
rect 3007 20893 3019 20896
rect 2961 20887 3019 20893
rect 3789 20893 3801 20896
rect 3835 20893 3847 20927
rect 3789 20887 3847 20893
rect 4338 20884 4344 20936
rect 4396 20884 4402 20936
rect 35526 20884 35532 20936
rect 35584 20924 35590 20936
rect 35693 20927 35751 20933
rect 35693 20924 35705 20927
rect 35584 20896 35705 20924
rect 35584 20884 35590 20896
rect 35693 20893 35705 20896
rect 35739 20893 35751 20927
rect 35693 20887 35751 20893
rect 2317 20859 2375 20865
rect 2317 20825 2329 20859
rect 2363 20856 2375 20859
rect 2590 20856 2596 20868
rect 2363 20828 2596 20856
rect 2363 20825 2375 20828
rect 2317 20819 2375 20825
rect 2590 20816 2596 20828
rect 2648 20816 2654 20868
rect 35345 20859 35403 20865
rect 35345 20825 35357 20859
rect 35391 20856 35403 20859
rect 36446 20856 36452 20868
rect 35391 20828 36452 20856
rect 35391 20825 35403 20828
rect 35345 20819 35403 20825
rect 36446 20816 36452 20828
rect 36504 20816 36510 20868
rect 3510 20748 3516 20800
rect 3568 20748 3574 20800
rect 4522 20748 4528 20800
rect 4580 20748 4586 20800
rect 1104 20698 37812 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 37812 20698
rect 1104 20624 37812 20646
rect 2866 20544 2872 20596
rect 2924 20584 2930 20596
rect 3421 20587 3479 20593
rect 3421 20584 3433 20587
rect 2924 20556 3433 20584
rect 2924 20544 2930 20556
rect 3421 20553 3433 20556
rect 3467 20553 3479 20587
rect 3421 20547 3479 20553
rect 20257 20587 20315 20593
rect 20257 20553 20269 20587
rect 20303 20584 20315 20587
rect 20346 20584 20352 20596
rect 20303 20556 20352 20584
rect 20303 20553 20315 20556
rect 20257 20547 20315 20553
rect 20346 20544 20352 20556
rect 20404 20544 20410 20596
rect 2774 20516 2780 20528
rect 1964 20488 2780 20516
rect 1964 20392 1992 20488
rect 2774 20476 2780 20488
rect 2832 20476 2838 20528
rect 4522 20476 4528 20528
rect 4580 20476 4586 20528
rect 2216 20451 2274 20457
rect 2216 20417 2228 20451
rect 2262 20448 2274 20451
rect 4540 20448 4568 20476
rect 2262 20420 4568 20448
rect 20717 20451 20775 20457
rect 2262 20417 2274 20420
rect 2216 20411 2274 20417
rect 20717 20417 20729 20451
rect 20763 20448 20775 20451
rect 21085 20451 21143 20457
rect 21085 20448 21097 20451
rect 20763 20420 21097 20448
rect 20763 20417 20775 20420
rect 20717 20411 20775 20417
rect 21085 20417 21097 20420
rect 21131 20448 21143 20451
rect 35621 20451 35679 20457
rect 21131 20420 26234 20448
rect 21131 20417 21143 20420
rect 21085 20411 21143 20417
rect 1946 20340 1952 20392
rect 2004 20340 2010 20392
rect 3510 20340 3516 20392
rect 3568 20380 3574 20392
rect 3973 20383 4031 20389
rect 3973 20380 3985 20383
rect 3568 20352 3985 20380
rect 3568 20340 3574 20352
rect 3973 20349 3985 20352
rect 4019 20349 4031 20383
rect 3973 20343 4031 20349
rect 4338 20340 4344 20392
rect 4396 20340 4402 20392
rect 3329 20315 3387 20321
rect 3329 20281 3341 20315
rect 3375 20312 3387 20315
rect 4356 20312 4384 20340
rect 3375 20284 4384 20312
rect 20441 20315 20499 20321
rect 3375 20281 3387 20284
rect 3329 20275 3387 20281
rect 20441 20281 20453 20315
rect 20487 20312 20499 20315
rect 22002 20312 22008 20324
rect 20487 20284 22008 20312
rect 20487 20281 20499 20284
rect 20441 20275 20499 20281
rect 22002 20272 22008 20284
rect 22060 20272 22066 20324
rect 26206 20312 26234 20420
rect 35621 20417 35633 20451
rect 35667 20448 35679 20451
rect 35805 20451 35863 20457
rect 35805 20448 35817 20451
rect 35667 20420 35817 20448
rect 35667 20417 35679 20420
rect 35621 20411 35679 20417
rect 35805 20417 35817 20420
rect 35851 20417 35863 20451
rect 35805 20411 35863 20417
rect 36004 20420 37136 20448
rect 35069 20383 35127 20389
rect 35069 20349 35081 20383
rect 35115 20380 35127 20383
rect 36004 20380 36032 20420
rect 37108 20392 37136 20420
rect 35115 20352 36032 20380
rect 35115 20349 35127 20352
rect 35069 20343 35127 20349
rect 36078 20340 36084 20392
rect 36136 20340 36142 20392
rect 37090 20340 37096 20392
rect 37148 20340 37154 20392
rect 35986 20312 35992 20324
rect 26206 20284 35992 20312
rect 35986 20272 35992 20284
rect 36044 20272 36050 20324
rect 1104 20154 37812 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 37812 20154
rect 1104 20080 37812 20102
rect 25777 20043 25835 20049
rect 25777 20009 25789 20043
rect 25823 20040 25835 20043
rect 28350 20040 28356 20052
rect 25823 20012 28356 20040
rect 25823 20009 25835 20012
rect 25777 20003 25835 20009
rect 28350 20000 28356 20012
rect 28408 20000 28414 20052
rect 35437 20043 35495 20049
rect 35437 20009 35449 20043
rect 35483 20040 35495 20043
rect 35710 20040 35716 20052
rect 35483 20012 35716 20040
rect 35483 20009 35495 20012
rect 35437 20003 35495 20009
rect 934 19864 940 19916
rect 992 19904 998 19916
rect 1581 19907 1639 19913
rect 1581 19904 1593 19907
rect 992 19876 1593 19904
rect 992 19864 998 19876
rect 1581 19873 1593 19876
rect 1627 19873 1639 19907
rect 1581 19867 1639 19873
rect 2961 19907 3019 19913
rect 2961 19873 2973 19907
rect 3007 19904 3019 19907
rect 3050 19904 3056 19916
rect 3007 19876 3056 19904
rect 3007 19873 3019 19876
rect 2961 19867 3019 19873
rect 3050 19864 3056 19876
rect 3108 19864 3114 19916
rect 2590 19796 2596 19848
rect 2648 19796 2654 19848
rect 24394 19796 24400 19848
rect 24452 19836 24458 19848
rect 26053 19839 26111 19845
rect 26053 19836 26065 19839
rect 24452 19808 26065 19836
rect 24452 19796 24458 19808
rect 26053 19805 26065 19808
rect 26099 19805 26111 19839
rect 26053 19799 26111 19805
rect 34606 19796 34612 19848
rect 34664 19836 34670 19848
rect 35544 19845 35572 20012
rect 35710 20000 35716 20012
rect 35768 20000 35774 20052
rect 35805 19907 35863 19913
rect 35805 19873 35817 19907
rect 35851 19904 35863 19907
rect 35986 19904 35992 19916
rect 35851 19876 35992 19904
rect 35851 19873 35863 19876
rect 35805 19867 35863 19873
rect 35986 19864 35992 19876
rect 36044 19864 36050 19916
rect 36078 19864 36084 19916
rect 36136 19864 36142 19916
rect 37185 19907 37243 19913
rect 37185 19873 37197 19907
rect 37231 19904 37243 19907
rect 37274 19904 37280 19916
rect 37231 19876 37280 19904
rect 37231 19873 37243 19876
rect 37185 19867 37243 19873
rect 37274 19864 37280 19876
rect 37332 19864 37338 19916
rect 35529 19839 35587 19845
rect 35529 19836 35541 19839
rect 34664 19808 35541 19836
rect 34664 19796 34670 19808
rect 35529 19805 35541 19808
rect 35575 19805 35587 19839
rect 36096 19836 36124 19864
rect 36173 19839 36231 19845
rect 36173 19836 36185 19839
rect 36096 19808 36185 19836
rect 35529 19799 35587 19805
rect 36173 19805 36185 19808
rect 36219 19805 36231 19839
rect 36173 19799 36231 19805
rect 24670 19777 24676 19780
rect 24664 19731 24676 19777
rect 24670 19728 24676 19731
rect 24728 19728 24734 19780
rect 3234 19660 3240 19712
rect 3292 19700 3298 19712
rect 3513 19703 3571 19709
rect 3513 19700 3525 19703
rect 3292 19672 3525 19700
rect 3292 19660 3298 19672
rect 3513 19669 3525 19672
rect 3559 19669 3571 19703
rect 3513 19663 3571 19669
rect 1104 19610 37812 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 37812 19610
rect 1104 19536 37812 19558
rect 1673 19499 1731 19505
rect 1673 19465 1685 19499
rect 1719 19496 1731 19499
rect 3142 19496 3148 19508
rect 1719 19468 3148 19496
rect 1719 19465 1731 19468
rect 1673 19459 1731 19465
rect 3142 19456 3148 19468
rect 3200 19456 3206 19508
rect 3329 19499 3387 19505
rect 3329 19465 3341 19499
rect 3375 19496 3387 19499
rect 3418 19496 3424 19508
rect 3375 19468 3424 19496
rect 3375 19465 3387 19468
rect 3329 19459 3387 19465
rect 3418 19456 3424 19468
rect 3476 19456 3482 19508
rect 17310 19496 17316 19508
rect 6886 19468 17316 19496
rect 1765 19431 1823 19437
rect 1765 19397 1777 19431
rect 1811 19428 1823 19431
rect 1854 19428 1860 19440
rect 1811 19400 1860 19428
rect 1811 19397 1823 19400
rect 1765 19391 1823 19397
rect 1854 19388 1860 19400
rect 1912 19428 1918 19440
rect 6886 19428 6914 19468
rect 17310 19456 17316 19468
rect 17368 19456 17374 19508
rect 20254 19456 20260 19508
rect 20312 19496 20318 19508
rect 20349 19499 20407 19505
rect 20349 19496 20361 19499
rect 20312 19468 20361 19496
rect 20312 19456 20318 19468
rect 20349 19465 20361 19468
rect 20395 19465 20407 19499
rect 20349 19459 20407 19465
rect 1912 19400 3188 19428
rect 1912 19388 1918 19400
rect 2216 19363 2274 19369
rect 2216 19329 2228 19363
rect 2262 19360 2274 19363
rect 2958 19360 2964 19372
rect 2262 19332 2964 19360
rect 2262 19329 2274 19332
rect 2216 19323 2274 19329
rect 2958 19320 2964 19332
rect 3016 19320 3022 19372
rect 3160 19360 3188 19400
rect 3436 19400 6914 19428
rect 3436 19360 3464 19400
rect 3160 19332 3464 19360
rect 3881 19363 3939 19369
rect 3881 19329 3893 19363
rect 3927 19360 3939 19363
rect 4062 19360 4068 19372
rect 3927 19332 4068 19360
rect 3927 19329 3939 19332
rect 3881 19323 3939 19329
rect 1946 19252 1952 19304
rect 2004 19252 2010 19304
rect 3142 19252 3148 19304
rect 3200 19292 3206 19304
rect 3896 19292 3924 19323
rect 4062 19320 4068 19332
rect 4120 19320 4126 19372
rect 21634 19320 21640 19372
rect 21692 19320 21698 19372
rect 35805 19363 35863 19369
rect 35805 19329 35817 19363
rect 35851 19360 35863 19363
rect 36078 19360 36084 19372
rect 35851 19332 36084 19360
rect 35851 19329 35863 19332
rect 35805 19323 35863 19329
rect 36078 19320 36084 19332
rect 36136 19320 36142 19372
rect 3200 19264 3924 19292
rect 3200 19252 3206 19264
rect 22462 19252 22468 19304
rect 22520 19292 22526 19304
rect 27525 19295 27583 19301
rect 27525 19292 27537 19295
rect 22520 19264 27537 19292
rect 22520 19252 22526 19264
rect 27525 19261 27537 19264
rect 27571 19261 27583 19295
rect 27525 19255 27583 19261
rect 34790 19252 34796 19304
rect 34848 19292 34854 19304
rect 34977 19295 35035 19301
rect 34977 19292 34989 19295
rect 34848 19264 34989 19292
rect 34848 19252 34854 19264
rect 34977 19261 34989 19264
rect 35023 19261 35035 19295
rect 34977 19255 35035 19261
rect 36906 19252 36912 19304
rect 36964 19252 36970 19304
rect 1964 19156 1992 19252
rect 3510 19184 3516 19236
rect 3568 19184 3574 19236
rect 2314 19156 2320 19168
rect 1964 19128 2320 19156
rect 2314 19116 2320 19128
rect 2372 19116 2378 19168
rect 3418 19116 3424 19168
rect 3476 19116 3482 19168
rect 26970 19116 26976 19168
rect 27028 19116 27034 19168
rect 35618 19116 35624 19168
rect 35676 19116 35682 19168
rect 1104 19066 37812 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 37812 19066
rect 1104 18992 37812 19014
rect 1854 18912 1860 18964
rect 1912 18912 1918 18964
rect 35437 18887 35495 18893
rect 35437 18853 35449 18887
rect 35483 18853 35495 18887
rect 35437 18847 35495 18853
rect 3329 18819 3387 18825
rect 3329 18785 3341 18819
rect 3375 18816 3387 18819
rect 35253 18819 35311 18825
rect 3375 18788 4660 18816
rect 3375 18785 3387 18788
rect 3329 18779 3387 18785
rect 2314 18708 2320 18760
rect 2372 18748 2378 18760
rect 3344 18748 3372 18779
rect 4632 18760 4660 18788
rect 35253 18785 35265 18819
rect 35299 18816 35311 18819
rect 35452 18816 35480 18847
rect 37090 18844 37096 18896
rect 37148 18844 37154 18896
rect 35299 18788 35480 18816
rect 35299 18785 35311 18788
rect 35253 18779 35311 18785
rect 2372 18720 3372 18748
rect 2372 18708 2378 18720
rect 3602 18708 3608 18760
rect 3660 18708 3666 18760
rect 4338 18708 4344 18760
rect 4396 18708 4402 18760
rect 4614 18708 4620 18760
rect 4672 18708 4678 18760
rect 35342 18708 35348 18760
rect 35400 18748 35406 18760
rect 36817 18751 36875 18757
rect 36817 18748 36829 18751
rect 35400 18720 36829 18748
rect 35400 18708 35406 18720
rect 36817 18717 36829 18720
rect 36863 18717 36875 18751
rect 36817 18711 36875 18717
rect 3084 18683 3142 18689
rect 3084 18649 3096 18683
rect 3130 18680 3142 18683
rect 3620 18680 3648 18708
rect 3130 18652 3648 18680
rect 36572 18683 36630 18689
rect 3130 18649 3142 18652
rect 3084 18643 3142 18649
rect 36572 18649 36584 18683
rect 36618 18680 36630 18683
rect 36618 18652 36952 18680
rect 36618 18649 36630 18652
rect 36572 18643 36630 18649
rect 1946 18572 1952 18624
rect 2004 18572 2010 18624
rect 3326 18572 3332 18624
rect 3384 18612 3390 18624
rect 3789 18615 3847 18621
rect 3789 18612 3801 18615
rect 3384 18584 3801 18612
rect 3384 18572 3390 18584
rect 3789 18581 3801 18584
rect 3835 18581 3847 18615
rect 3789 18575 3847 18581
rect 34698 18572 34704 18624
rect 34756 18572 34762 18624
rect 36924 18621 36952 18652
rect 36998 18640 37004 18692
rect 37056 18680 37062 18692
rect 37369 18683 37427 18689
rect 37369 18680 37381 18683
rect 37056 18652 37381 18680
rect 37056 18640 37062 18652
rect 37369 18649 37381 18652
rect 37415 18649 37427 18683
rect 37369 18643 37427 18649
rect 36909 18615 36967 18621
rect 36909 18581 36921 18615
rect 36955 18581 36967 18615
rect 36909 18575 36967 18581
rect 1104 18522 37812 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 37812 18522
rect 1104 18448 37812 18470
rect 1946 18368 1952 18420
rect 2004 18368 2010 18420
rect 3605 18411 3663 18417
rect 3605 18377 3617 18411
rect 3651 18408 3663 18411
rect 4338 18408 4344 18420
rect 3651 18380 4344 18408
rect 3651 18377 3663 18380
rect 3605 18371 3663 18377
rect 4338 18368 4344 18380
rect 4396 18368 4402 18420
rect 22462 18368 22468 18420
rect 22520 18368 22526 18420
rect 24118 18368 24124 18420
rect 24176 18368 24182 18420
rect 34698 18368 34704 18420
rect 34756 18368 34762 18420
rect 34790 18368 34796 18420
rect 34848 18408 34854 18420
rect 34977 18411 35035 18417
rect 34977 18408 34989 18411
rect 34848 18380 34989 18408
rect 34848 18368 34854 18380
rect 34977 18377 34989 18380
rect 35023 18377 35035 18411
rect 34977 18371 35035 18377
rect 35986 18368 35992 18420
rect 36044 18408 36050 18420
rect 36725 18411 36783 18417
rect 36725 18408 36737 18411
rect 36044 18380 36737 18408
rect 36044 18368 36050 18380
rect 36725 18377 36737 18380
rect 36771 18408 36783 18411
rect 36998 18408 37004 18420
rect 36771 18380 37004 18408
rect 36771 18377 36783 18380
rect 36725 18371 36783 18377
rect 36998 18368 37004 18380
rect 37056 18368 37062 18420
rect 1581 18275 1639 18281
rect 1581 18241 1593 18275
rect 1627 18272 1639 18275
rect 1964 18272 1992 18368
rect 2492 18343 2550 18349
rect 2492 18309 2504 18343
rect 2538 18340 2550 18343
rect 3418 18340 3424 18352
rect 2538 18312 3424 18340
rect 2538 18309 2550 18312
rect 2492 18303 2550 18309
rect 3418 18300 3424 18312
rect 3476 18300 3482 18352
rect 34333 18343 34391 18349
rect 34333 18309 34345 18343
rect 34379 18340 34391 18343
rect 34425 18343 34483 18349
rect 34425 18340 34437 18343
rect 34379 18312 34437 18340
rect 34379 18309 34391 18312
rect 34333 18303 34391 18309
rect 34425 18309 34437 18312
rect 34471 18340 34483 18343
rect 34606 18340 34612 18352
rect 34471 18312 34612 18340
rect 34471 18309 34483 18312
rect 34425 18303 34483 18309
rect 34606 18300 34612 18312
rect 34664 18300 34670 18352
rect 1627 18244 1992 18272
rect 2225 18275 2283 18281
rect 1627 18241 1639 18244
rect 1581 18235 1639 18241
rect 2225 18241 2237 18275
rect 2271 18272 2283 18275
rect 2314 18272 2320 18284
rect 2271 18244 2320 18272
rect 2271 18241 2283 18244
rect 2225 18235 2283 18241
rect 2314 18232 2320 18244
rect 2372 18232 2378 18284
rect 2958 18232 2964 18284
rect 3016 18272 3022 18284
rect 23937 18275 23995 18281
rect 23937 18272 23949 18275
rect 3016 18244 3280 18272
rect 3016 18232 3022 18244
rect 3252 18204 3280 18244
rect 23492 18244 23949 18272
rect 3697 18207 3755 18213
rect 3697 18204 3709 18207
rect 3252 18176 3709 18204
rect 3697 18173 3709 18176
rect 3743 18173 3755 18207
rect 3697 18167 3755 18173
rect 4157 18207 4215 18213
rect 4157 18173 4169 18207
rect 4203 18173 4215 18207
rect 4157 18167 4215 18173
rect 3786 18096 3792 18148
rect 3844 18096 3850 18148
rect 2133 18071 2191 18077
rect 2133 18037 2145 18071
rect 2179 18068 2191 18071
rect 2958 18068 2964 18080
rect 2179 18040 2964 18068
rect 2179 18037 2191 18040
rect 2133 18031 2191 18037
rect 2958 18028 2964 18040
rect 3016 18028 3022 18080
rect 4172 18068 4200 18167
rect 21818 18164 21824 18216
rect 21876 18164 21882 18216
rect 23492 18148 23520 18244
rect 23937 18241 23949 18244
rect 23983 18272 23995 18275
rect 26970 18272 26976 18284
rect 23983 18244 26976 18272
rect 23983 18241 23995 18244
rect 23937 18235 23995 18241
rect 26970 18232 26976 18244
rect 27028 18232 27034 18284
rect 34716 18272 34744 18368
rect 36078 18300 36084 18352
rect 36136 18340 36142 18352
rect 36173 18343 36231 18349
rect 36173 18340 36185 18343
rect 36136 18312 36185 18340
rect 36136 18300 36142 18312
rect 36173 18309 36185 18312
rect 36219 18309 36231 18343
rect 36173 18303 36231 18309
rect 35529 18275 35587 18281
rect 35529 18272 35541 18275
rect 34716 18244 35541 18272
rect 35529 18241 35541 18244
rect 35575 18241 35587 18275
rect 35529 18235 35587 18241
rect 35618 18232 35624 18284
rect 35676 18272 35682 18284
rect 35805 18275 35863 18281
rect 35805 18272 35817 18275
rect 35676 18244 35817 18272
rect 35676 18232 35682 18244
rect 35805 18241 35817 18244
rect 35851 18241 35863 18275
rect 35805 18235 35863 18241
rect 34790 18164 34796 18216
rect 34848 18164 34854 18216
rect 23474 18096 23480 18148
rect 23532 18096 23538 18148
rect 34701 18139 34759 18145
rect 34701 18105 34713 18139
rect 34747 18136 34759 18139
rect 34808 18136 34836 18164
rect 34747 18108 34836 18136
rect 34747 18105 34759 18108
rect 34701 18099 34759 18105
rect 4525 18071 4583 18077
rect 4525 18068 4537 18071
rect 4172 18040 4537 18068
rect 4525 18037 4537 18040
rect 4571 18068 4583 18071
rect 4706 18068 4712 18080
rect 4571 18040 4712 18068
rect 4571 18037 4583 18040
rect 4525 18031 4583 18037
rect 4706 18028 4712 18040
rect 4764 18028 4770 18080
rect 34885 18071 34943 18077
rect 34885 18037 34897 18071
rect 34931 18068 34943 18071
rect 35526 18068 35532 18080
rect 34931 18040 35532 18068
rect 34931 18037 34943 18040
rect 34885 18031 34943 18037
rect 35526 18028 35532 18040
rect 35584 18028 35590 18080
rect 1104 17978 37812 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 37812 17978
rect 1104 17904 37812 17926
rect 27522 17824 27528 17876
rect 27580 17824 27586 17876
rect 3513 17799 3571 17805
rect 3513 17765 3525 17799
rect 3559 17796 3571 17799
rect 27433 17799 27491 17805
rect 3559 17768 6914 17796
rect 3559 17765 3571 17768
rect 3513 17759 3571 17765
rect 1578 17688 1584 17740
rect 1636 17688 1642 17740
rect 2958 17688 2964 17740
rect 3016 17728 3022 17740
rect 3789 17731 3847 17737
rect 3789 17728 3801 17731
rect 3016 17700 3801 17728
rect 3016 17688 3022 17700
rect 3789 17697 3801 17700
rect 3835 17697 3847 17731
rect 3789 17691 3847 17697
rect 2590 17620 2596 17672
rect 2648 17620 2654 17672
rect 2869 17663 2927 17669
rect 2869 17629 2881 17663
rect 2915 17660 2927 17663
rect 3326 17660 3332 17672
rect 2915 17632 3332 17660
rect 2915 17629 2927 17632
rect 2869 17623 2927 17629
rect 3326 17620 3332 17632
rect 3384 17620 3390 17672
rect 6886 17660 6914 17768
rect 27433 17765 27445 17799
rect 27479 17796 27491 17799
rect 27890 17796 27896 17808
rect 27479 17768 27896 17796
rect 27479 17765 27491 17768
rect 27433 17759 27491 17765
rect 27890 17756 27896 17768
rect 27948 17756 27954 17808
rect 8205 17663 8263 17669
rect 8205 17660 8217 17663
rect 6886 17632 8217 17660
rect 8205 17629 8217 17632
rect 8251 17660 8263 17663
rect 11882 17660 11888 17672
rect 8251 17632 11888 17660
rect 8251 17629 8263 17632
rect 8205 17623 8263 17629
rect 11882 17620 11888 17632
rect 11940 17620 11946 17672
rect 33965 17663 34023 17669
rect 33965 17629 33977 17663
rect 34011 17660 34023 17663
rect 34011 17632 34744 17660
rect 34011 17629 34023 17632
rect 33965 17623 34023 17629
rect 27065 17595 27123 17601
rect 27065 17561 27077 17595
rect 27111 17561 27123 17595
rect 27065 17555 27123 17561
rect 3878 17484 3884 17536
rect 3936 17524 3942 17536
rect 4433 17527 4491 17533
rect 4433 17524 4445 17527
rect 3936 17496 4445 17524
rect 3936 17484 3942 17496
rect 4433 17493 4445 17496
rect 4479 17493 4491 17527
rect 4433 17487 4491 17493
rect 7558 17484 7564 17536
rect 7616 17484 7622 17536
rect 21910 17484 21916 17536
rect 21968 17524 21974 17536
rect 27080 17524 27108 17555
rect 34716 17536 34744 17632
rect 35250 17620 35256 17672
rect 35308 17620 35314 17672
rect 35342 17620 35348 17672
rect 35400 17660 35406 17672
rect 35437 17663 35495 17669
rect 35437 17660 35449 17663
rect 35400 17632 35449 17660
rect 35400 17620 35406 17632
rect 35437 17629 35449 17632
rect 35483 17629 35495 17663
rect 35437 17623 35495 17629
rect 35526 17620 35532 17672
rect 35584 17660 35590 17672
rect 35693 17663 35751 17669
rect 35693 17660 35705 17663
rect 35584 17632 35705 17660
rect 35584 17620 35590 17632
rect 35693 17629 35705 17632
rect 35739 17629 35751 17663
rect 35693 17623 35751 17629
rect 27893 17527 27951 17533
rect 27893 17524 27905 17527
rect 21968 17496 27905 17524
rect 21968 17484 21974 17496
rect 27893 17493 27905 17496
rect 27939 17524 27951 17527
rect 30190 17524 30196 17536
rect 27939 17496 30196 17524
rect 27939 17493 27951 17496
rect 27893 17487 27951 17493
rect 30190 17484 30196 17496
rect 30248 17484 30254 17536
rect 34514 17484 34520 17536
rect 34572 17484 34578 17536
rect 34698 17484 34704 17536
rect 34756 17484 34762 17536
rect 36814 17484 36820 17536
rect 36872 17484 36878 17536
rect 1104 17434 37812 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 37812 17434
rect 1104 17360 37812 17382
rect 2590 17320 2596 17332
rect 2332 17292 2596 17320
rect 2332 17261 2360 17292
rect 2590 17280 2596 17292
rect 2648 17280 2654 17332
rect 7558 17320 7564 17332
rect 2700 17292 7564 17320
rect 2317 17255 2375 17261
rect 2317 17221 2329 17255
rect 2363 17221 2375 17255
rect 2317 17215 2375 17221
rect 2700 17193 2728 17292
rect 7558 17280 7564 17292
rect 7616 17280 7622 17332
rect 34514 17280 34520 17332
rect 34572 17280 34578 17332
rect 34977 17323 35035 17329
rect 34977 17289 34989 17323
rect 35023 17320 35035 17323
rect 35250 17320 35256 17332
rect 35023 17292 35256 17320
rect 35023 17289 35035 17292
rect 34977 17283 35035 17289
rect 35250 17280 35256 17292
rect 35308 17280 35314 17332
rect 36814 17280 36820 17332
rect 36872 17280 36878 17332
rect 2685 17187 2743 17193
rect 2685 17153 2697 17187
rect 2731 17153 2743 17187
rect 2685 17147 2743 17153
rect 3694 17144 3700 17196
rect 3752 17184 3758 17196
rect 3982 17187 4040 17193
rect 3982 17184 3994 17187
rect 3752 17156 3994 17184
rect 3752 17144 3758 17156
rect 3982 17153 3994 17156
rect 4028 17153 4040 17187
rect 3982 17147 4040 17153
rect 4249 17187 4307 17193
rect 4249 17153 4261 17187
rect 4295 17184 4307 17187
rect 4614 17184 4620 17196
rect 4295 17156 4620 17184
rect 4295 17153 4307 17156
rect 4249 17147 4307 17153
rect 4614 17144 4620 17156
rect 4672 17144 4678 17196
rect 34532 17184 34560 17280
rect 35805 17187 35863 17193
rect 35805 17184 35817 17187
rect 34532 17156 35817 17184
rect 35805 17153 35817 17156
rect 35851 17153 35863 17187
rect 36832 17184 36860 17280
rect 35805 17147 35863 17153
rect 36096 17156 36860 17184
rect 4890 17076 4896 17128
rect 4948 17076 4954 17128
rect 35621 17119 35679 17125
rect 35621 17085 35633 17119
rect 35667 17116 35679 17119
rect 36096 17116 36124 17156
rect 35667 17088 36124 17116
rect 35667 17085 35679 17088
rect 35621 17079 35679 17085
rect 36262 17076 36268 17128
rect 36320 17076 36326 17128
rect 2866 16940 2872 16992
rect 2924 16940 2930 16992
rect 4341 16983 4399 16989
rect 4341 16949 4353 16983
rect 4387 16980 4399 16983
rect 4614 16980 4620 16992
rect 4387 16952 4620 16980
rect 4387 16949 4399 16952
rect 4341 16943 4399 16949
rect 4614 16940 4620 16952
rect 4672 16940 4678 16992
rect 20898 16940 20904 16992
rect 20956 16940 20962 16992
rect 1104 16890 37812 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 37812 16890
rect 1104 16816 37812 16838
rect 2866 16736 2872 16788
rect 2924 16776 2930 16788
rect 23474 16776 23480 16788
rect 2924 16748 3464 16776
rect 2924 16736 2930 16748
rect 3436 16649 3464 16748
rect 20548 16748 23480 16776
rect 20548 16717 20576 16748
rect 23474 16736 23480 16748
rect 23532 16736 23538 16788
rect 34517 16779 34575 16785
rect 34517 16745 34529 16779
rect 34563 16776 34575 16779
rect 34606 16776 34612 16788
rect 34563 16748 34612 16776
rect 34563 16745 34575 16748
rect 34517 16739 34575 16745
rect 34606 16736 34612 16748
rect 34664 16736 34670 16788
rect 20533 16711 20591 16717
rect 20533 16677 20545 16711
rect 20579 16677 20591 16711
rect 20533 16671 20591 16677
rect 20898 16668 20904 16720
rect 20956 16708 20962 16720
rect 21361 16711 21419 16717
rect 21361 16708 21373 16711
rect 20956 16680 21373 16708
rect 20956 16668 20962 16680
rect 21361 16677 21373 16680
rect 21407 16677 21419 16711
rect 21361 16671 21419 16677
rect 21450 16668 21456 16720
rect 21508 16708 21514 16720
rect 21910 16708 21916 16720
rect 21508 16680 21916 16708
rect 21508 16668 21514 16680
rect 21910 16668 21916 16680
rect 21968 16668 21974 16720
rect 3421 16643 3479 16649
rect 3421 16609 3433 16643
rect 3467 16609 3479 16643
rect 3421 16603 3479 16609
rect 3510 16600 3516 16652
rect 3568 16640 3574 16652
rect 4709 16643 4767 16649
rect 4709 16640 4721 16643
rect 3568 16612 4721 16640
rect 3568 16600 3574 16612
rect 4709 16609 4721 16612
rect 4755 16609 4767 16643
rect 4709 16603 4767 16609
rect 14274 16600 14280 16652
rect 14332 16640 14338 16652
rect 15473 16643 15531 16649
rect 15473 16640 15485 16643
rect 14332 16612 15485 16640
rect 14332 16600 14338 16612
rect 15473 16609 15485 16612
rect 15519 16609 15531 16643
rect 15473 16603 15531 16609
rect 20257 16643 20315 16649
rect 20257 16609 20269 16643
rect 20303 16640 20315 16643
rect 20809 16643 20867 16649
rect 20809 16640 20821 16643
rect 20303 16612 20821 16640
rect 20303 16609 20315 16612
rect 20257 16603 20315 16609
rect 20809 16609 20821 16612
rect 20855 16640 20867 16643
rect 21085 16643 21143 16649
rect 21085 16640 21097 16643
rect 20855 16612 21097 16640
rect 20855 16609 20867 16612
rect 20809 16603 20867 16609
rect 21085 16609 21097 16612
rect 21131 16640 21143 16643
rect 21468 16640 21496 16668
rect 21131 16612 21496 16640
rect 34624 16640 34652 16736
rect 34698 16668 34704 16720
rect 34756 16708 34762 16720
rect 35069 16711 35127 16717
rect 35069 16708 35081 16711
rect 34756 16680 35081 16708
rect 34756 16668 34762 16680
rect 35069 16677 35081 16680
rect 35115 16677 35127 16711
rect 35069 16671 35127 16677
rect 34793 16643 34851 16649
rect 34793 16640 34805 16643
rect 34624 16612 34805 16640
rect 21131 16609 21143 16612
rect 21085 16603 21143 16609
rect 34793 16609 34805 16612
rect 34839 16609 34851 16643
rect 34793 16603 34851 16609
rect 37182 16600 37188 16652
rect 37240 16600 37246 16652
rect 1578 16532 1584 16584
rect 1636 16532 1642 16584
rect 2590 16532 2596 16584
rect 2648 16532 2654 16584
rect 3878 16532 3884 16584
rect 3936 16572 3942 16584
rect 4341 16575 4399 16581
rect 4341 16572 4353 16575
rect 3936 16544 4353 16572
rect 3936 16532 3942 16544
rect 4341 16541 4353 16544
rect 4387 16541 4399 16575
rect 24670 16572 24676 16584
rect 4341 16535 4399 16541
rect 21652 16544 24676 16572
rect 4246 16464 4252 16516
rect 4304 16504 4310 16516
rect 4954 16507 5012 16513
rect 4954 16504 4966 16507
rect 4304 16476 4966 16504
rect 4304 16464 4310 16476
rect 4954 16473 4966 16476
rect 5000 16473 5012 16507
rect 4954 16467 5012 16473
rect 13262 16464 13268 16516
rect 13320 16504 13326 16516
rect 15718 16507 15776 16513
rect 15718 16504 15730 16507
rect 13320 16476 15730 16504
rect 13320 16464 13326 16476
rect 15718 16473 15730 16476
rect 15764 16473 15776 16507
rect 15718 16467 15776 16473
rect 16868 16476 20760 16504
rect 2866 16396 2872 16448
rect 2924 16396 2930 16448
rect 3234 16396 3240 16448
rect 3292 16436 3298 16448
rect 3789 16439 3847 16445
rect 3789 16436 3801 16439
rect 3292 16408 3801 16436
rect 3292 16396 3298 16408
rect 3789 16405 3801 16408
rect 3835 16405 3847 16439
rect 3789 16399 3847 16405
rect 6089 16439 6147 16445
rect 6089 16405 6101 16439
rect 6135 16436 6147 16439
rect 6546 16436 6552 16448
rect 6135 16408 6552 16436
rect 6135 16405 6147 16408
rect 6089 16399 6147 16405
rect 6546 16396 6552 16408
rect 6604 16396 6610 16448
rect 16868 16445 16896 16476
rect 20732 16448 20760 16476
rect 16853 16439 16911 16445
rect 16853 16405 16865 16439
rect 16899 16405 16911 16439
rect 16853 16399 16911 16405
rect 20349 16439 20407 16445
rect 20349 16405 20361 16439
rect 20395 16436 20407 16439
rect 20438 16436 20444 16448
rect 20395 16408 20444 16436
rect 20395 16405 20407 16408
rect 20349 16399 20407 16405
rect 20438 16396 20444 16408
rect 20496 16396 20502 16448
rect 20714 16396 20720 16448
rect 20772 16396 20778 16448
rect 21545 16439 21603 16445
rect 21545 16405 21557 16439
rect 21591 16436 21603 16439
rect 21652 16436 21680 16544
rect 24670 16532 24676 16544
rect 24728 16532 24734 16584
rect 35986 16532 35992 16584
rect 36044 16532 36050 16584
rect 36262 16532 36268 16584
rect 36320 16532 36326 16584
rect 35268 16476 35572 16504
rect 21591 16408 21680 16436
rect 21591 16405 21603 16408
rect 21545 16399 21603 16405
rect 22278 16396 22284 16448
rect 22336 16436 22342 16448
rect 24394 16436 24400 16448
rect 22336 16408 24400 16436
rect 22336 16396 22342 16408
rect 24394 16396 24400 16408
rect 24452 16396 24458 16448
rect 35268 16445 35296 16476
rect 35544 16448 35572 16476
rect 35253 16439 35311 16445
rect 35253 16405 35265 16439
rect 35299 16405 35311 16439
rect 35253 16399 35311 16405
rect 35345 16439 35403 16445
rect 35345 16405 35357 16439
rect 35391 16436 35403 16439
rect 35434 16436 35440 16448
rect 35391 16408 35440 16436
rect 35391 16405 35403 16408
rect 35345 16399 35403 16405
rect 35434 16396 35440 16408
rect 35492 16396 35498 16448
rect 35526 16396 35532 16448
rect 35584 16396 35590 16448
rect 1104 16346 37812 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 37812 16346
rect 1104 16272 37812 16294
rect 2590 16232 2596 16244
rect 2332 16204 2596 16232
rect 2332 16173 2360 16204
rect 2590 16192 2596 16204
rect 2648 16192 2654 16244
rect 2866 16192 2872 16244
rect 2924 16192 2930 16244
rect 4246 16192 4252 16244
rect 4304 16192 4310 16244
rect 13262 16192 13268 16244
rect 13320 16192 13326 16244
rect 13633 16235 13691 16241
rect 13633 16201 13645 16235
rect 13679 16232 13691 16235
rect 16114 16232 16120 16244
rect 13679 16204 16120 16232
rect 13679 16201 13691 16204
rect 13633 16195 13691 16201
rect 2317 16167 2375 16173
rect 2317 16133 2329 16167
rect 2363 16133 2375 16167
rect 2317 16127 2375 16133
rect 2884 16105 2912 16192
rect 3789 16167 3847 16173
rect 3789 16133 3801 16167
rect 3835 16164 3847 16167
rect 4062 16164 4068 16176
rect 3835 16136 4068 16164
rect 3835 16133 3847 16136
rect 3789 16127 3847 16133
rect 4062 16124 4068 16136
rect 4120 16164 4126 16176
rect 4525 16167 4583 16173
rect 4525 16164 4537 16167
rect 4120 16136 4537 16164
rect 4120 16124 4126 16136
rect 4525 16133 4537 16136
rect 4571 16164 4583 16167
rect 4706 16164 4712 16176
rect 4571 16136 4712 16164
rect 4571 16133 4583 16136
rect 4525 16127 4583 16133
rect 4706 16124 4712 16136
rect 4764 16124 4770 16176
rect 12802 16124 12808 16176
rect 12860 16164 12866 16176
rect 13648 16164 13676 16195
rect 16114 16192 16120 16204
rect 16172 16232 16178 16244
rect 17862 16232 17868 16244
rect 16172 16204 17868 16232
rect 16172 16192 16178 16204
rect 17862 16192 17868 16204
rect 17920 16192 17926 16244
rect 20714 16192 20720 16244
rect 20772 16232 20778 16244
rect 21818 16232 21824 16244
rect 20772 16204 21824 16232
rect 20772 16192 20778 16204
rect 21818 16192 21824 16204
rect 21876 16192 21882 16244
rect 22278 16192 22284 16244
rect 22336 16192 22342 16244
rect 35434 16192 35440 16244
rect 35492 16192 35498 16244
rect 35986 16192 35992 16244
rect 36044 16232 36050 16244
rect 36817 16235 36875 16241
rect 36817 16232 36829 16235
rect 36044 16204 36829 16232
rect 36044 16192 36050 16204
rect 36817 16201 36829 16204
rect 36863 16201 36875 16235
rect 36817 16195 36875 16201
rect 22296 16164 22324 16192
rect 35452 16164 35480 16192
rect 12860 16136 13676 16164
rect 20180 16136 22324 16164
rect 35268 16136 35480 16164
rect 12860 16124 12866 16136
rect 2685 16099 2743 16105
rect 2685 16065 2697 16099
rect 2731 16065 2743 16099
rect 2685 16059 2743 16065
rect 2869 16099 2927 16105
rect 2869 16065 2881 16099
rect 2915 16065 2927 16099
rect 4614 16096 4620 16108
rect 2869 16059 2927 16065
rect 3712 16068 4620 16096
rect 2700 16028 2728 16059
rect 3712 16028 3740 16068
rect 4614 16056 4620 16068
rect 4672 16056 4678 16108
rect 20180 16105 20208 16136
rect 20438 16105 20444 16108
rect 20165 16099 20223 16105
rect 20165 16065 20177 16099
rect 20211 16065 20223 16099
rect 20165 16059 20223 16065
rect 20432 16059 20444 16105
rect 20438 16056 20444 16059
rect 20496 16056 20502 16108
rect 21836 16105 21864 16136
rect 21821 16099 21879 16105
rect 21821 16065 21833 16099
rect 21867 16065 21879 16099
rect 21821 16059 21879 16065
rect 21910 16056 21916 16108
rect 21968 16096 21974 16108
rect 35268 16105 35296 16136
rect 35526 16124 35532 16176
rect 35584 16164 35590 16176
rect 35682 16167 35740 16173
rect 35682 16164 35694 16167
rect 35584 16136 35694 16164
rect 35584 16124 35590 16136
rect 35682 16133 35694 16136
rect 35728 16133 35740 16167
rect 35682 16127 35740 16133
rect 22077 16099 22135 16105
rect 22077 16096 22089 16099
rect 21968 16068 22089 16096
rect 21968 16056 21974 16068
rect 22077 16065 22089 16068
rect 22123 16065 22135 16099
rect 22077 16059 22135 16065
rect 35253 16099 35311 16105
rect 35253 16065 35265 16099
rect 35299 16065 35311 16099
rect 35253 16059 35311 16065
rect 35342 16056 35348 16108
rect 35400 16096 35406 16108
rect 35437 16099 35495 16105
rect 35437 16096 35449 16099
rect 35400 16068 35449 16096
rect 35400 16056 35406 16068
rect 35437 16065 35449 16068
rect 35483 16065 35495 16099
rect 35437 16059 35495 16065
rect 2700 16000 3740 16028
rect 3513 15963 3571 15969
rect 3513 15929 3525 15963
rect 3559 15960 3571 15963
rect 4065 15963 4123 15969
rect 4065 15960 4077 15963
rect 3559 15932 4077 15960
rect 3559 15929 3571 15932
rect 3513 15923 3571 15929
rect 4065 15929 4077 15932
rect 4111 15960 4123 15963
rect 4890 15960 4896 15972
rect 4111 15932 4896 15960
rect 4111 15929 4123 15932
rect 4065 15923 4123 15929
rect 4890 15920 4896 15932
rect 4948 15920 4954 15972
rect 13078 15920 13084 15972
rect 13136 15920 13142 15972
rect 25314 15960 25320 15972
rect 23124 15932 25320 15960
rect 21545 15895 21603 15901
rect 21545 15861 21557 15895
rect 21591 15892 21603 15895
rect 23124 15892 23152 15932
rect 25314 15920 25320 15932
rect 25372 15920 25378 15972
rect 21591 15864 23152 15892
rect 21591 15861 21603 15864
rect 21545 15855 21603 15861
rect 23198 15852 23204 15904
rect 23256 15852 23262 15904
rect 23569 15895 23627 15901
rect 23569 15861 23581 15895
rect 23615 15892 23627 15895
rect 24394 15892 24400 15904
rect 23615 15864 24400 15892
rect 23615 15861 23627 15864
rect 23569 15855 23627 15861
rect 24394 15852 24400 15864
rect 24452 15852 24458 15904
rect 34698 15852 34704 15904
rect 34756 15852 34762 15904
rect 1104 15802 37812 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 37812 15802
rect 1104 15728 37812 15750
rect 3234 15688 3240 15700
rect 2700 15660 3240 15688
rect 2700 15493 2728 15660
rect 3234 15648 3240 15660
rect 3292 15648 3298 15700
rect 3329 15691 3387 15697
rect 3329 15657 3341 15691
rect 3375 15688 3387 15691
rect 3694 15688 3700 15700
rect 3375 15660 3700 15688
rect 3375 15657 3387 15660
rect 3329 15651 3387 15657
rect 3694 15648 3700 15660
rect 3752 15648 3758 15700
rect 12621 15691 12679 15697
rect 12621 15657 12633 15691
rect 12667 15688 12679 15691
rect 12802 15688 12808 15700
rect 12667 15660 12808 15688
rect 12667 15657 12679 15660
rect 12621 15651 12679 15657
rect 2866 15580 2872 15632
rect 2924 15620 2930 15632
rect 3145 15623 3203 15629
rect 3145 15620 3157 15623
rect 2924 15592 3157 15620
rect 2924 15580 2930 15592
rect 3145 15589 3157 15592
rect 3191 15589 3203 15623
rect 3145 15583 3203 15589
rect 3160 15552 3188 15583
rect 11882 15580 11888 15632
rect 11940 15580 11946 15632
rect 3160 15524 4476 15552
rect 4448 15493 4476 15524
rect 2685 15487 2743 15493
rect 2685 15453 2697 15487
rect 2731 15453 2743 15487
rect 4433 15487 4491 15493
rect 2685 15447 2743 15453
rect 2792 15456 4292 15484
rect 2317 15419 2375 15425
rect 2317 15385 2329 15419
rect 2363 15416 2375 15419
rect 2590 15416 2596 15428
rect 2363 15388 2596 15416
rect 2363 15385 2375 15388
rect 2317 15379 2375 15385
rect 2590 15376 2596 15388
rect 2648 15376 2654 15428
rect 2682 15308 2688 15360
rect 2740 15348 2746 15360
rect 2792 15348 2820 15456
rect 2869 15419 2927 15425
rect 2869 15385 2881 15419
rect 2915 15416 2927 15419
rect 2915 15388 3096 15416
rect 2915 15385 2927 15388
rect 2869 15379 2927 15385
rect 2740 15320 2820 15348
rect 3068 15348 3096 15388
rect 4062 15348 4068 15360
rect 3068 15320 4068 15348
rect 2740 15308 2746 15320
rect 4062 15308 4068 15320
rect 4120 15308 4126 15360
rect 4264 15357 4292 15456
rect 4433 15453 4445 15487
rect 4479 15453 4491 15487
rect 4433 15447 4491 15453
rect 12253 15487 12311 15493
rect 12253 15453 12265 15487
rect 12299 15484 12311 15487
rect 12636 15484 12664 15651
rect 12802 15648 12808 15660
rect 12860 15648 12866 15700
rect 21910 15648 21916 15700
rect 21968 15648 21974 15700
rect 21821 15623 21879 15629
rect 21821 15589 21833 15623
rect 21867 15620 21879 15623
rect 24854 15620 24860 15632
rect 21867 15592 24860 15620
rect 21867 15589 21879 15592
rect 21821 15583 21879 15589
rect 24854 15580 24860 15592
rect 24912 15580 24918 15632
rect 21450 15512 21456 15564
rect 21508 15512 21514 15564
rect 34698 15512 34704 15564
rect 34756 15552 34762 15564
rect 35345 15555 35403 15561
rect 35345 15552 35357 15555
rect 34756 15524 35357 15552
rect 34756 15512 34762 15524
rect 35345 15521 35357 15524
rect 35391 15521 35403 15555
rect 35345 15515 35403 15521
rect 12299 15456 12664 15484
rect 12299 15453 12311 15456
rect 12253 15447 12311 15453
rect 22002 15444 22008 15496
rect 22060 15484 22066 15496
rect 22922 15484 22928 15496
rect 22060 15456 22928 15484
rect 22060 15444 22066 15456
rect 22922 15444 22928 15456
rect 22980 15444 22986 15496
rect 35989 15487 36047 15493
rect 35989 15453 36001 15487
rect 36035 15484 36047 15487
rect 36173 15487 36231 15493
rect 36173 15484 36185 15487
rect 36035 15456 36185 15484
rect 36035 15453 36047 15456
rect 35989 15447 36047 15453
rect 36173 15453 36185 15456
rect 36219 15453 36231 15487
rect 36173 15447 36231 15453
rect 36538 15376 36544 15428
rect 36596 15376 36602 15428
rect 4249 15351 4307 15357
rect 4249 15317 4261 15351
rect 4295 15317 4307 15351
rect 4249 15311 4307 15317
rect 11793 15351 11851 15357
rect 11793 15317 11805 15351
rect 11839 15348 11851 15351
rect 13814 15348 13820 15360
rect 11839 15320 13820 15348
rect 11839 15317 11851 15320
rect 11793 15311 11851 15317
rect 13814 15308 13820 15320
rect 13872 15308 13878 15360
rect 22649 15351 22707 15357
rect 22649 15317 22661 15351
rect 22695 15348 22707 15351
rect 23382 15348 23388 15360
rect 22695 15320 23388 15348
rect 22695 15317 22707 15320
rect 22649 15311 22707 15317
rect 23382 15308 23388 15320
rect 23440 15308 23446 15360
rect 34514 15308 34520 15360
rect 34572 15348 34578 15360
rect 34977 15351 35035 15357
rect 34977 15348 34989 15351
rect 34572 15320 34989 15348
rect 34572 15308 34578 15320
rect 34977 15317 34989 15320
rect 35023 15317 35035 15351
rect 34977 15311 35035 15317
rect 1104 15258 37812 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 37812 15258
rect 1104 15184 37812 15206
rect 21450 15104 21456 15156
rect 21508 15144 21514 15156
rect 22097 15147 22155 15153
rect 22097 15144 22109 15147
rect 21508 15116 22109 15144
rect 21508 15104 21514 15116
rect 22097 15113 22109 15116
rect 22143 15113 22155 15147
rect 22097 15107 22155 15113
rect 1578 15036 1584 15088
rect 1636 15036 1642 15088
rect 36906 15036 36912 15088
rect 36964 15036 36970 15088
rect 2590 14968 2596 15020
rect 2648 14968 2654 15020
rect 35805 15011 35863 15017
rect 35805 14977 35817 15011
rect 35851 15008 35863 15011
rect 36538 15008 36544 15020
rect 35851 14980 36544 15008
rect 35851 14977 35863 14980
rect 35805 14971 35863 14977
rect 36538 14968 36544 14980
rect 36596 14968 36602 15020
rect 1946 14900 1952 14952
rect 2004 14940 2010 14952
rect 2869 14943 2927 14949
rect 2869 14940 2881 14943
rect 2004 14912 2881 14940
rect 2004 14900 2010 14912
rect 2869 14909 2881 14912
rect 2915 14909 2927 14943
rect 2869 14903 2927 14909
rect 3513 14943 3571 14949
rect 3513 14909 3525 14943
rect 3559 14940 3571 14943
rect 3970 14940 3976 14952
rect 3559 14912 3976 14940
rect 3559 14909 3571 14912
rect 3513 14903 3571 14909
rect 3970 14900 3976 14912
rect 4028 14900 4034 14952
rect 4065 14943 4123 14949
rect 4065 14909 4077 14943
rect 4111 14909 4123 14943
rect 4065 14903 4123 14909
rect 3789 14875 3847 14881
rect 3789 14841 3801 14875
rect 3835 14872 3847 14875
rect 3878 14872 3884 14884
rect 3835 14844 3884 14872
rect 3835 14841 3847 14844
rect 3789 14835 3847 14841
rect 3878 14832 3884 14844
rect 3936 14832 3942 14884
rect 4080 14816 4108 14903
rect 34422 14900 34428 14952
rect 34480 14900 34486 14952
rect 35069 14943 35127 14949
rect 35069 14909 35081 14943
rect 35115 14940 35127 14943
rect 35434 14940 35440 14952
rect 35115 14912 35440 14940
rect 35115 14909 35127 14912
rect 35069 14903 35127 14909
rect 35434 14900 35440 14912
rect 35492 14900 35498 14952
rect 34698 14832 34704 14884
rect 34756 14832 34762 14884
rect 3602 14764 3608 14816
rect 3660 14764 3666 14816
rect 4062 14764 4068 14816
rect 4120 14804 4126 14816
rect 4341 14807 4399 14813
rect 4341 14804 4353 14807
rect 4120 14776 4353 14804
rect 4120 14764 4126 14776
rect 4341 14773 4353 14776
rect 4387 14773 4399 14807
rect 4341 14767 4399 14773
rect 34885 14807 34943 14813
rect 34885 14773 34897 14807
rect 34931 14804 34943 14807
rect 35526 14804 35532 14816
rect 34931 14776 35532 14804
rect 34931 14773 34943 14776
rect 34885 14767 34943 14773
rect 35526 14764 35532 14776
rect 35584 14764 35590 14816
rect 35621 14807 35679 14813
rect 35621 14773 35633 14807
rect 35667 14804 35679 14807
rect 35710 14804 35716 14816
rect 35667 14776 35716 14804
rect 35667 14773 35679 14776
rect 35621 14767 35679 14773
rect 35710 14764 35716 14776
rect 35768 14764 35774 14816
rect 1104 14714 37812 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 37812 14714
rect 1104 14640 37812 14662
rect 1946 14560 1952 14612
rect 2004 14560 2010 14612
rect 3602 14560 3608 14612
rect 3660 14560 3666 14612
rect 3970 14560 3976 14612
rect 4028 14560 4034 14612
rect 35345 14603 35403 14609
rect 35345 14569 35357 14603
rect 35391 14600 35403 14603
rect 35434 14600 35440 14612
rect 35391 14572 35440 14600
rect 35391 14569 35403 14572
rect 35345 14563 35403 14569
rect 35434 14560 35440 14572
rect 35492 14560 35498 14612
rect 3329 14467 3387 14473
rect 3329 14433 3341 14467
rect 3375 14464 3387 14467
rect 3510 14464 3516 14476
rect 3375 14436 3516 14464
rect 3375 14433 3387 14436
rect 3329 14427 3387 14433
rect 3510 14424 3516 14436
rect 3568 14424 3574 14476
rect 3073 14399 3131 14405
rect 3073 14365 3085 14399
rect 3119 14396 3131 14399
rect 3620 14396 3648 14560
rect 3988 14464 4016 14560
rect 4341 14467 4399 14473
rect 4341 14464 4353 14467
rect 3988 14436 4353 14464
rect 4341 14433 4353 14436
rect 4387 14433 4399 14467
rect 4341 14427 4399 14433
rect 35342 14424 35348 14476
rect 35400 14464 35406 14476
rect 35437 14467 35495 14473
rect 35437 14464 35449 14467
rect 35400 14436 35449 14464
rect 35400 14424 35406 14436
rect 35437 14433 35449 14436
rect 35483 14433 35495 14467
rect 35437 14427 35495 14433
rect 3119 14368 3648 14396
rect 3119 14365 3131 14368
rect 3073 14359 3131 14365
rect 34790 14356 34796 14408
rect 34848 14356 34854 14408
rect 35526 14356 35532 14408
rect 35584 14396 35590 14408
rect 35693 14399 35751 14405
rect 35693 14396 35705 14399
rect 35584 14368 35705 14396
rect 35584 14356 35590 14368
rect 35693 14365 35705 14368
rect 35739 14365 35751 14399
rect 35693 14359 35751 14365
rect 3786 14220 3792 14272
rect 3844 14220 3850 14272
rect 35802 14220 35808 14272
rect 35860 14260 35866 14272
rect 36817 14263 36875 14269
rect 36817 14260 36829 14263
rect 35860 14232 36829 14260
rect 35860 14220 35866 14232
rect 36817 14229 36829 14232
rect 36863 14229 36875 14263
rect 36817 14223 36875 14229
rect 1104 14170 37812 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 37812 14170
rect 1104 14096 37812 14118
rect 34790 14016 34796 14068
rect 34848 14056 34854 14068
rect 34977 14059 35035 14065
rect 34977 14056 34989 14059
rect 34848 14028 34989 14056
rect 34848 14016 34854 14028
rect 34977 14025 34989 14028
rect 35023 14025 35035 14059
rect 34977 14019 35035 14025
rect 35802 14016 35808 14068
rect 35860 14016 35866 14068
rect 35820 13988 35848 14016
rect 35636 13960 35848 13988
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13920 2743 13923
rect 2869 13923 2927 13929
rect 2869 13920 2881 13923
rect 2731 13892 2881 13920
rect 2731 13889 2743 13892
rect 2685 13883 2743 13889
rect 2869 13889 2881 13892
rect 2915 13889 2927 13923
rect 2869 13883 2927 13889
rect 25314 13880 25320 13932
rect 25372 13880 25378 13932
rect 35636 13929 35664 13960
rect 35621 13923 35679 13929
rect 35621 13889 35633 13923
rect 35667 13889 35679 13923
rect 35621 13883 35679 13889
rect 35710 13880 35716 13932
rect 35768 13920 35774 13932
rect 35805 13923 35863 13929
rect 35805 13920 35817 13923
rect 35768 13892 35817 13920
rect 35768 13880 35774 13892
rect 35805 13889 35817 13892
rect 35851 13889 35863 13923
rect 35805 13883 35863 13889
rect 2409 13855 2467 13861
rect 2409 13821 2421 13855
rect 2455 13852 2467 13855
rect 2590 13852 2596 13864
rect 2455 13824 2596 13852
rect 2455 13821 2467 13824
rect 2409 13815 2467 13821
rect 2590 13812 2596 13824
rect 2648 13812 2654 13864
rect 3513 13855 3571 13861
rect 3513 13821 3525 13855
rect 3559 13821 3571 13855
rect 3513 13815 3571 13821
rect 3528 13784 3556 13815
rect 4062 13812 4068 13864
rect 4120 13852 4126 13864
rect 4341 13855 4399 13861
rect 4341 13852 4353 13855
rect 4120 13824 4353 13852
rect 4120 13812 4126 13824
rect 4341 13821 4353 13824
rect 4387 13821 4399 13855
rect 4341 13815 4399 13821
rect 25961 13855 26019 13861
rect 25961 13821 25973 13855
rect 26007 13852 26019 13855
rect 29454 13852 29460 13864
rect 26007 13824 29460 13852
rect 26007 13821 26019 13824
rect 25961 13815 26019 13821
rect 29454 13812 29460 13824
rect 29512 13812 29518 13864
rect 36262 13812 36268 13864
rect 36320 13812 36326 13864
rect 3786 13784 3792 13796
rect 3528 13756 3792 13784
rect 3786 13744 3792 13756
rect 3844 13744 3850 13796
rect 2958 13676 2964 13728
rect 3016 13716 3022 13728
rect 3605 13719 3663 13725
rect 3605 13716 3617 13719
rect 3016 13688 3617 13716
rect 3016 13676 3022 13688
rect 3605 13685 3617 13688
rect 3651 13685 3663 13719
rect 3605 13679 3663 13685
rect 1104 13626 37812 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 37812 13626
rect 1104 13552 37812 13574
rect 2866 13472 2872 13524
rect 2924 13472 2930 13524
rect 35161 13447 35219 13453
rect 35161 13413 35173 13447
rect 35207 13444 35219 13447
rect 35434 13444 35440 13456
rect 35207 13416 35440 13444
rect 35207 13413 35219 13416
rect 35161 13407 35219 13413
rect 35434 13404 35440 13416
rect 35492 13404 35498 13456
rect 934 13336 940 13388
rect 992 13376 998 13388
rect 1581 13379 1639 13385
rect 1581 13376 1593 13379
rect 992 13348 1593 13376
rect 992 13336 998 13348
rect 1581 13345 1593 13348
rect 1627 13345 1639 13379
rect 1581 13339 1639 13345
rect 3418 13336 3424 13388
rect 3476 13336 3482 13388
rect 6546 13336 6552 13388
rect 6604 13336 6610 13388
rect 23198 13336 23204 13388
rect 23256 13336 23262 13388
rect 37185 13379 37243 13385
rect 37185 13345 37197 13379
rect 37231 13376 37243 13379
rect 37274 13376 37280 13388
rect 37231 13348 37280 13376
rect 37231 13345 37243 13348
rect 37185 13339 37243 13345
rect 37274 13336 37280 13348
rect 37332 13336 37338 13388
rect 2590 13268 2596 13320
rect 2648 13268 2654 13320
rect 3786 13268 3792 13320
rect 3844 13268 3850 13320
rect 11054 13268 11060 13320
rect 11112 13308 11118 13320
rect 13078 13308 13084 13320
rect 11112 13280 13084 13308
rect 11112 13268 11118 13280
rect 13078 13268 13084 13280
rect 13136 13268 13142 13320
rect 24854 13268 24860 13320
rect 24912 13308 24918 13320
rect 25777 13311 25835 13317
rect 25777 13308 25789 13311
rect 24912 13280 25789 13308
rect 24912 13268 24918 13280
rect 25777 13277 25789 13280
rect 25823 13308 25835 13311
rect 28902 13308 28908 13320
rect 25823 13280 28908 13308
rect 25823 13277 25835 13280
rect 25777 13271 25835 13277
rect 28902 13268 28908 13280
rect 28960 13268 28966 13320
rect 35986 13268 35992 13320
rect 36044 13268 36050 13320
rect 36262 13268 36268 13320
rect 36320 13268 36326 13320
rect 34793 13243 34851 13249
rect 34793 13240 34805 13243
rect 34532 13212 34805 13240
rect 34532 13184 34560 13212
rect 34793 13209 34805 13212
rect 34839 13209 34851 13243
rect 35526 13240 35532 13252
rect 34793 13203 34851 13209
rect 35268 13212 35532 13240
rect 4430 13132 4436 13184
rect 4488 13132 4494 13184
rect 7190 13132 7196 13184
rect 7248 13132 7254 13184
rect 10410 13132 10416 13184
rect 10468 13132 10474 13184
rect 23750 13132 23756 13184
rect 23808 13132 23814 13184
rect 25958 13132 25964 13184
rect 26016 13132 26022 13184
rect 34514 13132 34520 13184
rect 34572 13132 34578 13184
rect 35268 13181 35296 13212
rect 35526 13200 35532 13212
rect 35584 13200 35590 13252
rect 35253 13175 35311 13181
rect 35253 13141 35265 13175
rect 35299 13141 35311 13175
rect 35253 13135 35311 13141
rect 35345 13175 35403 13181
rect 35345 13141 35357 13175
rect 35391 13172 35403 13175
rect 35434 13172 35440 13184
rect 35391 13144 35440 13172
rect 35391 13141 35403 13144
rect 35345 13135 35403 13141
rect 35434 13132 35440 13144
rect 35492 13132 35498 13184
rect 1104 13082 37812 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 37812 13082
rect 1104 13008 37812 13030
rect 3329 12971 3387 12977
rect 3329 12937 3341 12971
rect 3375 12968 3387 12971
rect 3786 12968 3792 12980
rect 3375 12940 3792 12968
rect 3375 12937 3387 12940
rect 3329 12931 3387 12937
rect 3786 12928 3792 12940
rect 3844 12928 3850 12980
rect 4430 12928 4436 12980
rect 4488 12928 4494 12980
rect 35434 12928 35440 12980
rect 35492 12928 35498 12980
rect 35526 12928 35532 12980
rect 35584 12928 35590 12980
rect 35986 12928 35992 12980
rect 36044 12968 36050 12980
rect 36817 12971 36875 12977
rect 36817 12968 36829 12971
rect 36044 12940 36829 12968
rect 36044 12928 36050 12940
rect 36817 12937 36829 12940
rect 36863 12937 36875 12971
rect 36817 12931 36875 12937
rect 1964 12872 3556 12900
rect 1964 12844 1992 12872
rect 3528 12844 3556 12872
rect 1946 12792 1952 12844
rect 2004 12792 2010 12844
rect 2216 12835 2274 12841
rect 2216 12801 2228 12835
rect 2262 12832 2274 12835
rect 2958 12832 2964 12844
rect 2262 12804 2964 12832
rect 2262 12801 2274 12804
rect 2216 12795 2274 12801
rect 2958 12792 2964 12804
rect 3016 12792 3022 12844
rect 3510 12792 3516 12844
rect 3568 12792 3574 12844
rect 4065 12835 4123 12841
rect 4065 12801 4077 12835
rect 4111 12832 4123 12835
rect 4448 12832 4476 12928
rect 13814 12860 13820 12912
rect 13872 12900 13878 12912
rect 14430 12903 14488 12909
rect 14430 12900 14442 12903
rect 13872 12872 14442 12900
rect 13872 12860 13878 12872
rect 14430 12869 14442 12872
rect 14476 12869 14488 12903
rect 35452 12900 35480 12928
rect 14430 12863 14488 12869
rect 35268 12872 35480 12900
rect 35544 12900 35572 12928
rect 35682 12903 35740 12909
rect 35682 12900 35694 12903
rect 35544 12872 35694 12900
rect 4111 12804 4476 12832
rect 14185 12835 14243 12841
rect 4111 12801 4123 12804
rect 4065 12795 4123 12801
rect 14185 12801 14197 12835
rect 14231 12832 14243 12835
rect 14274 12832 14280 12844
rect 14231 12804 14280 12832
rect 14231 12801 14243 12804
rect 14185 12795 14243 12801
rect 14274 12792 14280 12804
rect 14332 12792 14338 12844
rect 35268 12841 35296 12872
rect 35682 12869 35694 12872
rect 35728 12869 35740 12903
rect 35682 12863 35740 12869
rect 35253 12835 35311 12841
rect 35253 12801 35265 12835
rect 35299 12801 35311 12835
rect 35253 12795 35311 12801
rect 35342 12792 35348 12844
rect 35400 12832 35406 12844
rect 35437 12835 35495 12841
rect 35437 12832 35449 12835
rect 35400 12804 35449 12832
rect 35400 12792 35406 12804
rect 35437 12801 35449 12804
rect 35483 12801 35495 12835
rect 35437 12795 35495 12801
rect 3418 12588 3424 12640
rect 3476 12588 3482 12640
rect 15565 12631 15623 12637
rect 15565 12597 15577 12631
rect 15611 12628 15623 12631
rect 17218 12628 17224 12640
rect 15611 12600 17224 12628
rect 15611 12597 15623 12600
rect 15565 12591 15623 12597
rect 17218 12588 17224 12600
rect 17276 12588 17282 12640
rect 34698 12588 34704 12640
rect 34756 12588 34762 12640
rect 1104 12538 37812 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 37812 12538
rect 1104 12464 37812 12486
rect 3418 12248 3424 12300
rect 3476 12248 3482 12300
rect 34698 12248 34704 12300
rect 34756 12288 34762 12300
rect 35345 12291 35403 12297
rect 35345 12288 35357 12291
rect 34756 12260 35357 12288
rect 34756 12248 34762 12260
rect 35345 12257 35357 12260
rect 35391 12257 35403 12291
rect 35345 12251 35403 12257
rect 2685 12223 2743 12229
rect 2685 12189 2697 12223
rect 2731 12220 2743 12223
rect 2869 12223 2927 12229
rect 2869 12220 2881 12223
rect 2731 12192 2881 12220
rect 2731 12189 2743 12192
rect 2685 12183 2743 12189
rect 2869 12189 2881 12192
rect 2915 12189 2927 12223
rect 2869 12183 2927 12189
rect 35989 12223 36047 12229
rect 35989 12189 36001 12223
rect 36035 12220 36047 12223
rect 36173 12223 36231 12229
rect 36173 12220 36185 12223
rect 36035 12192 36185 12220
rect 36035 12189 36047 12192
rect 35989 12183 36047 12189
rect 36173 12189 36185 12192
rect 36219 12189 36231 12223
rect 36173 12183 36231 12189
rect 2317 12155 2375 12161
rect 2317 12121 2329 12155
rect 2363 12121 2375 12155
rect 2317 12115 2375 12121
rect 2332 12084 2360 12115
rect 36538 12112 36544 12164
rect 36596 12112 36602 12164
rect 2590 12084 2596 12096
rect 2332 12056 2596 12084
rect 2590 12044 2596 12056
rect 2648 12044 2654 12096
rect 34514 12044 34520 12096
rect 34572 12084 34578 12096
rect 34977 12087 35035 12093
rect 34977 12084 34989 12087
rect 34572 12056 34989 12084
rect 34572 12044 34578 12056
rect 34977 12053 34989 12056
rect 35023 12053 35035 12087
rect 34977 12047 35035 12053
rect 1104 11994 37812 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 37812 11994
rect 1104 11920 37812 11942
rect 36538 11840 36544 11892
rect 36596 11840 36602 11892
rect 934 11772 940 11824
rect 992 11812 998 11824
rect 1581 11815 1639 11821
rect 1581 11812 1593 11815
rect 992 11784 1593 11812
rect 992 11772 998 11784
rect 1581 11781 1593 11784
rect 1627 11781 1639 11815
rect 1581 11775 1639 11781
rect 2590 11704 2596 11756
rect 2648 11704 2654 11756
rect 3513 11747 3571 11753
rect 3513 11713 3525 11747
rect 3559 11744 3571 11747
rect 3694 11744 3700 11756
rect 3559 11716 3700 11744
rect 3559 11713 3571 11716
rect 3513 11707 3571 11713
rect 3694 11704 3700 11716
rect 3752 11704 3758 11756
rect 35897 11747 35955 11753
rect 35897 11713 35909 11747
rect 35943 11744 35955 11747
rect 36556 11744 36584 11840
rect 36909 11815 36967 11821
rect 36909 11781 36921 11815
rect 36955 11812 36967 11815
rect 37458 11812 37464 11824
rect 36955 11784 37464 11812
rect 36955 11781 36967 11784
rect 36909 11775 36967 11781
rect 37458 11772 37464 11784
rect 37516 11772 37522 11824
rect 35943 11716 36584 11744
rect 35943 11713 35955 11716
rect 35897 11707 35955 11713
rect 4065 11679 4123 11685
rect 4065 11645 4077 11679
rect 4111 11645 4123 11679
rect 4065 11639 4123 11645
rect 34425 11679 34483 11685
rect 34425 11645 34437 11679
rect 34471 11676 34483 11679
rect 34514 11676 34520 11688
rect 34471 11648 34520 11676
rect 34471 11645 34483 11648
rect 34425 11639 34483 11645
rect 3697 11611 3755 11617
rect 3697 11608 3709 11611
rect 3436 11580 3709 11608
rect 3436 11552 3464 11580
rect 3697 11577 3709 11580
rect 3743 11577 3755 11611
rect 3697 11571 3755 11577
rect 4080 11552 4108 11639
rect 34514 11636 34520 11648
rect 34572 11636 34578 11688
rect 35069 11679 35127 11685
rect 35069 11645 35081 11679
rect 35115 11676 35127 11679
rect 35434 11676 35440 11688
rect 35115 11648 35440 11676
rect 35115 11645 35127 11648
rect 35069 11639 35127 11645
rect 35434 11636 35440 11648
rect 35492 11636 35498 11688
rect 34698 11568 34704 11620
rect 34756 11568 34762 11620
rect 2866 11500 2872 11552
rect 2924 11500 2930 11552
rect 3418 11500 3424 11552
rect 3476 11500 3482 11552
rect 3602 11500 3608 11552
rect 3660 11500 3666 11552
rect 4062 11500 4068 11552
rect 4120 11540 4126 11552
rect 4341 11543 4399 11549
rect 4341 11540 4353 11543
rect 4120 11512 4353 11540
rect 4120 11500 4126 11512
rect 4341 11509 4353 11512
rect 4387 11509 4399 11543
rect 4341 11503 4399 11509
rect 34885 11543 34943 11549
rect 34885 11509 34897 11543
rect 34931 11540 34943 11543
rect 35526 11540 35532 11552
rect 34931 11512 35532 11540
rect 34931 11509 34943 11512
rect 34885 11503 34943 11509
rect 35526 11500 35532 11512
rect 35584 11500 35590 11552
rect 35618 11500 35624 11552
rect 35676 11500 35682 11552
rect 1104 11450 37812 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 37812 11450
rect 1104 11376 37812 11398
rect 3602 11336 3608 11348
rect 2976 11308 3608 11336
rect 1946 11160 1952 11212
rect 2004 11160 2010 11212
rect 2216 11135 2274 11141
rect 2216 11101 2228 11135
rect 2262 11132 2274 11135
rect 2976 11132 3004 11308
rect 3602 11296 3608 11308
rect 3660 11296 3666 11348
rect 35345 11339 35403 11345
rect 35345 11305 35357 11339
rect 35391 11336 35403 11339
rect 35434 11336 35440 11348
rect 35391 11308 35440 11336
rect 35391 11305 35403 11308
rect 35345 11299 35403 11305
rect 35434 11296 35440 11308
rect 35492 11296 35498 11348
rect 3329 11271 3387 11277
rect 3329 11237 3341 11271
rect 3375 11268 3387 11271
rect 3375 11240 4384 11268
rect 3375 11237 3387 11240
rect 3329 11231 3387 11237
rect 4356 11209 4384 11240
rect 4341 11203 4399 11209
rect 4341 11169 4353 11203
rect 4387 11169 4399 11203
rect 4341 11163 4399 11169
rect 35342 11160 35348 11212
rect 35400 11200 35406 11212
rect 35437 11203 35495 11209
rect 35437 11200 35449 11203
rect 35400 11172 35449 11200
rect 35400 11160 35406 11172
rect 35437 11169 35449 11172
rect 35483 11169 35495 11203
rect 35437 11163 35495 11169
rect 2262 11104 3004 11132
rect 2262 11101 2274 11104
rect 2216 11095 2274 11101
rect 34790 11092 34796 11144
rect 34848 11092 34854 11144
rect 35526 11092 35532 11144
rect 35584 11132 35590 11144
rect 35693 11135 35751 11141
rect 35693 11132 35705 11135
rect 35584 11104 35705 11132
rect 35584 11092 35590 11104
rect 35693 11101 35705 11104
rect 35739 11101 35751 11135
rect 35693 11095 35751 11101
rect 3510 10956 3516 11008
rect 3568 10996 3574 11008
rect 3789 10999 3847 11005
rect 3789 10996 3801 10999
rect 3568 10968 3801 10996
rect 3568 10956 3574 10968
rect 3789 10965 3801 10968
rect 3835 10965 3847 10999
rect 3789 10959 3847 10965
rect 36814 10956 36820 11008
rect 36872 10956 36878 11008
rect 1104 10906 37812 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 37812 10906
rect 1104 10832 37812 10854
rect 28902 10752 28908 10804
rect 28960 10752 28966 10804
rect 34790 10752 34796 10804
rect 34848 10792 34854 10804
rect 34977 10795 35035 10801
rect 34977 10792 34989 10795
rect 34848 10764 34989 10792
rect 34848 10752 34854 10764
rect 34977 10761 34989 10764
rect 35023 10761 35035 10795
rect 34977 10755 35035 10761
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10656 2743 10659
rect 2869 10659 2927 10665
rect 2869 10656 2881 10659
rect 2731 10628 2881 10656
rect 2731 10625 2743 10628
rect 2685 10619 2743 10625
rect 2869 10625 2881 10628
rect 2915 10625 2927 10659
rect 2869 10619 2927 10625
rect 17218 10616 17224 10668
rect 17276 10616 17282 10668
rect 27890 10616 27896 10668
rect 27948 10656 27954 10668
rect 28534 10656 28540 10668
rect 27948 10628 28540 10656
rect 27948 10616 27954 10628
rect 28534 10616 28540 10628
rect 28592 10616 28598 10668
rect 29454 10616 29460 10668
rect 29512 10616 29518 10668
rect 35618 10616 35624 10668
rect 35676 10656 35682 10668
rect 35805 10659 35863 10665
rect 35805 10656 35817 10659
rect 35676 10628 35817 10656
rect 35676 10616 35682 10628
rect 35805 10625 35817 10628
rect 35851 10625 35863 10659
rect 36814 10656 36820 10668
rect 35805 10619 35863 10625
rect 36004 10628 36820 10656
rect 2409 10591 2467 10597
rect 2409 10557 2421 10591
rect 2455 10588 2467 10591
rect 3421 10591 3479 10597
rect 3421 10588 3433 10591
rect 2455 10560 2636 10588
rect 2455 10557 2467 10560
rect 2409 10551 2467 10557
rect 2608 10464 2636 10560
rect 2884 10560 3433 10588
rect 2884 10464 2912 10560
rect 3421 10557 3433 10560
rect 3467 10588 3479 10591
rect 4065 10591 4123 10597
rect 3467 10560 3740 10588
rect 3467 10557 3479 10560
rect 3421 10551 3479 10557
rect 3712 10529 3740 10560
rect 4065 10557 4077 10591
rect 4111 10557 4123 10591
rect 4065 10551 4123 10557
rect 35529 10591 35587 10597
rect 35529 10557 35541 10591
rect 35575 10588 35587 10591
rect 36004 10588 36032 10628
rect 36814 10616 36820 10628
rect 36872 10616 36878 10668
rect 35575 10560 36032 10588
rect 35575 10557 35587 10560
rect 35529 10551 35587 10557
rect 3697 10523 3755 10529
rect 3697 10489 3709 10523
rect 3743 10489 3755 10523
rect 3697 10483 3755 10489
rect 4080 10464 4108 10551
rect 36078 10548 36084 10600
rect 36136 10548 36142 10600
rect 2590 10412 2596 10464
rect 2648 10412 2654 10464
rect 2866 10412 2872 10464
rect 2924 10412 2930 10464
rect 3602 10412 3608 10464
rect 3660 10412 3666 10464
rect 4062 10412 4068 10464
rect 4120 10452 4126 10464
rect 4341 10455 4399 10461
rect 4341 10452 4353 10455
rect 4120 10424 4353 10452
rect 4120 10412 4126 10424
rect 4341 10421 4353 10424
rect 4387 10421 4399 10455
rect 4341 10415 4399 10421
rect 17865 10455 17923 10461
rect 17865 10421 17877 10455
rect 17911 10452 17923 10455
rect 19334 10452 19340 10464
rect 17911 10424 19340 10452
rect 17911 10421 17923 10424
rect 17865 10415 17923 10421
rect 19334 10412 19340 10424
rect 19392 10412 19398 10464
rect 27338 10412 27344 10464
rect 27396 10412 27402 10464
rect 1104 10362 37812 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 37812 10362
rect 1104 10288 37812 10310
rect 2866 10208 2872 10260
rect 2924 10208 2930 10260
rect 7561 10251 7619 10257
rect 7561 10217 7573 10251
rect 7607 10248 7619 10251
rect 11054 10248 11060 10260
rect 7607 10220 11060 10248
rect 7607 10217 7619 10220
rect 7561 10211 7619 10217
rect 11054 10208 11060 10220
rect 11112 10208 11118 10260
rect 22922 10208 22928 10260
rect 22980 10208 22986 10260
rect 35161 10183 35219 10189
rect 35161 10149 35173 10183
rect 35207 10180 35219 10183
rect 35434 10180 35440 10192
rect 35207 10152 35440 10180
rect 35207 10149 35219 10152
rect 35161 10143 35219 10149
rect 35434 10140 35440 10152
rect 35492 10140 35498 10192
rect 934 10072 940 10124
rect 992 10112 998 10124
rect 1581 10115 1639 10121
rect 1581 10112 1593 10115
rect 992 10084 1593 10112
rect 992 10072 998 10084
rect 1581 10081 1593 10084
rect 1627 10081 1639 10115
rect 1581 10075 1639 10081
rect 7009 10115 7067 10121
rect 7009 10081 7021 10115
rect 7055 10112 7067 10115
rect 7190 10112 7196 10124
rect 7055 10084 7196 10112
rect 7055 10081 7067 10084
rect 7009 10075 7067 10081
rect 7190 10072 7196 10084
rect 7248 10072 7254 10124
rect 23569 10115 23627 10121
rect 23569 10081 23581 10115
rect 23615 10112 23627 10115
rect 23750 10112 23756 10124
rect 23615 10084 23756 10112
rect 23615 10081 23627 10084
rect 23569 10075 23627 10081
rect 23750 10072 23756 10084
rect 23808 10072 23814 10124
rect 35253 10115 35311 10121
rect 35253 10081 35265 10115
rect 35299 10112 35311 10115
rect 35526 10112 35532 10124
rect 35299 10084 35532 10112
rect 35299 10081 35311 10084
rect 35253 10075 35311 10081
rect 35526 10072 35532 10084
rect 35584 10072 35590 10124
rect 36078 10072 36084 10124
rect 36136 10072 36142 10124
rect 37185 10115 37243 10121
rect 37185 10081 37197 10115
rect 37231 10112 37243 10115
rect 37274 10112 37280 10124
rect 37231 10084 37280 10112
rect 37231 10081 37243 10084
rect 37185 10075 37243 10081
rect 37274 10072 37280 10084
rect 37332 10072 37338 10124
rect 2590 10004 2596 10056
rect 2648 10004 2654 10056
rect 3510 10004 3516 10056
rect 3568 10004 3574 10056
rect 3786 10004 3792 10056
rect 3844 10004 3850 10056
rect 16850 10004 16856 10056
rect 16908 10044 16914 10056
rect 17037 10047 17095 10053
rect 17037 10044 17049 10047
rect 16908 10016 17049 10044
rect 16908 10004 16914 10016
rect 17037 10013 17049 10016
rect 17083 10044 17095 10047
rect 17313 10047 17371 10053
rect 17313 10044 17325 10047
rect 17083 10016 17325 10044
rect 17083 10013 17095 10016
rect 17037 10007 17095 10013
rect 17313 10013 17325 10016
rect 17359 10044 17371 10047
rect 20898 10044 20904 10056
rect 17359 10016 20904 10044
rect 17359 10013 17371 10016
rect 17313 10007 17371 10013
rect 20898 10004 20904 10016
rect 20956 10004 20962 10056
rect 32953 10047 33011 10053
rect 32953 10013 32965 10047
rect 32999 10044 33011 10047
rect 35342 10044 35348 10056
rect 32999 10016 35348 10044
rect 32999 10013 33011 10016
rect 32953 10007 33011 10013
rect 35342 10004 35348 10016
rect 35400 10004 35406 10056
rect 35986 10004 35992 10056
rect 36044 10004 36050 10056
rect 36096 10044 36124 10072
rect 36173 10047 36231 10053
rect 36173 10044 36185 10047
rect 36096 10016 36185 10044
rect 36173 10013 36185 10016
rect 36219 10013 36231 10047
rect 36173 10007 36231 10013
rect 31205 9979 31263 9985
rect 31205 9945 31217 9979
rect 31251 9945 31263 9979
rect 31205 9939 31263 9945
rect 4430 9868 4436 9920
rect 4488 9868 4494 9920
rect 17126 9868 17132 9920
rect 17184 9868 17190 9920
rect 31018 9868 31024 9920
rect 31076 9908 31082 9920
rect 31220 9908 31248 9939
rect 34514 9936 34520 9988
rect 34572 9976 34578 9988
rect 34793 9979 34851 9985
rect 34793 9976 34805 9979
rect 34572 9948 34805 9976
rect 34572 9936 34578 9948
rect 34793 9945 34805 9948
rect 34839 9976 34851 9979
rect 35802 9976 35808 9988
rect 34839 9948 35808 9976
rect 34839 9945 34851 9948
rect 34793 9939 34851 9945
rect 35802 9936 35808 9948
rect 35860 9936 35866 9988
rect 31076 9880 31248 9908
rect 35345 9911 35403 9917
rect 31076 9868 31082 9880
rect 35345 9877 35357 9911
rect 35391 9908 35403 9911
rect 35434 9908 35440 9920
rect 35391 9880 35440 9908
rect 35391 9877 35403 9880
rect 35345 9871 35403 9877
rect 35434 9868 35440 9880
rect 35492 9868 35498 9920
rect 1104 9818 37812 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 37812 9818
rect 1104 9744 37812 9766
rect 3329 9707 3387 9713
rect 3329 9673 3341 9707
rect 3375 9704 3387 9707
rect 3786 9704 3792 9716
rect 3375 9676 3792 9704
rect 3375 9673 3387 9676
rect 3329 9667 3387 9673
rect 3786 9664 3792 9676
rect 3844 9664 3850 9716
rect 8662 9664 8668 9716
rect 8720 9704 8726 9716
rect 17126 9704 17132 9716
rect 8720 9676 17132 9704
rect 8720 9664 8726 9676
rect 17126 9664 17132 9676
rect 17184 9664 17190 9716
rect 35434 9704 35440 9716
rect 35268 9676 35440 9704
rect 2216 9639 2274 9645
rect 2216 9605 2228 9639
rect 2262 9636 2274 9639
rect 3602 9636 3608 9648
rect 2262 9608 3608 9636
rect 2262 9605 2274 9608
rect 2216 9599 2274 9605
rect 3602 9596 3608 9608
rect 3660 9596 3666 9648
rect 1946 9528 1952 9580
rect 2004 9528 2010 9580
rect 4065 9571 4123 9577
rect 4065 9537 4077 9571
rect 4111 9568 4123 9571
rect 4430 9568 4436 9580
rect 4111 9540 4436 9568
rect 4111 9537 4123 9540
rect 4065 9531 4123 9537
rect 4430 9528 4436 9540
rect 4488 9528 4494 9580
rect 35268 9577 35296 9676
rect 35434 9664 35440 9676
rect 35492 9664 35498 9716
rect 35986 9664 35992 9716
rect 36044 9704 36050 9716
rect 36817 9707 36875 9713
rect 36817 9704 36829 9707
rect 36044 9676 36829 9704
rect 36044 9664 36050 9676
rect 36817 9673 36829 9676
rect 36863 9673 36875 9707
rect 36817 9667 36875 9673
rect 35526 9596 35532 9648
rect 35584 9636 35590 9648
rect 35682 9639 35740 9645
rect 35682 9636 35694 9639
rect 35584 9608 35694 9636
rect 35584 9596 35590 9608
rect 35682 9605 35694 9608
rect 35728 9605 35740 9639
rect 35682 9599 35740 9605
rect 35253 9571 35311 9577
rect 35253 9537 35265 9571
rect 35299 9537 35311 9571
rect 35253 9531 35311 9537
rect 35342 9528 35348 9580
rect 35400 9568 35406 9580
rect 35437 9571 35495 9577
rect 35437 9568 35449 9571
rect 35400 9540 35449 9568
rect 35400 9528 35406 9540
rect 35437 9537 35449 9540
rect 35483 9537 35495 9571
rect 35437 9531 35495 9537
rect 3418 9324 3424 9376
rect 3476 9324 3482 9376
rect 34698 9324 34704 9376
rect 34756 9324 34762 9376
rect 1104 9274 37812 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 37812 9274
rect 1104 9200 37812 9222
rect 3418 9120 3424 9172
rect 3476 9120 3482 9172
rect 34698 9120 34704 9172
rect 34756 9120 34762 9172
rect 3436 9033 3464 9120
rect 3421 9027 3479 9033
rect 3421 8993 3433 9027
rect 3467 8993 3479 9027
rect 34716 9024 34744 9120
rect 35345 9027 35403 9033
rect 35345 9024 35357 9027
rect 34716 8996 35357 9024
rect 3421 8987 3479 8993
rect 35345 8993 35357 8996
rect 35391 8993 35403 9027
rect 35345 8987 35403 8993
rect 2685 8959 2743 8965
rect 2685 8925 2697 8959
rect 2731 8956 2743 8959
rect 2869 8959 2927 8965
rect 2869 8956 2881 8959
rect 2731 8928 2881 8956
rect 2731 8925 2743 8928
rect 2685 8919 2743 8925
rect 2869 8925 2881 8928
rect 2915 8925 2927 8959
rect 2869 8919 2927 8925
rect 35989 8959 36047 8965
rect 35989 8925 36001 8959
rect 36035 8956 36047 8959
rect 36173 8959 36231 8965
rect 36173 8956 36185 8959
rect 36035 8928 36185 8956
rect 36035 8925 36047 8928
rect 35989 8919 36047 8925
rect 36173 8925 36185 8928
rect 36219 8925 36231 8959
rect 36173 8919 36231 8925
rect 2317 8891 2375 8897
rect 2317 8857 2329 8891
rect 2363 8857 2375 8891
rect 2317 8851 2375 8857
rect 2332 8820 2360 8851
rect 36538 8848 36544 8900
rect 36596 8848 36602 8900
rect 2590 8820 2596 8832
rect 2332 8792 2596 8820
rect 2590 8780 2596 8792
rect 2648 8780 2654 8832
rect 34514 8780 34520 8832
rect 34572 8820 34578 8832
rect 34977 8823 35035 8829
rect 34977 8820 34989 8823
rect 34572 8792 34989 8820
rect 34572 8780 34578 8792
rect 34977 8789 34989 8792
rect 35023 8789 35035 8823
rect 34977 8783 35035 8789
rect 1104 8730 37812 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 37812 8730
rect 1104 8656 37812 8678
rect 3418 8576 3424 8628
rect 3476 8576 3482 8628
rect 34698 8576 34704 8628
rect 34756 8576 34762 8628
rect 36538 8576 36544 8628
rect 36596 8576 36602 8628
rect 934 8508 940 8560
rect 992 8548 998 8560
rect 1581 8551 1639 8557
rect 1581 8548 1593 8551
rect 992 8520 1593 8548
rect 992 8508 998 8520
rect 1581 8517 1593 8520
rect 1627 8517 1639 8551
rect 1581 8511 1639 8517
rect 2590 8440 2596 8492
rect 2648 8440 2654 8492
rect 3436 8480 3464 8576
rect 3252 8452 3464 8480
rect 3053 8347 3111 8353
rect 3053 8313 3065 8347
rect 3099 8344 3111 8347
rect 3252 8344 3280 8452
rect 3329 8415 3387 8421
rect 3329 8381 3341 8415
rect 3375 8412 3387 8415
rect 34425 8415 34483 8421
rect 3375 8384 3556 8412
rect 3375 8381 3387 8384
rect 3329 8375 3387 8381
rect 3099 8316 3280 8344
rect 3528 8344 3556 8384
rect 34425 8381 34437 8415
rect 34471 8412 34483 8415
rect 34514 8412 34520 8424
rect 34471 8384 34520 8412
rect 34471 8381 34483 8384
rect 34425 8375 34483 8381
rect 34514 8372 34520 8384
rect 34572 8372 34578 8424
rect 3697 8347 3755 8353
rect 3697 8344 3709 8347
rect 3528 8316 3709 8344
rect 3099 8313 3111 8316
rect 3053 8307 3111 8313
rect 3697 8313 3709 8316
rect 3743 8344 3755 8347
rect 4062 8344 4068 8356
rect 3743 8316 4068 8344
rect 3743 8313 3755 8316
rect 3697 8307 3755 8313
rect 4062 8304 4068 8316
rect 4120 8344 4126 8356
rect 34716 8353 34744 8576
rect 35897 8483 35955 8489
rect 35897 8449 35909 8483
rect 35943 8480 35955 8483
rect 36556 8480 36584 8576
rect 36909 8551 36967 8557
rect 36909 8517 36921 8551
rect 36955 8548 36967 8551
rect 37458 8548 37464 8560
rect 36955 8520 37464 8548
rect 36955 8517 36967 8520
rect 36909 8511 36967 8517
rect 37458 8508 37464 8520
rect 37516 8508 37522 8560
rect 35943 8452 36584 8480
rect 35943 8449 35955 8452
rect 35897 8443 35955 8449
rect 35069 8415 35127 8421
rect 35069 8381 35081 8415
rect 35115 8412 35127 8415
rect 35434 8412 35440 8424
rect 35115 8384 35440 8412
rect 35115 8381 35127 8384
rect 35069 8375 35127 8381
rect 35434 8372 35440 8384
rect 35492 8372 35498 8424
rect 34701 8347 34759 8353
rect 4120 8316 5488 8344
rect 4120 8304 4126 8316
rect 5460 8288 5488 8316
rect 34701 8313 34713 8347
rect 34747 8313 34759 8347
rect 34701 8307 34759 8313
rect 2774 8236 2780 8288
rect 2832 8276 2838 8288
rect 2869 8279 2927 8285
rect 2869 8276 2881 8279
rect 2832 8248 2881 8276
rect 2832 8236 2838 8248
rect 2869 8245 2881 8248
rect 2915 8245 2927 8279
rect 2869 8239 2927 8245
rect 5442 8236 5448 8288
rect 5500 8236 5506 8288
rect 34885 8279 34943 8285
rect 34885 8245 34897 8279
rect 34931 8276 34943 8279
rect 35526 8276 35532 8288
rect 34931 8248 35532 8276
rect 34931 8245 34943 8248
rect 34885 8239 34943 8245
rect 35526 8236 35532 8248
rect 35584 8236 35590 8288
rect 35618 8236 35624 8288
rect 35676 8236 35682 8288
rect 1104 8186 37812 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 37812 8186
rect 1104 8112 37812 8134
rect 11885 8075 11943 8081
rect 11885 8041 11897 8075
rect 11931 8072 11943 8075
rect 12066 8072 12072 8084
rect 11931 8044 12072 8072
rect 11931 8041 11943 8044
rect 11885 8035 11943 8041
rect 12066 8032 12072 8044
rect 12124 8072 12130 8084
rect 14274 8072 14280 8084
rect 12124 8044 14280 8072
rect 12124 8032 12130 8044
rect 14274 8032 14280 8044
rect 14332 8032 14338 8084
rect 35345 8075 35403 8081
rect 35345 8041 35357 8075
rect 35391 8072 35403 8075
rect 35434 8072 35440 8084
rect 35391 8044 35440 8072
rect 35391 8041 35403 8044
rect 35345 8035 35403 8041
rect 35434 8032 35440 8044
rect 35492 8032 35498 8084
rect 3329 8007 3387 8013
rect 3329 7973 3341 8007
rect 3375 7973 3387 8007
rect 3329 7967 3387 7973
rect 1946 7896 1952 7948
rect 2004 7896 2010 7948
rect 3344 7936 3372 7967
rect 3789 7939 3847 7945
rect 3789 7936 3801 7939
rect 3344 7908 3801 7936
rect 3789 7905 3801 7908
rect 3835 7905 3847 7939
rect 3789 7899 3847 7905
rect 19334 7896 19340 7948
rect 19392 7936 19398 7948
rect 19797 7939 19855 7945
rect 19797 7936 19809 7939
rect 19392 7908 19809 7936
rect 19392 7896 19398 7908
rect 19797 7905 19809 7908
rect 19843 7905 19855 7939
rect 19797 7899 19855 7905
rect 35342 7896 35348 7948
rect 35400 7936 35406 7948
rect 35437 7939 35495 7945
rect 35437 7936 35449 7939
rect 35400 7908 35449 7936
rect 35400 7896 35406 7908
rect 35437 7905 35449 7908
rect 35483 7905 35495 7939
rect 35437 7899 35495 7905
rect 2216 7871 2274 7877
rect 2216 7837 2228 7871
rect 2262 7868 2274 7871
rect 2774 7868 2780 7880
rect 2262 7840 2780 7868
rect 2262 7837 2274 7840
rect 2216 7831 2274 7837
rect 2774 7828 2780 7840
rect 2832 7828 2838 7880
rect 34517 7871 34575 7877
rect 34517 7837 34529 7871
rect 34563 7868 34575 7871
rect 34698 7868 34704 7880
rect 34563 7840 34704 7868
rect 34563 7837 34575 7840
rect 34517 7831 34575 7837
rect 34698 7828 34704 7840
rect 34756 7828 34762 7880
rect 34790 7828 34796 7880
rect 34848 7828 34854 7880
rect 35526 7828 35532 7880
rect 35584 7868 35590 7880
rect 35693 7871 35751 7877
rect 35693 7868 35705 7871
rect 35584 7840 35705 7868
rect 35584 7828 35590 7840
rect 35693 7837 35705 7840
rect 35739 7837 35751 7871
rect 35693 7831 35751 7837
rect 10410 7760 10416 7812
rect 10468 7800 10474 7812
rect 12529 7803 12587 7809
rect 12529 7800 12541 7803
rect 10468 7772 12541 7800
rect 10468 7760 10474 7772
rect 12529 7769 12541 7772
rect 12575 7800 12587 7803
rect 20254 7800 20260 7812
rect 12575 7772 20260 7800
rect 12575 7769 12587 7772
rect 12529 7763 12587 7769
rect 20254 7760 20260 7772
rect 20312 7800 20318 7812
rect 20622 7800 20628 7812
rect 20312 7772 20628 7800
rect 20312 7760 20318 7772
rect 20622 7760 20628 7772
rect 20680 7760 20686 7812
rect 37274 7760 37280 7812
rect 37332 7760 37338 7812
rect 4430 7692 4436 7744
rect 4488 7692 4494 7744
rect 19242 7692 19248 7744
rect 19300 7692 19306 7744
rect 33686 7692 33692 7744
rect 33744 7732 33750 7744
rect 33873 7735 33931 7741
rect 33873 7732 33885 7735
rect 33744 7704 33885 7732
rect 33744 7692 33750 7704
rect 33873 7701 33885 7704
rect 33919 7701 33931 7735
rect 33873 7695 33931 7701
rect 36814 7692 36820 7744
rect 36872 7692 36878 7744
rect 36906 7692 36912 7744
rect 36964 7732 36970 7744
rect 37001 7735 37059 7741
rect 37001 7732 37013 7735
rect 36964 7704 37013 7732
rect 36964 7692 36970 7704
rect 37001 7701 37013 7704
rect 37047 7701 37059 7735
rect 37001 7695 37059 7701
rect 1104 7642 37812 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 37812 7642
rect 1104 7568 37812 7590
rect 9953 7531 10011 7537
rect 9953 7497 9965 7531
rect 9999 7528 10011 7531
rect 10410 7528 10416 7540
rect 9999 7500 10416 7528
rect 9999 7497 10011 7500
rect 9953 7491 10011 7497
rect 3084 7463 3142 7469
rect 3084 7429 3096 7463
rect 3130 7460 3142 7463
rect 4706 7460 4712 7472
rect 3130 7432 4712 7460
rect 3130 7429 3142 7432
rect 3084 7423 3142 7429
rect 4706 7420 4712 7432
rect 4764 7420 4770 7472
rect 9585 7463 9643 7469
rect 9585 7429 9597 7463
rect 9631 7460 9643 7463
rect 9968 7460 9996 7491
rect 10410 7488 10416 7500
rect 10468 7488 10474 7540
rect 20622 7488 20628 7540
rect 20680 7528 20686 7540
rect 28445 7531 28503 7537
rect 28445 7528 28457 7531
rect 20680 7500 28457 7528
rect 20680 7488 20686 7500
rect 28445 7497 28457 7500
rect 28491 7497 28503 7531
rect 28445 7491 28503 7497
rect 9631 7432 9996 7460
rect 28460 7460 28488 7491
rect 34790 7488 34796 7540
rect 34848 7528 34854 7540
rect 34977 7531 35035 7537
rect 34977 7528 34989 7531
rect 34848 7500 34989 7528
rect 34848 7488 34854 7500
rect 34977 7497 34989 7500
rect 35023 7497 35035 7531
rect 36814 7528 36820 7540
rect 34977 7491 35035 7497
rect 35544 7500 36820 7528
rect 28629 7463 28687 7469
rect 28629 7460 28641 7463
rect 28460 7432 28641 7460
rect 9631 7429 9643 7432
rect 9585 7423 9643 7429
rect 28629 7429 28641 7432
rect 28675 7460 28687 7463
rect 31018 7460 31024 7472
rect 28675 7432 31024 7460
rect 28675 7429 28687 7432
rect 28629 7423 28687 7429
rect 31018 7420 31024 7432
rect 31076 7420 31082 7472
rect 1946 7352 1952 7404
rect 2004 7392 2010 7404
rect 3326 7392 3332 7404
rect 2004 7364 3332 7392
rect 2004 7352 2010 7364
rect 3326 7352 3332 7364
rect 3384 7392 3390 7404
rect 35544 7401 35572 7500
rect 36814 7488 36820 7500
rect 36872 7488 36878 7540
rect 7837 7395 7895 7401
rect 7837 7392 7849 7395
rect 3384 7364 7849 7392
rect 3384 7352 3390 7364
rect 7837 7361 7849 7364
rect 7883 7361 7895 7395
rect 7837 7355 7895 7361
rect 35529 7395 35587 7401
rect 35529 7361 35541 7395
rect 35575 7361 35587 7395
rect 35529 7355 35587 7361
rect 35618 7352 35624 7404
rect 35676 7392 35682 7404
rect 35805 7395 35863 7401
rect 35805 7392 35817 7395
rect 35676 7364 35817 7392
rect 35676 7352 35682 7364
rect 35805 7361 35817 7364
rect 35851 7361 35863 7395
rect 35805 7355 35863 7361
rect 4341 7327 4399 7333
rect 4341 7293 4353 7327
rect 4387 7293 4399 7327
rect 4341 7287 4399 7293
rect 4356 7256 4384 7287
rect 4982 7284 4988 7336
rect 5040 7284 5046 7336
rect 5442 7284 5448 7336
rect 5500 7324 5506 7336
rect 5629 7327 5687 7333
rect 5629 7324 5641 7327
rect 5500 7296 5641 7324
rect 5500 7284 5506 7296
rect 5629 7293 5641 7296
rect 5675 7324 5687 7327
rect 5905 7327 5963 7333
rect 5905 7324 5917 7327
rect 5675 7296 5917 7324
rect 5675 7293 5687 7296
rect 5629 7287 5687 7293
rect 5905 7293 5917 7296
rect 5951 7293 5963 7327
rect 5905 7287 5963 7293
rect 33502 7284 33508 7336
rect 33560 7284 33566 7336
rect 34330 7284 34336 7336
rect 34388 7324 34394 7336
rect 34793 7327 34851 7333
rect 34793 7324 34805 7327
rect 34388 7296 34805 7324
rect 34388 7284 34394 7296
rect 34793 7293 34805 7296
rect 34839 7293 34851 7327
rect 34793 7287 34851 7293
rect 36170 7284 36176 7336
rect 36228 7284 36234 7336
rect 4798 7256 4804 7268
rect 4356 7228 4804 7256
rect 4798 7216 4804 7228
rect 4856 7256 4862 7268
rect 5261 7259 5319 7265
rect 5261 7256 5273 7259
rect 4856 7228 5273 7256
rect 4856 7216 4862 7228
rect 5261 7225 5273 7228
rect 5307 7225 5319 7259
rect 5261 7219 5319 7225
rect 26206 7228 29592 7256
rect 1949 7191 2007 7197
rect 1949 7157 1961 7191
rect 1995 7188 2007 7191
rect 3418 7188 3424 7200
rect 1995 7160 3424 7188
rect 1995 7157 2007 7160
rect 1949 7151 2007 7157
rect 3418 7148 3424 7160
rect 3476 7148 3482 7200
rect 3694 7148 3700 7200
rect 3752 7148 3758 7200
rect 3786 7148 3792 7200
rect 3844 7188 3850 7200
rect 4433 7191 4491 7197
rect 4433 7188 4445 7191
rect 3844 7160 4445 7188
rect 3844 7148 3850 7160
rect 4433 7157 4445 7160
rect 4479 7157 4491 7191
rect 4433 7151 4491 7157
rect 5166 7148 5172 7200
rect 5224 7148 5230 7200
rect 24394 7148 24400 7200
rect 24452 7188 24458 7200
rect 26206 7188 26234 7228
rect 29564 7200 29592 7228
rect 24452 7160 26234 7188
rect 24452 7148 24458 7160
rect 29546 7148 29552 7200
rect 29604 7188 29610 7200
rect 29917 7191 29975 7197
rect 29917 7188 29929 7191
rect 29604 7160 29929 7188
rect 29604 7148 29610 7160
rect 29917 7157 29929 7160
rect 29963 7157 29975 7191
rect 29917 7151 29975 7157
rect 33962 7148 33968 7200
rect 34020 7188 34026 7200
rect 34149 7191 34207 7197
rect 34149 7188 34161 7191
rect 34020 7160 34161 7188
rect 34020 7148 34026 7160
rect 34149 7157 34161 7160
rect 34195 7157 34207 7191
rect 34149 7151 34207 7157
rect 34238 7148 34244 7200
rect 34296 7148 34302 7200
rect 1104 7098 37812 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 37812 7098
rect 1104 7024 37812 7046
rect 4798 6984 4804 6996
rect 4356 6956 4804 6984
rect 3326 6808 3332 6860
rect 3384 6808 3390 6860
rect 3789 6851 3847 6857
rect 3789 6817 3801 6851
rect 3835 6848 3847 6851
rect 4356 6848 4384 6956
rect 4798 6944 4804 6956
rect 4856 6944 4862 6996
rect 4709 6919 4767 6925
rect 4709 6885 4721 6919
rect 4755 6916 4767 6919
rect 4982 6916 4988 6928
rect 4755 6888 4988 6916
rect 4755 6885 4767 6888
rect 4709 6879 4767 6885
rect 4982 6876 4988 6888
rect 5040 6876 5046 6928
rect 35161 6919 35219 6925
rect 35161 6885 35173 6919
rect 35207 6916 35219 6919
rect 35434 6916 35440 6928
rect 35207 6888 35440 6916
rect 35207 6885 35219 6888
rect 35161 6879 35219 6885
rect 35434 6876 35440 6888
rect 35492 6876 35498 6928
rect 3835 6820 4384 6848
rect 4433 6851 4491 6857
rect 3835 6817 3847 6820
rect 3789 6811 3847 6817
rect 4433 6817 4445 6851
rect 4479 6848 4491 6851
rect 4614 6848 4620 6860
rect 4479 6820 4620 6848
rect 4479 6817 4491 6820
rect 4433 6811 4491 6817
rect 4614 6808 4620 6820
rect 4672 6808 4678 6860
rect 33686 6808 33692 6860
rect 33744 6808 33750 6860
rect 33781 6851 33839 6857
rect 33781 6817 33793 6851
rect 33827 6848 33839 6851
rect 34238 6848 34244 6860
rect 33827 6820 34244 6848
rect 33827 6817 33839 6820
rect 33781 6811 33839 6817
rect 34238 6808 34244 6820
rect 34296 6808 34302 6860
rect 37182 6808 37188 6860
rect 37240 6808 37246 6860
rect 3073 6783 3131 6789
rect 3073 6749 3085 6783
rect 3119 6780 3131 6783
rect 5166 6780 5172 6792
rect 3119 6752 5172 6780
rect 3119 6749 3131 6752
rect 3073 6743 3131 6749
rect 5166 6740 5172 6752
rect 5224 6740 5230 6792
rect 33045 6783 33103 6789
rect 33045 6749 33057 6783
rect 33091 6780 33103 6783
rect 33704 6780 33732 6808
rect 33091 6752 33732 6780
rect 34517 6783 34575 6789
rect 33091 6749 33103 6752
rect 33045 6743 33103 6749
rect 34517 6749 34529 6783
rect 34563 6780 34575 6783
rect 35345 6783 35403 6789
rect 35345 6780 35357 6783
rect 34563 6752 35357 6780
rect 34563 6749 34575 6752
rect 34517 6743 34575 6749
rect 35345 6749 35357 6752
rect 35391 6749 35403 6783
rect 35345 6743 35403 6749
rect 35986 6740 35992 6792
rect 36044 6740 36050 6792
rect 36170 6740 36176 6792
rect 36228 6740 36234 6792
rect 4706 6712 4712 6724
rect 4540 6684 4712 6712
rect 1949 6647 2007 6653
rect 1949 6613 1961 6647
rect 1995 6644 2007 6647
rect 2774 6644 2780 6656
rect 1995 6616 2780 6644
rect 1995 6613 2007 6616
rect 1949 6607 2007 6613
rect 2774 6604 2780 6616
rect 2832 6604 2838 6656
rect 4540 6653 4568 6684
rect 4706 6672 4712 6684
rect 4764 6672 4770 6724
rect 4985 6715 5043 6721
rect 4985 6681 4997 6715
rect 5031 6712 5043 6715
rect 34793 6715 34851 6721
rect 34793 6712 34805 6715
rect 5031 6684 5396 6712
rect 5031 6681 5043 6684
rect 4985 6675 5043 6681
rect 5368 6653 5396 6684
rect 34532 6684 34805 6712
rect 34532 6656 34560 6684
rect 34793 6681 34805 6684
rect 34839 6681 34851 6715
rect 34793 6675 34851 6681
rect 4525 6647 4583 6653
rect 4525 6613 4537 6647
rect 4571 6613 4583 6647
rect 4525 6607 4583 6613
rect 5353 6647 5411 6653
rect 5353 6613 5365 6647
rect 5399 6644 5411 6647
rect 5442 6644 5448 6656
rect 5399 6616 5448 6644
rect 5399 6613 5411 6616
rect 5353 6607 5411 6613
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 32398 6604 32404 6656
rect 32456 6604 32462 6656
rect 33042 6604 33048 6656
rect 33100 6644 33106 6656
rect 33137 6647 33195 6653
rect 33137 6644 33149 6647
rect 33100 6616 33149 6644
rect 33100 6604 33106 6616
rect 33137 6613 33149 6616
rect 33183 6613 33195 6647
rect 33137 6607 33195 6613
rect 33873 6647 33931 6653
rect 33873 6613 33885 6647
rect 33919 6644 33931 6647
rect 34146 6644 34152 6656
rect 33919 6616 34152 6644
rect 33919 6613 33931 6616
rect 33873 6607 33931 6613
rect 34146 6604 34152 6616
rect 34204 6604 34210 6656
rect 34514 6604 34520 6656
rect 34572 6604 34578 6656
rect 35250 6604 35256 6656
rect 35308 6604 35314 6656
rect 1104 6554 37812 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 37812 6554
rect 1104 6480 37812 6502
rect 4249 6443 4307 6449
rect 4249 6409 4261 6443
rect 4295 6440 4307 6443
rect 4982 6440 4988 6452
rect 4295 6412 4988 6440
rect 4295 6409 4307 6412
rect 4249 6403 4307 6409
rect 4982 6400 4988 6412
rect 5040 6400 5046 6452
rect 33137 6443 33195 6449
rect 33137 6409 33149 6443
rect 33183 6440 33195 6443
rect 33502 6440 33508 6452
rect 33183 6412 33508 6440
rect 33183 6409 33195 6412
rect 33137 6403 33195 6409
rect 33502 6400 33508 6412
rect 33560 6400 33566 6452
rect 35250 6400 35256 6452
rect 35308 6400 35314 6452
rect 35986 6400 35992 6452
rect 36044 6440 36050 6452
rect 36817 6443 36875 6449
rect 36817 6440 36829 6443
rect 36044 6412 36829 6440
rect 36044 6400 36050 6412
rect 36817 6409 36829 6412
rect 36863 6409 36875 6443
rect 36817 6403 36875 6409
rect 1578 6332 1584 6384
rect 1636 6332 1642 6384
rect 35268 6372 35296 6400
rect 35682 6375 35740 6381
rect 35682 6372 35694 6375
rect 35268 6344 35694 6372
rect 35682 6341 35694 6344
rect 35728 6341 35740 6375
rect 35682 6335 35740 6341
rect 2590 6264 2596 6316
rect 2648 6264 2654 6316
rect 3418 6264 3424 6316
rect 3476 6264 3482 6316
rect 34054 6264 34060 6316
rect 34112 6304 34118 6316
rect 34112 6276 34836 6304
rect 34112 6264 34118 6276
rect 3602 6196 3608 6248
rect 3660 6196 3666 6248
rect 18506 6196 18512 6248
rect 18564 6236 18570 6248
rect 19242 6236 19248 6248
rect 18564 6208 19248 6236
rect 18564 6196 18570 6208
rect 19242 6196 19248 6208
rect 19300 6196 19306 6248
rect 32585 6239 32643 6245
rect 32585 6205 32597 6239
rect 32631 6205 32643 6239
rect 32585 6199 32643 6205
rect 33321 6239 33379 6245
rect 33321 6205 33333 6239
rect 33367 6236 33379 6239
rect 34146 6236 34152 6248
rect 33367 6208 34152 6236
rect 33367 6205 33379 6208
rect 33321 6199 33379 6205
rect 32600 6168 32628 6199
rect 34146 6196 34152 6208
rect 34204 6196 34210 6248
rect 34514 6196 34520 6248
rect 34572 6196 34578 6248
rect 34698 6196 34704 6248
rect 34756 6196 34762 6248
rect 34808 6236 34836 6276
rect 35250 6264 35256 6316
rect 35308 6264 35314 6316
rect 35342 6264 35348 6316
rect 35400 6304 35406 6316
rect 35437 6307 35495 6313
rect 35437 6304 35449 6307
rect 35400 6276 35449 6304
rect 35400 6264 35406 6276
rect 35437 6273 35449 6276
rect 35483 6273 35495 6307
rect 35437 6267 35495 6273
rect 35360 6236 35388 6264
rect 34808 6208 35388 6236
rect 32600 6140 34560 6168
rect 2866 6060 2872 6112
rect 2924 6060 2930 6112
rect 13998 6060 14004 6112
rect 14056 6060 14062 6112
rect 19153 6103 19211 6109
rect 19153 6069 19165 6103
rect 19199 6100 19211 6103
rect 20714 6100 20720 6112
rect 19199 6072 20720 6100
rect 19199 6069 19211 6072
rect 19153 6063 19211 6069
rect 20714 6060 20720 6072
rect 20772 6060 20778 6112
rect 33870 6060 33876 6112
rect 33928 6060 33934 6112
rect 34532 6100 34560 6140
rect 36170 6100 36176 6112
rect 34532 6072 36176 6100
rect 36170 6060 36176 6072
rect 36228 6060 36234 6112
rect 1104 6010 37812 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 37812 6010
rect 1104 5936 37812 5958
rect 2590 5856 2596 5908
rect 2648 5856 2654 5908
rect 3513 5899 3571 5905
rect 3513 5865 3525 5899
rect 3559 5896 3571 5899
rect 3602 5896 3608 5908
rect 3559 5868 3608 5896
rect 3559 5865 3571 5868
rect 3513 5859 3571 5865
rect 3602 5856 3608 5868
rect 3660 5856 3666 5908
rect 30190 5856 30196 5908
rect 30248 5856 30254 5908
rect 33870 5856 33876 5908
rect 33928 5896 33934 5908
rect 33928 5868 35848 5896
rect 33928 5856 33934 5868
rect 2409 5763 2467 5769
rect 2409 5729 2421 5763
rect 2455 5760 2467 5763
rect 2608 5760 2636 5856
rect 13538 5788 13544 5840
rect 13596 5788 13602 5840
rect 14458 5788 14464 5840
rect 14516 5788 14522 5840
rect 15381 5831 15439 5837
rect 15381 5797 15393 5831
rect 15427 5828 15439 5831
rect 16482 5828 16488 5840
rect 15427 5800 16488 5828
rect 15427 5797 15439 5800
rect 15381 5791 15439 5797
rect 16482 5788 16488 5800
rect 16540 5788 16546 5840
rect 34146 5788 34152 5840
rect 34204 5828 34210 5840
rect 35529 5831 35587 5837
rect 35529 5828 35541 5831
rect 34204 5800 35541 5828
rect 34204 5788 34210 5800
rect 35529 5797 35541 5800
rect 35575 5797 35587 5831
rect 35529 5791 35587 5797
rect 2455 5732 2636 5760
rect 2455 5729 2467 5732
rect 2409 5723 2467 5729
rect 2774 5720 2780 5772
rect 2832 5760 2838 5772
rect 2869 5763 2927 5769
rect 2869 5760 2881 5763
rect 2832 5732 2881 5760
rect 2832 5720 2838 5732
rect 2869 5729 2881 5732
rect 2915 5729 2927 5763
rect 2869 5723 2927 5729
rect 10888 5732 11652 5760
rect 10888 5704 10916 5732
rect 2685 5695 2743 5701
rect 2685 5661 2697 5695
rect 2731 5692 2743 5695
rect 3694 5692 3700 5704
rect 2731 5664 3700 5692
rect 2731 5661 2743 5664
rect 2685 5655 2743 5661
rect 3694 5652 3700 5664
rect 3752 5652 3758 5704
rect 10870 5652 10876 5704
rect 10928 5652 10934 5704
rect 10962 5652 10968 5704
rect 11020 5652 11026 5704
rect 11624 5692 11652 5732
rect 11882 5720 11888 5772
rect 11940 5760 11946 5772
rect 13449 5763 13507 5769
rect 13449 5760 13461 5763
rect 11940 5732 13461 5760
rect 11940 5720 11946 5732
rect 13449 5729 13461 5732
rect 13495 5729 13507 5763
rect 13449 5723 13507 5729
rect 31021 5763 31079 5769
rect 31021 5729 31033 5763
rect 31067 5760 31079 5763
rect 32398 5760 32404 5772
rect 31067 5732 32404 5760
rect 31067 5729 31079 5732
rect 31021 5723 31079 5729
rect 32398 5720 32404 5732
rect 32456 5720 32462 5772
rect 34057 5763 34115 5769
rect 34057 5729 34069 5763
rect 34103 5729 34115 5763
rect 34057 5723 34115 5729
rect 11624 5664 11928 5692
rect 9306 5584 9312 5636
rect 9364 5624 9370 5636
rect 11793 5627 11851 5633
rect 11793 5624 11805 5627
rect 9364 5596 11805 5624
rect 9364 5584 9370 5596
rect 11793 5593 11805 5596
rect 11839 5593 11851 5627
rect 11900 5624 11928 5664
rect 12158 5652 12164 5704
rect 12216 5692 12222 5704
rect 12345 5695 12403 5701
rect 12345 5692 12357 5695
rect 12216 5664 12357 5692
rect 12216 5652 12222 5664
rect 12345 5661 12357 5664
rect 12391 5661 12403 5695
rect 12345 5655 12403 5661
rect 13078 5652 13084 5704
rect 13136 5652 13142 5704
rect 31665 5695 31723 5701
rect 31665 5661 31677 5695
rect 31711 5692 31723 5695
rect 33045 5695 33103 5701
rect 31711 5664 32996 5692
rect 31711 5661 31723 5664
rect 31665 5655 31723 5661
rect 13909 5627 13967 5633
rect 13909 5624 13921 5627
rect 11900 5596 13921 5624
rect 11793 5587 11851 5593
rect 13909 5593 13921 5596
rect 13955 5624 13967 5627
rect 13998 5624 14004 5636
rect 13955 5596 14004 5624
rect 13955 5593 13967 5596
rect 13909 5587 13967 5593
rect 13998 5584 14004 5596
rect 14056 5624 14062 5636
rect 14093 5627 14151 5633
rect 14093 5624 14105 5627
rect 14056 5596 14105 5624
rect 14056 5584 14062 5596
rect 14093 5593 14105 5596
rect 14139 5624 14151 5627
rect 14829 5627 14887 5633
rect 14829 5624 14841 5627
rect 14139 5596 14841 5624
rect 14139 5593 14151 5596
rect 14093 5587 14151 5593
rect 14829 5593 14841 5596
rect 14875 5624 14887 5627
rect 15657 5627 15715 5633
rect 15657 5624 15669 5627
rect 14875 5596 15669 5624
rect 14875 5593 14887 5596
rect 14829 5587 14887 5593
rect 15657 5593 15669 5596
rect 15703 5624 15715 5627
rect 15746 5624 15752 5636
rect 15703 5596 15752 5624
rect 15703 5593 15715 5596
rect 15657 5587 15715 5593
rect 15746 5584 15752 5596
rect 15804 5624 15810 5636
rect 15933 5627 15991 5633
rect 15933 5624 15945 5627
rect 15804 5596 15945 5624
rect 15804 5584 15810 5596
rect 15933 5593 15945 5596
rect 15979 5593 15991 5627
rect 15933 5587 15991 5593
rect 31386 5584 31392 5636
rect 31444 5624 31450 5636
rect 32401 5627 32459 5633
rect 32401 5624 32413 5627
rect 31444 5596 32413 5624
rect 31444 5584 31450 5596
rect 32401 5593 32413 5596
rect 32447 5593 32459 5627
rect 32968 5624 32996 5664
rect 33045 5661 33057 5695
rect 33091 5692 33103 5695
rect 33870 5692 33876 5704
rect 33091 5664 33876 5692
rect 33091 5661 33103 5664
rect 33045 5655 33103 5661
rect 33870 5652 33876 5664
rect 33928 5652 33934 5704
rect 33962 5652 33968 5704
rect 34020 5652 34026 5704
rect 33980 5624 34008 5652
rect 32968 5596 34008 5624
rect 34072 5624 34100 5723
rect 34238 5720 34244 5772
rect 34296 5760 34302 5772
rect 35437 5763 35495 5769
rect 35437 5760 35449 5763
rect 34296 5732 35449 5760
rect 34296 5720 34302 5732
rect 35437 5729 35449 5732
rect 35483 5729 35495 5763
rect 35437 5723 35495 5729
rect 34517 5695 34575 5701
rect 34517 5661 34529 5695
rect 34563 5692 34575 5695
rect 34606 5692 34612 5704
rect 34563 5664 34612 5692
rect 34563 5661 34575 5664
rect 34517 5655 34575 5661
rect 34606 5652 34612 5664
rect 34664 5652 34670 5704
rect 35345 5695 35403 5701
rect 35345 5661 35357 5695
rect 35391 5692 35403 5695
rect 35710 5692 35716 5704
rect 35391 5664 35716 5692
rect 35391 5661 35403 5664
rect 35345 5655 35403 5661
rect 35710 5652 35716 5664
rect 35768 5652 35774 5704
rect 35820 5692 35848 5868
rect 36173 5695 36231 5701
rect 36173 5692 36185 5695
rect 35820 5664 36185 5692
rect 36173 5661 36185 5664
rect 36219 5661 36231 5695
rect 36173 5655 36231 5661
rect 34422 5624 34428 5636
rect 34072 5596 34428 5624
rect 32401 5587 32459 5593
rect 34422 5584 34428 5596
rect 34480 5584 34486 5636
rect 35618 5624 35624 5636
rect 34532 5596 35624 5624
rect 9950 5516 9956 5568
rect 10008 5556 10014 5568
rect 10689 5559 10747 5565
rect 10689 5556 10701 5559
rect 10008 5528 10701 5556
rect 10008 5516 10014 5528
rect 10689 5525 10701 5528
rect 10735 5556 10747 5559
rect 10870 5556 10876 5568
rect 10735 5528 10876 5556
rect 10735 5525 10747 5528
rect 10689 5519 10747 5525
rect 10870 5516 10876 5528
rect 10928 5516 10934 5568
rect 11238 5516 11244 5568
rect 11296 5556 11302 5568
rect 11609 5559 11667 5565
rect 11609 5556 11621 5559
rect 11296 5528 11621 5556
rect 11296 5516 11302 5528
rect 11609 5525 11621 5528
rect 11655 5525 11667 5559
rect 11609 5519 11667 5525
rect 11974 5516 11980 5568
rect 12032 5556 12038 5568
rect 12529 5559 12587 5565
rect 12529 5556 12541 5559
rect 12032 5528 12541 5556
rect 12032 5516 12038 5528
rect 12529 5525 12541 5528
rect 12575 5525 12587 5559
rect 12529 5519 12587 5525
rect 14366 5516 14372 5568
rect 14424 5556 14430 5568
rect 14553 5559 14611 5565
rect 14553 5556 14565 5559
rect 14424 5528 14565 5556
rect 14424 5516 14430 5528
rect 14553 5525 14565 5528
rect 14599 5525 14611 5559
rect 14553 5519 14611 5525
rect 15194 5516 15200 5568
rect 15252 5516 15258 5568
rect 29086 5516 29092 5568
rect 29144 5556 29150 5568
rect 29546 5556 29552 5568
rect 29144 5528 29552 5556
rect 29144 5516 29150 5528
rect 29546 5516 29552 5528
rect 29604 5556 29610 5568
rect 29733 5559 29791 5565
rect 29733 5556 29745 5559
rect 29604 5528 29745 5556
rect 29604 5516 29610 5528
rect 29733 5525 29745 5528
rect 29779 5525 29791 5559
rect 29733 5519 29791 5525
rect 31573 5559 31631 5565
rect 31573 5525 31585 5559
rect 31619 5556 31631 5559
rect 32214 5556 32220 5568
rect 31619 5528 32220 5556
rect 31619 5525 31631 5528
rect 31573 5519 31631 5525
rect 32214 5516 32220 5528
rect 32272 5516 32278 5568
rect 32309 5559 32367 5565
rect 32309 5525 32321 5559
rect 32355 5556 32367 5559
rect 34532 5556 34560 5596
rect 35618 5584 35624 5596
rect 35676 5584 35682 5636
rect 35894 5584 35900 5636
rect 35952 5584 35958 5636
rect 36538 5584 36544 5636
rect 36596 5584 36602 5636
rect 32355 5528 34560 5556
rect 34701 5559 34759 5565
rect 32355 5525 32367 5528
rect 32309 5519 32367 5525
rect 34701 5525 34713 5559
rect 34747 5556 34759 5559
rect 34882 5556 34888 5568
rect 34747 5528 34888 5556
rect 34747 5525 34759 5528
rect 34701 5519 34759 5525
rect 34882 5516 34888 5528
rect 34940 5516 34946 5568
rect 35912 5556 35940 5584
rect 37093 5559 37151 5565
rect 37093 5556 37105 5559
rect 35912 5528 37105 5556
rect 37093 5525 37105 5528
rect 37139 5525 37151 5559
rect 37093 5519 37151 5525
rect 1104 5466 37812 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 37812 5466
rect 1104 5392 37812 5414
rect 3510 5312 3516 5364
rect 3568 5312 3574 5364
rect 11701 5355 11759 5361
rect 11701 5321 11713 5355
rect 11747 5352 11759 5355
rect 13078 5352 13084 5364
rect 11747 5324 13084 5352
rect 11747 5321 11759 5324
rect 11701 5315 11759 5321
rect 3786 5284 3792 5296
rect 2700 5256 3792 5284
rect 2700 5225 2728 5256
rect 3786 5244 3792 5256
rect 3844 5244 3850 5296
rect 2685 5219 2743 5225
rect 2685 5185 2697 5219
rect 2731 5185 2743 5219
rect 2685 5179 2743 5185
rect 2866 5176 2872 5228
rect 2924 5176 2930 5228
rect 2409 5151 2467 5157
rect 2409 5117 2421 5151
rect 2455 5148 2467 5151
rect 2455 5120 2636 5148
rect 2455 5117 2467 5120
rect 2409 5111 2467 5117
rect 2608 5024 2636 5120
rect 9950 5108 9956 5160
rect 10008 5148 10014 5160
rect 10137 5151 10195 5157
rect 10137 5148 10149 5151
rect 10008 5120 10149 5148
rect 10008 5108 10014 5120
rect 10137 5117 10149 5120
rect 10183 5117 10195 5151
rect 11238 5148 11244 5160
rect 10137 5111 10195 5117
rect 10336 5120 11244 5148
rect 10336 5080 10364 5120
rect 11238 5108 11244 5120
rect 11296 5108 11302 5160
rect 9784 5052 10364 5080
rect 10505 5083 10563 5089
rect 9784 5024 9812 5052
rect 10505 5049 10517 5083
rect 10551 5080 10563 5083
rect 11716 5080 11744 5315
rect 13078 5312 13084 5324
rect 13136 5312 13142 5364
rect 14458 5312 14464 5364
rect 14516 5352 14522 5364
rect 14918 5352 14924 5364
rect 14516 5324 14924 5352
rect 14516 5312 14522 5324
rect 14918 5312 14924 5324
rect 14976 5312 14982 5364
rect 15746 5312 15752 5364
rect 15804 5352 15810 5364
rect 15841 5355 15899 5361
rect 15841 5352 15853 5355
rect 15804 5324 15853 5352
rect 15804 5312 15810 5324
rect 15841 5321 15853 5324
rect 15887 5321 15899 5355
rect 35253 5355 35311 5361
rect 35253 5352 35265 5355
rect 15841 5315 15899 5321
rect 31726 5324 34376 5352
rect 16114 5244 16120 5296
rect 16172 5284 16178 5296
rect 31726 5284 31754 5324
rect 34238 5284 34244 5296
rect 16172 5256 16574 5284
rect 16172 5244 16178 5256
rect 12345 5219 12403 5225
rect 12345 5185 12357 5219
rect 12391 5216 12403 5219
rect 13909 5219 13967 5225
rect 13909 5216 13921 5219
rect 12391 5188 13921 5216
rect 12391 5185 12403 5188
rect 12345 5179 12403 5185
rect 13909 5185 13921 5188
rect 13955 5185 13967 5219
rect 13909 5179 13967 5185
rect 13078 5108 13084 5160
rect 13136 5108 13142 5160
rect 13722 5108 13728 5160
rect 13780 5108 13786 5160
rect 14458 5108 14464 5160
rect 14516 5108 14522 5160
rect 15470 5108 15476 5160
rect 15528 5108 15534 5160
rect 16546 5148 16574 5256
rect 26206 5256 31754 5284
rect 33040 5256 34244 5284
rect 25958 5176 25964 5228
rect 26016 5216 26022 5228
rect 26206 5216 26234 5256
rect 26016 5188 26234 5216
rect 26016 5176 26022 5188
rect 31386 5176 31392 5228
rect 31444 5176 31450 5228
rect 33040 5225 33068 5256
rect 34238 5244 34244 5256
rect 34296 5244 34302 5296
rect 34348 5225 34376 5324
rect 34532 5324 35265 5352
rect 34532 5296 34560 5324
rect 35253 5321 35265 5324
rect 35299 5352 35311 5355
rect 35894 5352 35900 5364
rect 35299 5324 35900 5352
rect 35299 5321 35311 5324
rect 35253 5315 35311 5321
rect 35894 5312 35900 5324
rect 35952 5312 35958 5364
rect 34514 5244 34520 5296
rect 34572 5244 34578 5296
rect 34606 5244 34612 5296
rect 34664 5284 34670 5296
rect 34701 5287 34759 5293
rect 34701 5284 34713 5287
rect 34664 5256 34713 5284
rect 34664 5244 34670 5256
rect 34701 5253 34713 5256
rect 34747 5253 34759 5287
rect 34701 5247 34759 5253
rect 33036 5219 33094 5225
rect 33036 5185 33048 5219
rect 33082 5185 33094 5219
rect 33036 5179 33094 5185
rect 34333 5219 34391 5225
rect 34333 5185 34345 5219
rect 34379 5185 34391 5219
rect 35805 5219 35863 5225
rect 35805 5216 35817 5219
rect 34333 5179 34391 5185
rect 34900 5188 35817 5216
rect 16945 5151 17003 5157
rect 16945 5148 16957 5151
rect 16546 5120 16957 5148
rect 16945 5117 16957 5120
rect 16991 5148 17003 5151
rect 17129 5151 17187 5157
rect 17129 5148 17141 5151
rect 16991 5120 17141 5148
rect 16991 5117 17003 5120
rect 16945 5111 17003 5117
rect 17129 5117 17141 5120
rect 17175 5148 17187 5151
rect 17175 5120 18644 5148
rect 17175 5117 17187 5120
rect 17129 5111 17187 5117
rect 10551 5052 11744 5080
rect 10551 5049 10563 5052
rect 10505 5043 10563 5049
rect 12250 5040 12256 5092
rect 12308 5080 12314 5092
rect 13173 5083 13231 5089
rect 13173 5080 13185 5083
rect 12308 5052 13185 5080
rect 12308 5040 12314 5052
rect 13173 5049 13185 5052
rect 13219 5049 13231 5083
rect 13173 5043 13231 5049
rect 17497 5083 17555 5089
rect 17497 5049 17509 5083
rect 17543 5080 17555 5083
rect 18506 5080 18512 5092
rect 17543 5052 18512 5080
rect 17543 5049 17555 5052
rect 17497 5043 17555 5049
rect 18506 5040 18512 5052
rect 18564 5040 18570 5092
rect 2590 4972 2596 5024
rect 2648 4972 2654 5024
rect 9766 4972 9772 5024
rect 9824 4972 9830 5024
rect 9950 4972 9956 5024
rect 10008 4972 10014 5024
rect 10594 4972 10600 5024
rect 10652 4972 10658 5024
rect 10686 4972 10692 5024
rect 10744 4972 10750 5024
rect 12437 5015 12495 5021
rect 12437 4981 12449 5015
rect 12483 5012 12495 5015
rect 12618 5012 12624 5024
rect 12483 4984 12624 5012
rect 12483 4981 12495 4984
rect 12437 4975 12495 4981
rect 12618 4972 12624 4984
rect 12676 4972 12682 5024
rect 17589 5015 17647 5021
rect 17589 4981 17601 5015
rect 17635 5012 17647 5015
rect 17678 5012 17684 5024
rect 17635 4984 17684 5012
rect 17635 4981 17647 4984
rect 17589 4975 17647 4981
rect 17678 4972 17684 4984
rect 17736 4972 17742 5024
rect 17957 5015 18015 5021
rect 17957 4981 17969 5015
rect 18003 5012 18015 5015
rect 18616 5012 18644 5120
rect 27154 5108 27160 5160
rect 27212 5108 27218 5160
rect 28166 5108 28172 5160
rect 28224 5148 28230 5160
rect 28905 5151 28963 5157
rect 28905 5148 28917 5151
rect 28224 5120 28917 5148
rect 28224 5108 28230 5120
rect 28905 5117 28917 5120
rect 28951 5117 28963 5151
rect 28905 5111 28963 5117
rect 29454 5108 29460 5160
rect 29512 5108 29518 5160
rect 29546 5108 29552 5160
rect 29604 5148 29610 5160
rect 29641 5151 29699 5157
rect 29641 5148 29653 5151
rect 29604 5120 29653 5148
rect 29604 5108 29610 5120
rect 29641 5117 29653 5120
rect 29687 5117 29699 5151
rect 29641 5111 29699 5117
rect 30190 5108 30196 5160
rect 30248 5108 30254 5160
rect 30469 5151 30527 5157
rect 30469 5117 30481 5151
rect 30515 5148 30527 5151
rect 30650 5148 30656 5160
rect 30515 5120 30656 5148
rect 30515 5117 30527 5120
rect 30469 5111 30527 5117
rect 30650 5108 30656 5120
rect 30708 5108 30714 5160
rect 32217 5151 32275 5157
rect 32217 5117 32229 5151
rect 32263 5117 32275 5151
rect 32217 5111 32275 5117
rect 28813 5083 28871 5089
rect 28813 5049 28825 5083
rect 28859 5080 28871 5083
rect 29362 5080 29368 5092
rect 28859 5052 29368 5080
rect 28859 5049 28871 5052
rect 28813 5043 28871 5049
rect 29362 5040 29368 5052
rect 29420 5040 29426 5092
rect 30208 5080 30236 5108
rect 31846 5080 31852 5092
rect 30208 5052 31852 5080
rect 31846 5040 31852 5052
rect 31904 5080 31910 5092
rect 32232 5080 32260 5111
rect 32766 5108 32772 5160
rect 32824 5108 32830 5160
rect 34790 5108 34796 5160
rect 34848 5108 34854 5160
rect 31904 5052 32260 5080
rect 31904 5040 31910 5052
rect 32398 5040 32404 5092
rect 32456 5080 32462 5092
rect 32493 5083 32551 5089
rect 32493 5080 32505 5083
rect 32456 5052 32505 5080
rect 32456 5040 32462 5052
rect 32493 5049 32505 5052
rect 32539 5049 32551 5083
rect 34149 5083 34207 5089
rect 32493 5043 32551 5049
rect 32600 5052 32812 5080
rect 19334 5012 19340 5024
rect 18003 4984 19340 5012
rect 18003 4981 18015 4984
rect 17957 4975 18015 4981
rect 19334 4972 19340 4984
rect 19392 4972 19398 5024
rect 26234 4972 26240 5024
rect 26292 5012 26298 5024
rect 26329 5015 26387 5021
rect 26329 5012 26341 5015
rect 26292 4984 26341 5012
rect 26292 4972 26298 4984
rect 26329 4981 26341 4984
rect 26375 4981 26387 5015
rect 26329 4975 26387 4981
rect 27798 4972 27804 5024
rect 27856 4972 27862 5024
rect 30282 4972 30288 5024
rect 30340 4972 30346 5024
rect 31021 5015 31079 5021
rect 31021 4981 31033 5015
rect 31067 5012 31079 5015
rect 31754 5012 31760 5024
rect 31067 4984 31760 5012
rect 31067 4981 31079 4984
rect 31021 4975 31079 4981
rect 31754 4972 31760 4984
rect 31812 4972 31818 5024
rect 31938 4972 31944 5024
rect 31996 4972 32002 5024
rect 32214 4972 32220 5024
rect 32272 5012 32278 5024
rect 32600 5012 32628 5052
rect 32272 4984 32628 5012
rect 32272 4972 32278 4984
rect 32674 4972 32680 5024
rect 32732 4972 32738 5024
rect 32784 5012 32812 5052
rect 34149 5049 34161 5083
rect 34195 5080 34207 5083
rect 34808 5080 34836 5108
rect 34195 5052 34836 5080
rect 34195 5049 34207 5052
rect 34149 5043 34207 5049
rect 34900 5012 34928 5188
rect 35805 5185 35817 5188
rect 35851 5185 35863 5219
rect 35805 5179 35863 5185
rect 36078 5108 36084 5160
rect 36136 5108 36142 5160
rect 32784 4984 34928 5012
rect 36817 5015 36875 5021
rect 36817 4981 36829 5015
rect 36863 5012 36875 5015
rect 37090 5012 37096 5024
rect 36863 4984 37096 5012
rect 36863 4981 36875 4984
rect 36817 4975 36875 4981
rect 37090 4972 37096 4984
rect 37148 4972 37154 5024
rect 1104 4922 37812 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 37812 4922
rect 1104 4848 37812 4870
rect 10597 4811 10655 4817
rect 10597 4777 10609 4811
rect 10643 4808 10655 4811
rect 10962 4808 10968 4820
rect 10643 4780 10968 4808
rect 10643 4777 10655 4780
rect 10597 4771 10655 4777
rect 10962 4768 10968 4780
rect 11020 4768 11026 4820
rect 13078 4768 13084 4820
rect 13136 4808 13142 4820
rect 13265 4811 13323 4817
rect 13265 4808 13277 4811
rect 13136 4780 13277 4808
rect 13136 4768 13142 4780
rect 13265 4777 13277 4780
rect 13311 4777 13323 4811
rect 13265 4771 13323 4777
rect 29181 4811 29239 4817
rect 29181 4777 29193 4811
rect 29227 4808 29239 4811
rect 29454 4808 29460 4820
rect 29227 4780 29460 4808
rect 29227 4777 29239 4780
rect 29181 4771 29239 4777
rect 29454 4768 29460 4780
rect 29512 4768 29518 4820
rect 33870 4768 33876 4820
rect 33928 4808 33934 4820
rect 34701 4811 34759 4817
rect 34701 4808 34713 4811
rect 33928 4780 34713 4808
rect 33928 4768 33934 4780
rect 34701 4777 34713 4780
rect 34747 4777 34759 4811
rect 34701 4771 34759 4777
rect 36078 4768 36084 4820
rect 36136 4768 36142 4820
rect 9766 4700 9772 4752
rect 9824 4700 9830 4752
rect 10689 4743 10747 4749
rect 10689 4709 10701 4743
rect 10735 4709 10747 4743
rect 10689 4703 10747 4709
rect 18785 4743 18843 4749
rect 18785 4709 18797 4743
rect 18831 4740 18843 4743
rect 19242 4740 19248 4752
rect 18831 4712 19248 4740
rect 18831 4709 18843 4712
rect 18785 4703 18843 4709
rect 934 4632 940 4684
rect 992 4672 998 4684
rect 1581 4675 1639 4681
rect 1581 4672 1593 4675
rect 992 4644 1593 4672
rect 992 4632 998 4644
rect 1581 4641 1593 4644
rect 1627 4641 1639 4675
rect 1581 4635 1639 4641
rect 10045 4675 10103 4681
rect 10045 4641 10057 4675
rect 10091 4672 10103 4675
rect 10704 4672 10732 4703
rect 19242 4700 19248 4712
rect 19300 4700 19306 4752
rect 26142 4700 26148 4752
rect 26200 4700 26206 4752
rect 30009 4743 30067 4749
rect 30009 4709 30021 4743
rect 30055 4740 30067 4743
rect 31386 4740 31392 4752
rect 30055 4712 31392 4740
rect 30055 4709 30067 4712
rect 30009 4703 30067 4709
rect 31386 4700 31392 4712
rect 31444 4700 31450 4752
rect 36096 4740 36124 4768
rect 31726 4712 36124 4740
rect 10091 4644 10732 4672
rect 10091 4641 10103 4644
rect 10045 4635 10103 4641
rect 12066 4632 12072 4684
rect 12124 4632 12130 4684
rect 13538 4672 13544 4684
rect 12452 4644 13544 4672
rect 12452 4616 12480 4644
rect 13538 4632 13544 4644
rect 13596 4672 13602 4684
rect 14645 4675 14703 4681
rect 14645 4672 14657 4675
rect 13596 4644 14657 4672
rect 13596 4632 13602 4644
rect 14645 4641 14657 4644
rect 14691 4641 14703 4675
rect 14645 4635 14703 4641
rect 14918 4632 14924 4684
rect 14976 4672 14982 4684
rect 15013 4675 15071 4681
rect 15013 4672 15025 4675
rect 14976 4644 15025 4672
rect 14976 4632 14982 4644
rect 15013 4641 15025 4644
rect 15059 4641 15071 4675
rect 15013 4635 15071 4641
rect 16666 4632 16672 4684
rect 16724 4632 16730 4684
rect 2590 4564 2596 4616
rect 2648 4564 2654 4616
rect 10594 4564 10600 4616
rect 10652 4564 10658 4616
rect 12434 4564 12440 4616
rect 12492 4564 12498 4616
rect 13170 4564 13176 4616
rect 13228 4564 13234 4616
rect 13814 4564 13820 4616
rect 13872 4564 13878 4616
rect 16482 4564 16488 4616
rect 16540 4564 16546 4616
rect 18230 4564 18236 4616
rect 18288 4564 18294 4616
rect 5442 4496 5448 4548
rect 5500 4536 5506 4548
rect 9401 4539 9459 4545
rect 9401 4536 9413 4539
rect 5500 4508 9413 4536
rect 5500 4496 5506 4508
rect 9401 4505 9413 4508
rect 9447 4536 9459 4539
rect 9950 4536 9956 4548
rect 9447 4508 9956 4536
rect 9447 4505 9459 4508
rect 9401 4499 9459 4505
rect 9950 4496 9956 4508
rect 10008 4496 10014 4548
rect 10612 4536 10640 4564
rect 11802 4539 11860 4545
rect 11802 4536 11814 4539
rect 10612 4508 11814 4536
rect 11802 4505 11814 4508
rect 11848 4505 11860 4539
rect 11802 4499 11860 4505
rect 18417 4539 18475 4545
rect 18417 4505 18429 4539
rect 18463 4536 18475 4539
rect 25501 4539 25559 4545
rect 18463 4508 19380 4536
rect 18463 4505 18475 4508
rect 18417 4499 18475 4505
rect 19352 4480 19380 4508
rect 25501 4505 25513 4539
rect 25547 4536 25559 4539
rect 25777 4539 25835 4545
rect 25777 4536 25789 4539
rect 25547 4508 25789 4536
rect 25547 4505 25559 4508
rect 25501 4499 25559 4505
rect 25777 4505 25789 4508
rect 25823 4505 25835 4539
rect 26160 4536 26188 4700
rect 26237 4675 26295 4681
rect 26237 4641 26249 4675
rect 26283 4672 26295 4675
rect 27706 4672 27712 4684
rect 26283 4644 27712 4672
rect 26283 4641 26295 4644
rect 26237 4635 26295 4641
rect 27706 4632 27712 4644
rect 27764 4632 27770 4684
rect 27893 4675 27951 4681
rect 27893 4641 27905 4675
rect 27939 4672 27951 4675
rect 27939 4644 28764 4672
rect 27939 4641 27951 4644
rect 27893 4635 27951 4641
rect 28736 4616 28764 4644
rect 29454 4632 29460 4684
rect 29512 4672 29518 4684
rect 29641 4675 29699 4681
rect 29641 4672 29653 4675
rect 29512 4644 29653 4672
rect 29512 4632 29518 4644
rect 29641 4641 29653 4644
rect 29687 4672 29699 4675
rect 30190 4672 30196 4684
rect 29687 4644 30196 4672
rect 29687 4641 29699 4644
rect 29641 4635 29699 4641
rect 30190 4632 30196 4644
rect 30248 4632 30254 4684
rect 31110 4632 31116 4684
rect 31168 4632 31174 4684
rect 31726 4672 31754 4712
rect 31588 4644 31754 4672
rect 32585 4675 32643 4681
rect 26326 4564 26332 4616
rect 26384 4564 26390 4616
rect 27617 4607 27675 4613
rect 27617 4573 27629 4607
rect 27663 4573 27675 4607
rect 27617 4567 27675 4573
rect 27632 4536 27660 4567
rect 28626 4564 28632 4616
rect 28684 4564 28690 4616
rect 28718 4564 28724 4616
rect 28776 4564 28782 4616
rect 31588 4613 31616 4644
rect 32585 4641 32597 4675
rect 32631 4672 32643 4675
rect 33870 4672 33876 4684
rect 32631 4644 33876 4672
rect 32631 4641 32643 4644
rect 32585 4635 32643 4641
rect 33870 4632 33876 4644
rect 33928 4632 33934 4684
rect 34054 4632 34060 4684
rect 34112 4632 34118 4684
rect 35802 4672 35808 4684
rect 35452 4644 35808 4672
rect 31573 4607 31631 4613
rect 31573 4573 31585 4607
rect 31619 4573 31631 4607
rect 31573 4567 31631 4573
rect 33045 4607 33103 4613
rect 33045 4573 33057 4607
rect 33091 4604 33103 4607
rect 33502 4604 33508 4616
rect 33091 4576 33508 4604
rect 33091 4573 33103 4576
rect 33045 4567 33103 4573
rect 33502 4564 33508 4576
rect 33560 4564 33566 4616
rect 34425 4607 34483 4613
rect 34425 4573 34437 4607
rect 34471 4604 34483 4607
rect 34790 4604 34796 4616
rect 34471 4576 34796 4604
rect 34471 4573 34483 4576
rect 34425 4567 34483 4573
rect 34790 4564 34796 4576
rect 34848 4564 34854 4616
rect 35452 4613 35480 4644
rect 35802 4632 35808 4644
rect 35860 4672 35866 4684
rect 37185 4675 37243 4681
rect 35860 4644 37136 4672
rect 35860 4632 35866 4644
rect 37108 4616 37136 4644
rect 37185 4641 37197 4675
rect 37231 4672 37243 4675
rect 37642 4672 37648 4684
rect 37231 4644 37648 4672
rect 37231 4641 37243 4644
rect 37185 4635 37243 4641
rect 37642 4632 37648 4644
rect 37700 4632 37706 4684
rect 35253 4607 35311 4613
rect 35253 4573 35265 4607
rect 35299 4573 35311 4607
rect 35253 4567 35311 4573
rect 35437 4607 35495 4613
rect 35437 4573 35449 4607
rect 35483 4573 35495 4607
rect 35437 4567 35495 4573
rect 36265 4607 36323 4613
rect 36265 4573 36277 4607
rect 36311 4604 36323 4607
rect 36538 4604 36544 4616
rect 36311 4576 36544 4604
rect 36311 4573 36323 4576
rect 36265 4567 36323 4573
rect 26160 4508 27660 4536
rect 25777 4499 25835 4505
rect 9861 4471 9919 4477
rect 9861 4437 9873 4471
rect 9907 4468 9919 4471
rect 11054 4468 11060 4480
rect 9907 4440 11060 4468
rect 9907 4437 9919 4440
rect 9861 4431 9919 4437
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 12526 4428 12532 4480
rect 12584 4428 12590 4480
rect 14090 4428 14096 4480
rect 14148 4428 14154 4480
rect 15654 4428 15660 4480
rect 15712 4428 15718 4480
rect 15838 4428 15844 4480
rect 15896 4428 15902 4480
rect 17218 4428 17224 4480
rect 17276 4428 17282 4480
rect 17310 4428 17316 4480
rect 17368 4468 17374 4480
rect 17681 4471 17739 4477
rect 17681 4468 17693 4471
rect 17368 4440 17693 4468
rect 17368 4428 17374 4440
rect 17681 4437 17693 4440
rect 17727 4437 17739 4471
rect 17681 4431 17739 4437
rect 18782 4428 18788 4480
rect 18840 4468 18846 4480
rect 18877 4471 18935 4477
rect 18877 4468 18889 4471
rect 18840 4440 18889 4468
rect 18840 4428 18846 4440
rect 18877 4437 18889 4440
rect 18923 4437 18935 4471
rect 18877 4431 18935 4437
rect 19334 4428 19340 4480
rect 19392 4468 19398 4480
rect 19429 4471 19487 4477
rect 19429 4468 19441 4471
rect 19392 4440 19441 4468
rect 19392 4428 19398 4440
rect 19429 4437 19441 4440
rect 19475 4437 19487 4471
rect 25792 4468 25820 4499
rect 33686 4496 33692 4548
rect 33744 4536 33750 4548
rect 35268 4536 35296 4567
rect 36538 4564 36544 4576
rect 36596 4564 36602 4616
rect 37090 4564 37096 4616
rect 37148 4564 37154 4616
rect 33744 4508 35296 4536
rect 35713 4539 35771 4545
rect 33744 4496 33750 4508
rect 35713 4505 35725 4539
rect 35759 4505 35771 4539
rect 35713 4499 35771 4505
rect 26234 4468 26240 4480
rect 25792 4440 26240 4468
rect 19429 4431 19487 4437
rect 26234 4428 26240 4440
rect 26292 4428 26298 4480
rect 26694 4428 26700 4480
rect 26752 4468 26758 4480
rect 26973 4471 27031 4477
rect 26973 4468 26985 4471
rect 26752 4440 26985 4468
rect 26752 4428 26758 4440
rect 26973 4437 26985 4440
rect 27019 4437 27031 4471
rect 26973 4431 27031 4437
rect 27062 4428 27068 4480
rect 27120 4428 27126 4480
rect 28442 4428 28448 4480
rect 28500 4428 28506 4480
rect 30098 4428 30104 4480
rect 30156 4428 30162 4480
rect 34514 4428 34520 4480
rect 34572 4468 34578 4480
rect 35728 4468 35756 4499
rect 34572 4440 35756 4468
rect 34572 4428 34578 4440
rect 1104 4378 37812 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 37812 4378
rect 1104 4304 37812 4326
rect 12066 4224 12072 4276
rect 12124 4224 12130 4276
rect 13170 4224 13176 4276
rect 13228 4264 13234 4276
rect 13265 4267 13323 4273
rect 13265 4264 13277 4267
rect 13228 4236 13277 4264
rect 13228 4224 13234 4236
rect 13265 4233 13277 4236
rect 13311 4233 13323 4267
rect 26970 4264 26976 4276
rect 13265 4227 13323 4233
rect 26252 4236 26976 4264
rect 12084 4196 12112 4224
rect 26252 4208 26280 4236
rect 26970 4224 26976 4236
rect 27028 4224 27034 4276
rect 28626 4224 28632 4276
rect 28684 4264 28690 4276
rect 28905 4267 28963 4273
rect 28905 4264 28917 4267
rect 28684 4236 28917 4264
rect 28684 4224 28690 4236
rect 28905 4233 28917 4236
rect 28951 4233 28963 4267
rect 28905 4227 28963 4233
rect 31110 4224 31116 4276
rect 31168 4264 31174 4276
rect 36998 4264 37004 4276
rect 31168 4236 37004 4264
rect 31168 4224 31174 4236
rect 36998 4224 37004 4236
rect 37056 4224 37062 4276
rect 25317 4199 25375 4205
rect 11808 4168 12388 4196
rect 2685 4131 2743 4137
rect 2685 4097 2697 4131
rect 2731 4128 2743 4131
rect 2958 4128 2964 4140
rect 2731 4100 2964 4128
rect 2731 4097 2743 4100
rect 2685 4091 2743 4097
rect 2958 4088 2964 4100
rect 3016 4088 3022 4140
rect 9306 4088 9312 4140
rect 9364 4088 9370 4140
rect 10134 4088 10140 4140
rect 10192 4088 10198 4140
rect 11808 4137 11836 4168
rect 11793 4131 11851 4137
rect 11793 4097 11805 4131
rect 11839 4097 11851 4131
rect 11793 4091 11851 4097
rect 11882 4088 11888 4140
rect 11940 4128 11946 4140
rect 12049 4131 12107 4137
rect 12049 4128 12061 4131
rect 11940 4100 12061 4128
rect 11940 4088 11946 4100
rect 12049 4097 12061 4100
rect 12095 4097 12107 4131
rect 12360 4128 12388 4168
rect 14292 4168 14596 4196
rect 14292 4128 14320 4168
rect 12360 4100 14320 4128
rect 12049 4091 12107 4097
rect 14366 4088 14372 4140
rect 14424 4137 14430 4140
rect 14424 4128 14436 4137
rect 14568 4128 14596 4168
rect 25317 4165 25329 4199
rect 25363 4196 25375 4199
rect 26234 4196 26240 4208
rect 25363 4168 26240 4196
rect 25363 4165 25375 4168
rect 25317 4159 25375 4165
rect 26234 4156 26240 4168
rect 26292 4156 26298 4208
rect 26712 4168 28764 4196
rect 14642 4128 14648 4140
rect 14424 4100 14469 4128
rect 14568 4100 14648 4128
rect 14424 4091 14436 4100
rect 14424 4088 14430 4091
rect 14642 4088 14648 4100
rect 14700 4088 14706 4140
rect 15286 4088 15292 4140
rect 15344 4088 15350 4140
rect 17589 4131 17647 4137
rect 17589 4097 17601 4131
rect 17635 4128 17647 4131
rect 17773 4131 17831 4137
rect 17773 4128 17785 4131
rect 17635 4100 17785 4128
rect 17635 4097 17647 4100
rect 17589 4091 17647 4097
rect 17773 4097 17785 4100
rect 17819 4097 17831 4131
rect 17773 4091 17831 4097
rect 2409 4063 2467 4069
rect 2409 4029 2421 4063
rect 2455 4060 2467 4063
rect 2455 4032 2636 4060
rect 2455 4029 2467 4032
rect 2409 4023 2467 4029
rect 2608 3936 2636 4032
rect 10594 4020 10600 4072
rect 10652 4020 10658 4072
rect 13630 4020 13636 4072
rect 13688 4020 13694 4072
rect 15010 4020 15016 4072
rect 15068 4060 15074 4072
rect 15565 4063 15623 4069
rect 15565 4060 15577 4063
rect 15068 4032 15577 4060
rect 15068 4020 15074 4032
rect 15565 4029 15577 4032
rect 15611 4029 15623 4063
rect 15565 4023 15623 4029
rect 16942 4020 16948 4072
rect 17000 4020 17006 4072
rect 18046 4020 18052 4072
rect 18104 4020 18110 4072
rect 19150 4020 19156 4072
rect 19208 4020 19214 4072
rect 25314 4020 25320 4072
rect 25372 4060 25378 4072
rect 25593 4063 25651 4069
rect 25593 4060 25605 4063
rect 25372 4032 25605 4060
rect 25372 4020 25378 4032
rect 25593 4029 25605 4032
rect 25639 4029 25651 4063
rect 25593 4023 25651 4029
rect 13648 3992 13676 4020
rect 12728 3964 13676 3992
rect 25041 3995 25099 4001
rect 2590 3884 2596 3936
rect 2648 3884 2654 3936
rect 9861 3927 9919 3933
rect 9861 3893 9873 3927
rect 9907 3924 9919 3927
rect 12728 3924 12756 3964
rect 25041 3961 25053 3995
rect 25087 3992 25099 3995
rect 26712 3992 26740 4168
rect 28736 4140 28764 4168
rect 32766 4156 32772 4208
rect 32824 4196 32830 4208
rect 34146 4196 34152 4208
rect 32824 4168 34152 4196
rect 32824 4156 32830 4168
rect 26789 4131 26847 4137
rect 26789 4097 26801 4131
rect 26835 4128 26847 4131
rect 26835 4100 26924 4128
rect 26835 4097 26847 4100
rect 26789 4091 26847 4097
rect 25087 3964 26740 3992
rect 25087 3961 25099 3964
rect 25041 3955 25099 3961
rect 26896 3936 26924 4100
rect 26970 4088 26976 4140
rect 27028 4088 27034 4140
rect 27781 4131 27839 4137
rect 27781 4128 27793 4131
rect 27448 4100 27793 4128
rect 27448 4069 27476 4100
rect 27781 4097 27793 4100
rect 27827 4097 27839 4131
rect 27781 4091 27839 4097
rect 28718 4088 28724 4140
rect 28776 4088 28782 4140
rect 30466 4088 30472 4140
rect 30524 4088 30530 4140
rect 31941 4131 31999 4137
rect 31941 4097 31953 4131
rect 31987 4128 31999 4131
rect 32490 4128 32496 4140
rect 31987 4100 32496 4128
rect 31987 4097 31999 4100
rect 31941 4091 31999 4097
rect 32490 4088 32496 4100
rect 32548 4088 32554 4140
rect 33152 4137 33180 4168
rect 34146 4156 34152 4168
rect 34204 4156 34210 4208
rect 34790 4156 34796 4208
rect 34848 4196 34854 4208
rect 35345 4199 35403 4205
rect 35345 4196 35357 4199
rect 34848 4168 35357 4196
rect 34848 4156 34854 4168
rect 35345 4165 35357 4168
rect 35391 4165 35403 4199
rect 35345 4159 35403 4165
rect 33137 4131 33195 4137
rect 33137 4097 33149 4131
rect 33183 4097 33195 4131
rect 33137 4091 33195 4097
rect 33404 4131 33462 4137
rect 33404 4097 33416 4131
rect 33450 4128 33462 4131
rect 34238 4128 34244 4140
rect 33450 4100 34244 4128
rect 33450 4097 33462 4100
rect 33404 4091 33462 4097
rect 34238 4088 34244 4100
rect 34296 4088 34302 4140
rect 34514 4088 34520 4140
rect 34572 4088 34578 4140
rect 35434 4088 35440 4140
rect 35492 4088 35498 4140
rect 35894 4088 35900 4140
rect 35952 4088 35958 4140
rect 36630 4088 36636 4140
rect 36688 4088 36694 4140
rect 27433 4063 27491 4069
rect 27433 4029 27445 4063
rect 27479 4029 27491 4063
rect 27433 4023 27491 4029
rect 27522 4020 27528 4072
rect 27580 4020 27586 4072
rect 28626 4020 28632 4072
rect 28684 4060 28690 4072
rect 29273 4063 29331 4069
rect 29273 4060 29285 4063
rect 28684 4032 29285 4060
rect 28684 4020 28690 4032
rect 29273 4029 29285 4032
rect 29319 4029 29331 4063
rect 29273 4023 29331 4029
rect 29730 4020 29736 4072
rect 29788 4060 29794 4072
rect 30745 4063 30803 4069
rect 30745 4060 30757 4063
rect 29788 4032 30757 4060
rect 29788 4020 29794 4032
rect 30745 4029 30757 4032
rect 30791 4029 30803 4063
rect 30745 4023 30803 4029
rect 32122 4020 32128 4072
rect 32180 4020 32186 4072
rect 27341 3995 27399 4001
rect 27341 3961 27353 3995
rect 27387 3961 27399 3995
rect 27341 3955 27399 3961
rect 9907 3896 12756 3924
rect 13173 3927 13231 3933
rect 9907 3893 9919 3896
rect 9861 3887 9919 3893
rect 13173 3893 13185 3927
rect 13219 3924 13231 3927
rect 14458 3924 14464 3936
rect 13219 3896 14464 3924
rect 13219 3893 13231 3896
rect 13173 3887 13231 3893
rect 14458 3884 14464 3896
rect 14516 3884 14522 3936
rect 19797 3927 19855 3933
rect 19797 3893 19809 3927
rect 19843 3924 19855 3927
rect 19978 3924 19984 3936
rect 19843 3896 19984 3924
rect 19843 3893 19855 3896
rect 19797 3887 19855 3893
rect 19978 3884 19984 3896
rect 20036 3884 20042 3936
rect 24854 3884 24860 3936
rect 24912 3884 24918 3936
rect 26878 3884 26884 3936
rect 26936 3884 26942 3936
rect 27356 3924 27384 3955
rect 30650 3952 30656 4004
rect 30708 3952 30714 4004
rect 34532 3992 34560 4088
rect 35452 4060 35480 4088
rect 36081 4063 36139 4069
rect 36081 4060 36093 4063
rect 35452 4032 36093 4060
rect 36081 4029 36093 4032
rect 36127 4029 36139 4063
rect 36081 4023 36139 4029
rect 34793 3995 34851 4001
rect 34793 3992 34805 3995
rect 34440 3964 34805 3992
rect 30668 3924 30696 3952
rect 34440 3936 34468 3964
rect 34793 3961 34805 3964
rect 34839 3961 34851 3995
rect 34793 3955 34851 3961
rect 27356 3896 30696 3924
rect 32769 3927 32827 3933
rect 32769 3893 32781 3927
rect 32815 3924 32827 3927
rect 33134 3924 33140 3936
rect 32815 3896 33140 3924
rect 32815 3893 32827 3896
rect 32769 3887 32827 3893
rect 33134 3884 33140 3896
rect 33192 3884 33198 3936
rect 34422 3884 34428 3936
rect 34480 3884 34486 3936
rect 34517 3927 34575 3933
rect 34517 3893 34529 3927
rect 34563 3924 34575 3927
rect 34606 3924 34612 3936
rect 34563 3896 34612 3924
rect 34563 3893 34575 3896
rect 34517 3887 34575 3893
rect 34606 3884 34612 3896
rect 34664 3884 34670 3936
rect 36906 3884 36912 3936
rect 36964 3924 36970 3936
rect 37001 3927 37059 3933
rect 37001 3924 37013 3927
rect 36964 3896 37013 3924
rect 36964 3884 36970 3896
rect 37001 3893 37013 3896
rect 37047 3893 37059 3927
rect 37001 3887 37059 3893
rect 1104 3834 37812 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 37812 3834
rect 1104 3760 37812 3782
rect 12158 3680 12164 3732
rect 12216 3680 12222 3732
rect 13633 3723 13691 3729
rect 13633 3689 13645 3723
rect 13679 3720 13691 3723
rect 13814 3720 13820 3732
rect 13679 3692 13820 3720
rect 13679 3689 13691 3692
rect 13633 3683 13691 3689
rect 13814 3680 13820 3692
rect 13872 3680 13878 3732
rect 14642 3680 14648 3732
rect 14700 3720 14706 3732
rect 16025 3723 16083 3729
rect 14700 3692 15976 3720
rect 14700 3680 14706 3692
rect 10318 3652 10324 3664
rect 7208 3624 10324 3652
rect 934 3544 940 3596
rect 992 3584 998 3596
rect 1581 3587 1639 3593
rect 1581 3584 1593 3587
rect 992 3556 1593 3584
rect 992 3544 998 3556
rect 1581 3553 1593 3556
rect 1627 3553 1639 3587
rect 1581 3547 1639 3553
rect 2590 3476 2596 3528
rect 2648 3476 2654 3528
rect 7208 3525 7236 3624
rect 10318 3612 10324 3624
rect 10376 3612 10382 3664
rect 10134 3544 10140 3596
rect 10192 3544 10198 3596
rect 12066 3544 12072 3596
rect 12124 3584 12130 3596
rect 15948 3593 15976 3692
rect 16025 3689 16037 3723
rect 16071 3720 16083 3723
rect 16666 3720 16672 3732
rect 16071 3692 16672 3720
rect 16071 3689 16083 3692
rect 16025 3683 16083 3689
rect 16666 3680 16672 3692
rect 16724 3680 16730 3732
rect 17497 3723 17555 3729
rect 17497 3689 17509 3723
rect 17543 3720 17555 3723
rect 18230 3720 18236 3732
rect 17543 3692 18236 3720
rect 17543 3689 17555 3692
rect 17497 3683 17555 3689
rect 18230 3680 18236 3692
rect 18288 3680 18294 3732
rect 26053 3723 26111 3729
rect 26053 3689 26065 3723
rect 26099 3720 26111 3723
rect 26326 3720 26332 3732
rect 26099 3692 26332 3720
rect 26099 3689 26111 3692
rect 26053 3683 26111 3689
rect 26326 3680 26332 3692
rect 26384 3680 26390 3732
rect 26970 3680 26976 3732
rect 27028 3720 27034 3732
rect 28997 3723 29055 3729
rect 27028 3692 28856 3720
rect 27028 3680 27034 3692
rect 28828 3652 28856 3692
rect 28997 3689 29009 3723
rect 29043 3720 29055 3723
rect 29546 3720 29552 3732
rect 29043 3692 29552 3720
rect 29043 3689 29055 3692
rect 28997 3683 29055 3689
rect 29546 3680 29552 3692
rect 29604 3680 29610 3732
rect 30929 3723 30987 3729
rect 30929 3689 30941 3723
rect 30975 3720 30987 3723
rect 32122 3720 32128 3732
rect 30975 3692 32128 3720
rect 30975 3689 30987 3692
rect 30929 3683 30987 3689
rect 32122 3680 32128 3692
rect 32180 3680 32186 3732
rect 32766 3720 32772 3732
rect 32508 3692 32772 3720
rect 29365 3655 29423 3661
rect 29365 3652 29377 3655
rect 28828 3624 29377 3652
rect 29365 3621 29377 3624
rect 29411 3652 29423 3655
rect 29454 3652 29460 3664
rect 29411 3624 29460 3652
rect 29411 3621 29423 3624
rect 29365 3615 29423 3621
rect 29454 3612 29460 3624
rect 29512 3612 29518 3664
rect 12253 3587 12311 3593
rect 12253 3584 12265 3587
rect 12124 3556 12265 3584
rect 12124 3544 12130 3556
rect 12253 3553 12265 3556
rect 12299 3553 12311 3587
rect 12253 3547 12311 3553
rect 15933 3587 15991 3593
rect 15933 3553 15945 3587
rect 15979 3553 15991 3587
rect 15933 3547 15991 3553
rect 7193 3519 7251 3525
rect 7193 3485 7205 3519
rect 7239 3485 7251 3519
rect 7193 3479 7251 3485
rect 8662 3476 8668 3528
rect 8720 3476 8726 3528
rect 10597 3519 10655 3525
rect 10597 3485 10609 3519
rect 10643 3516 10655 3519
rect 10686 3516 10692 3528
rect 10643 3488 10692 3516
rect 10643 3485 10655 3488
rect 10597 3479 10655 3485
rect 10686 3476 10692 3488
rect 10744 3476 10750 3528
rect 10781 3519 10839 3525
rect 10781 3485 10793 3519
rect 10827 3516 10839 3519
rect 12084 3516 12112 3544
rect 10827 3488 12112 3516
rect 10827 3485 10839 3488
rect 10781 3479 10839 3485
rect 15194 3476 15200 3528
rect 15252 3516 15258 3528
rect 15666 3519 15724 3525
rect 15666 3516 15678 3519
rect 15252 3488 15678 3516
rect 15252 3476 15258 3488
rect 15666 3485 15678 3488
rect 15712 3485 15724 3519
rect 15948 3516 15976 3547
rect 19242 3544 19248 3596
rect 19300 3544 19306 3596
rect 26421 3587 26479 3593
rect 26421 3584 26433 3587
rect 26206 3556 26433 3584
rect 17402 3516 17408 3528
rect 15948 3488 17408 3516
rect 15666 3479 15724 3485
rect 17402 3476 17408 3488
rect 17460 3516 17466 3528
rect 18877 3519 18935 3525
rect 18877 3516 18889 3519
rect 17460 3488 18889 3516
rect 17460 3476 17466 3488
rect 18877 3485 18889 3488
rect 18923 3485 18935 3519
rect 18877 3479 18935 3485
rect 24673 3519 24731 3525
rect 24673 3485 24685 3519
rect 24719 3485 24731 3519
rect 24673 3479 24731 3485
rect 24940 3519 24998 3525
rect 24940 3485 24952 3519
rect 24986 3485 24998 3519
rect 24940 3479 24998 3485
rect 6638 3408 6644 3460
rect 6696 3408 6702 3460
rect 8294 3408 8300 3460
rect 8352 3408 8358 3460
rect 11054 3457 11060 3460
rect 11048 3448 11060 3457
rect 11015 3420 11060 3448
rect 11048 3411 11060 3420
rect 11054 3408 11060 3411
rect 11112 3408 11118 3460
rect 12066 3408 12072 3460
rect 12124 3448 12130 3460
rect 12498 3451 12556 3457
rect 12498 3448 12510 3451
rect 12124 3420 12510 3448
rect 12124 3408 12130 3420
rect 12498 3417 12510 3420
rect 12544 3417 12556 3451
rect 12498 3411 12556 3417
rect 17160 3451 17218 3457
rect 17160 3417 17172 3451
rect 17206 3448 17218 3451
rect 17954 3448 17960 3460
rect 17206 3420 17960 3448
rect 17206 3417 17218 3420
rect 17160 3411 17218 3417
rect 17954 3408 17960 3420
rect 18012 3408 18018 3460
rect 18632 3451 18690 3457
rect 18632 3417 18644 3451
rect 18678 3448 18690 3451
rect 18782 3448 18788 3460
rect 18678 3420 18788 3448
rect 18678 3417 18690 3420
rect 18632 3411 18690 3417
rect 18782 3408 18788 3420
rect 18840 3408 18846 3460
rect 14550 3340 14556 3392
rect 14608 3340 14614 3392
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 19889 3383 19947 3389
rect 19889 3380 19901 3383
rect 19484 3352 19901 3380
rect 19484 3340 19490 3352
rect 19889 3349 19901 3352
rect 19935 3349 19947 3383
rect 24688 3380 24716 3479
rect 24854 3408 24860 3460
rect 24912 3448 24918 3460
rect 24964 3448 24992 3479
rect 24912 3420 24992 3448
rect 24912 3408 24918 3420
rect 26206 3380 26234 3556
rect 26421 3553 26433 3556
rect 26467 3584 26479 3587
rect 27522 3584 27528 3596
rect 26467 3556 27528 3584
rect 26467 3553 26479 3556
rect 26421 3547 26479 3553
rect 27522 3544 27528 3556
rect 27580 3584 27586 3596
rect 32508 3593 32536 3692
rect 32766 3680 32772 3692
rect 32824 3680 32830 3732
rect 33873 3723 33931 3729
rect 33873 3689 33885 3723
rect 33919 3720 33931 3723
rect 34330 3720 34336 3732
rect 33919 3692 34336 3720
rect 33919 3689 33931 3692
rect 33873 3683 33931 3689
rect 34330 3680 34336 3692
rect 34388 3680 34394 3732
rect 34514 3720 34520 3732
rect 34440 3692 34520 3720
rect 33965 3655 34023 3661
rect 33965 3621 33977 3655
rect 34011 3621 34023 3655
rect 33965 3615 34023 3621
rect 34149 3655 34207 3661
rect 34149 3621 34161 3655
rect 34195 3652 34207 3655
rect 34440 3652 34468 3692
rect 34514 3680 34520 3692
rect 34572 3680 34578 3732
rect 34606 3680 34612 3732
rect 34664 3720 34670 3732
rect 34664 3692 36768 3720
rect 34664 3680 34670 3692
rect 34195 3624 34468 3652
rect 34532 3624 34744 3652
rect 34195 3621 34207 3624
rect 34149 3615 34207 3621
rect 32493 3587 32551 3593
rect 27580 3556 27660 3584
rect 27580 3544 27586 3556
rect 26878 3476 26884 3528
rect 26936 3476 26942 3528
rect 27062 3476 27068 3528
rect 27120 3516 27126 3528
rect 27632 3525 27660 3556
rect 32493 3553 32505 3587
rect 32539 3553 32551 3587
rect 32493 3547 32551 3553
rect 27433 3519 27491 3525
rect 27433 3516 27445 3519
rect 27120 3488 27445 3516
rect 27120 3476 27126 3488
rect 27433 3485 27445 3488
rect 27479 3485 27491 3519
rect 27433 3479 27491 3485
rect 27617 3519 27675 3525
rect 27617 3485 27629 3519
rect 27663 3516 27675 3519
rect 29086 3516 29092 3528
rect 27663 3488 29092 3516
rect 27663 3485 27675 3488
rect 27617 3479 27675 3485
rect 29086 3476 29092 3488
rect 29144 3516 29150 3528
rect 29546 3516 29552 3528
rect 29144 3488 29552 3516
rect 29144 3476 29150 3488
rect 29546 3476 29552 3488
rect 29604 3516 29610 3528
rect 31021 3519 31079 3525
rect 31021 3516 31033 3519
rect 29604 3488 31033 3516
rect 29604 3476 29610 3488
rect 31021 3485 31033 3488
rect 31067 3485 31079 3519
rect 31021 3479 31079 3485
rect 32760 3519 32818 3525
rect 32760 3485 32772 3519
rect 32806 3516 32818 3519
rect 33980 3516 34008 3615
rect 34422 3544 34428 3596
rect 34480 3544 34486 3596
rect 32806 3488 34008 3516
rect 32806 3485 32818 3488
rect 32760 3479 32818 3485
rect 26786 3408 26792 3460
rect 26844 3448 26850 3460
rect 27862 3451 27920 3457
rect 27862 3448 27874 3451
rect 26844 3420 27874 3448
rect 26844 3408 26850 3420
rect 27862 3417 27874 3420
rect 27908 3417 27920 3451
rect 27862 3411 27920 3417
rect 29816 3451 29874 3457
rect 29816 3417 29828 3451
rect 29862 3448 29874 3451
rect 30098 3448 30104 3460
rect 29862 3420 30104 3448
rect 29862 3417 29874 3420
rect 29816 3411 29874 3417
rect 30098 3408 30104 3420
rect 30156 3408 30162 3460
rect 31036 3392 31064 3479
rect 34146 3476 34152 3528
rect 34204 3516 34210 3528
rect 34532 3516 34560 3624
rect 34716 3593 34744 3624
rect 35710 3612 35716 3664
rect 35768 3652 35774 3664
rect 36173 3655 36231 3661
rect 36173 3652 36185 3655
rect 35768 3624 36185 3652
rect 35768 3612 35774 3624
rect 36173 3621 36185 3624
rect 36219 3621 36231 3655
rect 36173 3615 36231 3621
rect 36740 3593 36768 3692
rect 37090 3680 37096 3732
rect 37148 3680 37154 3732
rect 34701 3587 34759 3593
rect 34701 3553 34713 3587
rect 34747 3553 34759 3587
rect 34701 3547 34759 3553
rect 36725 3587 36783 3593
rect 36725 3553 36737 3587
rect 36771 3553 36783 3587
rect 36725 3547 36783 3553
rect 34204 3488 34560 3516
rect 34204 3476 34210 3488
rect 36170 3476 36176 3528
rect 36228 3476 36234 3528
rect 31288 3451 31346 3457
rect 31288 3417 31300 3451
rect 31334 3448 31346 3451
rect 31386 3448 31392 3460
rect 31334 3420 31392 3448
rect 31334 3417 31346 3420
rect 31288 3411 31346 3417
rect 31386 3408 31392 3420
rect 31444 3408 31450 3460
rect 32674 3408 32680 3460
rect 32732 3448 32738 3460
rect 34946 3451 35004 3457
rect 34946 3448 34958 3451
rect 32732 3420 34958 3448
rect 32732 3408 32738 3420
rect 34946 3417 34958 3420
rect 34992 3417 35004 3451
rect 34946 3411 35004 3417
rect 24688 3352 26234 3380
rect 19889 3343 19947 3349
rect 31018 3340 31024 3392
rect 31076 3340 31082 3392
rect 32401 3383 32459 3389
rect 32401 3349 32413 3383
rect 32447 3380 32459 3383
rect 33686 3380 33692 3392
rect 32447 3352 33692 3380
rect 32447 3349 32459 3352
rect 32401 3343 32459 3349
rect 33686 3340 33692 3352
rect 33744 3340 33750 3392
rect 34514 3340 34520 3392
rect 34572 3380 34578 3392
rect 34790 3380 34796 3392
rect 34572 3352 34796 3380
rect 34572 3340 34578 3352
rect 34790 3340 34796 3352
rect 34848 3340 34854 3392
rect 36081 3383 36139 3389
rect 36081 3349 36093 3383
rect 36127 3380 36139 3383
rect 36188 3380 36216 3476
rect 36262 3408 36268 3460
rect 36320 3448 36326 3460
rect 36906 3448 36912 3460
rect 36320 3420 36912 3448
rect 36320 3408 36326 3420
rect 36906 3408 36912 3420
rect 36964 3448 36970 3460
rect 37001 3451 37059 3457
rect 37001 3448 37013 3451
rect 36964 3420 37013 3448
rect 36964 3408 36970 3420
rect 37001 3417 37013 3420
rect 37047 3417 37059 3451
rect 37001 3411 37059 3417
rect 36127 3352 36216 3380
rect 36127 3349 36139 3352
rect 36081 3343 36139 3349
rect 1104 3290 37812 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 37812 3290
rect 1104 3216 37812 3238
rect 8294 3136 8300 3188
rect 8352 3136 8358 3188
rect 12066 3136 12072 3188
rect 12124 3136 12130 3188
rect 15838 3176 15844 3188
rect 14936 3148 15844 3176
rect 2590 3000 2596 3052
rect 2648 3000 2654 3052
rect 8312 3049 8340 3136
rect 9784 3080 12296 3108
rect 9784 3049 9812 3080
rect 12268 3052 12296 3080
rect 8297 3043 8355 3049
rect 8297 3009 8309 3043
rect 8343 3009 8355 3043
rect 8297 3003 8355 3009
rect 9769 3043 9827 3049
rect 9769 3009 9781 3043
rect 9815 3009 9827 3043
rect 9769 3003 9827 3009
rect 9950 3000 9956 3052
rect 10008 3000 10014 3052
rect 11241 3043 11299 3049
rect 11241 3009 11253 3043
rect 11287 3040 11299 3043
rect 11974 3040 11980 3052
rect 11287 3012 11980 3040
rect 11287 3009 11299 3012
rect 11241 3003 11299 3009
rect 11974 3000 11980 3012
rect 12032 3000 12038 3052
rect 12250 3000 12256 3052
rect 12308 3000 12314 3052
rect 13449 3043 13507 3049
rect 13449 3009 13461 3043
rect 13495 3040 13507 3043
rect 14090 3040 14096 3052
rect 13495 3012 14096 3040
rect 13495 3009 13507 3012
rect 13449 3003 13507 3009
rect 14090 3000 14096 3012
rect 14148 3000 14154 3052
rect 14936 3049 14964 3148
rect 15838 3136 15844 3148
rect 15896 3136 15902 3188
rect 17402 3136 17408 3188
rect 17460 3136 17466 3188
rect 17954 3136 17960 3188
rect 18012 3136 18018 3188
rect 18785 3179 18843 3185
rect 18785 3145 18797 3179
rect 18831 3176 18843 3179
rect 19150 3176 19156 3188
rect 18831 3148 19156 3176
rect 18831 3145 18843 3148
rect 18785 3139 18843 3145
rect 19150 3136 19156 3148
rect 19208 3136 19214 3188
rect 19426 3136 19432 3188
rect 19484 3136 19490 3188
rect 25317 3179 25375 3185
rect 25317 3145 25329 3179
rect 25363 3176 25375 3179
rect 26234 3176 26240 3188
rect 25363 3148 26240 3176
rect 25363 3145 25375 3148
rect 25317 3139 25375 3145
rect 26206 3136 26240 3148
rect 26292 3136 26298 3188
rect 26786 3136 26792 3188
rect 26844 3136 26850 3188
rect 26973 3179 27031 3185
rect 26973 3145 26985 3179
rect 27019 3176 27031 3179
rect 27154 3176 27160 3188
rect 27019 3148 27160 3176
rect 27019 3145 27031 3148
rect 26973 3139 27031 3145
rect 27154 3136 27160 3148
rect 27212 3136 27218 3188
rect 29546 3136 29552 3188
rect 29604 3136 29610 3188
rect 30466 3136 30472 3188
rect 30524 3136 30530 3188
rect 31018 3136 31024 3188
rect 31076 3176 31082 3188
rect 33137 3179 33195 3185
rect 33137 3176 33149 3179
rect 31076 3148 33149 3176
rect 31076 3136 31082 3148
rect 33137 3145 33149 3148
rect 33183 3145 33195 3179
rect 33137 3139 33195 3145
rect 34238 3136 34244 3188
rect 34296 3176 34302 3188
rect 35069 3179 35127 3185
rect 35069 3176 35081 3179
rect 34296 3148 35081 3176
rect 34296 3136 34302 3148
rect 35069 3145 35081 3148
rect 35115 3145 35127 3179
rect 35069 3139 35127 3145
rect 15286 3068 15292 3120
rect 15344 3068 15350 3120
rect 14921 3043 14979 3049
rect 14921 3009 14933 3043
rect 14967 3009 14979 3043
rect 14921 3003 14979 3009
rect 15654 3000 15660 3052
rect 15712 3040 15718 3052
rect 15749 3043 15807 3049
rect 15749 3040 15761 3043
rect 15712 3012 15761 3040
rect 15712 3000 15718 3012
rect 15749 3009 15761 3012
rect 15795 3009 15807 3043
rect 15749 3003 15807 3009
rect 17310 3000 17316 3052
rect 17368 3000 17374 3052
rect 17420 3049 17448 3136
rect 17678 3117 17684 3120
rect 17672 3071 17684 3117
rect 17736 3108 17742 3120
rect 17736 3080 17772 3108
rect 17678 3068 17684 3071
rect 17736 3068 17742 3080
rect 17405 3043 17463 3049
rect 17405 3009 17417 3043
rect 17451 3009 17463 3043
rect 17972 3040 18000 3136
rect 19444 3040 19472 3136
rect 20622 3108 20628 3120
rect 19720 3080 20628 3108
rect 19613 3043 19671 3049
rect 19613 3040 19625 3043
rect 17972 3012 18920 3040
rect 19444 3012 19625 3040
rect 17405 3003 17463 3009
rect 1578 2932 1584 2984
rect 1636 2932 1642 2984
rect 7650 2932 7656 2984
rect 7708 2932 7714 2984
rect 8754 2932 8760 2984
rect 8812 2972 8818 2984
rect 9217 2975 9275 2981
rect 9217 2972 9229 2975
rect 8812 2944 9229 2972
rect 8812 2932 8818 2944
rect 9217 2941 9229 2944
rect 9263 2941 9275 2975
rect 9217 2935 9275 2941
rect 9968 2904 9996 3000
rect 10965 2975 11023 2981
rect 10965 2941 10977 2975
rect 11011 2972 11023 2975
rect 11146 2972 11152 2984
rect 11011 2944 11152 2972
rect 11011 2941 11023 2944
rect 10965 2935 11023 2941
rect 11146 2932 11152 2944
rect 11204 2932 11210 2984
rect 11609 2975 11667 2981
rect 11609 2941 11621 2975
rect 11655 2972 11667 2975
rect 12345 2975 12403 2981
rect 12345 2972 12357 2975
rect 11655 2944 12357 2972
rect 11655 2941 11667 2944
rect 11609 2935 11667 2941
rect 12345 2941 12357 2944
rect 12391 2941 12403 2975
rect 12345 2935 12403 2941
rect 11624 2904 11652 2935
rect 12894 2932 12900 2984
rect 12952 2932 12958 2984
rect 14645 2975 14703 2981
rect 14645 2941 14657 2975
rect 14691 2972 14703 2975
rect 15194 2972 15200 2984
rect 14691 2944 15200 2972
rect 14691 2941 14703 2944
rect 14645 2935 14703 2941
rect 15194 2932 15200 2944
rect 15252 2932 15258 2984
rect 18892 2981 18920 3012
rect 19613 3009 19625 3012
rect 19659 3009 19671 3043
rect 19613 3003 19671 3009
rect 18877 2975 18935 2981
rect 18877 2941 18889 2975
rect 18923 2941 18935 2975
rect 18877 2935 18935 2941
rect 19334 2932 19340 2984
rect 19392 2972 19398 2984
rect 19720 2972 19748 3080
rect 20622 3068 20628 3080
rect 20680 3068 20686 3120
rect 26206 3108 26234 3136
rect 26329 3111 26387 3117
rect 26329 3108 26341 3111
rect 26206 3080 26341 3108
rect 26329 3077 26341 3080
rect 26375 3077 26387 3111
rect 26329 3071 26387 3077
rect 27706 3068 27712 3120
rect 27764 3108 27770 3120
rect 28086 3111 28144 3117
rect 28086 3108 28098 3111
rect 27764 3080 28098 3108
rect 27764 3068 27770 3080
rect 28086 3077 28098 3080
rect 28132 3077 28144 3111
rect 29564 3108 29592 3136
rect 28086 3071 28144 3077
rect 28368 3080 29592 3108
rect 30377 3111 30435 3117
rect 22005 3043 22063 3049
rect 22005 3009 22017 3043
rect 22051 3040 22063 3043
rect 22186 3040 22192 3052
rect 22051 3012 22192 3040
rect 22051 3009 22063 3012
rect 22005 3003 22063 3009
rect 22186 3000 22192 3012
rect 22244 3000 22250 3052
rect 23382 3000 23388 3052
rect 23440 3000 23446 3052
rect 26053 3043 26111 3049
rect 26053 3009 26065 3043
rect 26099 3040 26111 3043
rect 27338 3040 27344 3052
rect 26099 3012 27344 3040
rect 26099 3009 26111 3012
rect 26053 3003 26111 3009
rect 27338 3000 27344 3012
rect 27396 3000 27402 3052
rect 28368 3049 28396 3080
rect 30377 3077 30389 3111
rect 30423 3108 30435 3111
rect 30484 3108 30512 3136
rect 30423 3080 30512 3108
rect 30423 3077 30435 3080
rect 30377 3071 30435 3077
rect 31386 3068 31392 3120
rect 31444 3068 31450 3120
rect 31846 3068 31852 3120
rect 31904 3068 31910 3120
rect 33502 3068 33508 3120
rect 33560 3108 33566 3120
rect 36173 3111 36231 3117
rect 36173 3108 36185 3111
rect 33560 3080 36185 3108
rect 33560 3068 33566 3080
rect 36173 3077 36185 3080
rect 36219 3077 36231 3111
rect 36173 3071 36231 3077
rect 28353 3043 28411 3049
rect 28353 3009 28365 3043
rect 28399 3009 28411 3043
rect 28353 3003 28411 3009
rect 28442 3000 28448 3052
rect 28500 3040 28506 3052
rect 28537 3043 28595 3049
rect 28537 3040 28549 3043
rect 28500 3012 28549 3040
rect 28500 3000 28506 3012
rect 28537 3009 28549 3012
rect 28583 3009 28595 3043
rect 28537 3003 28595 3009
rect 29362 3000 29368 3052
rect 29420 3040 29426 3052
rect 30009 3043 30067 3049
rect 30009 3040 30021 3043
rect 29420 3012 30021 3040
rect 29420 3000 29426 3012
rect 30009 3009 30021 3012
rect 30055 3009 30067 3043
rect 30009 3003 30067 3009
rect 19392 2944 19748 2972
rect 19392 2932 19398 2944
rect 20070 2932 20076 2984
rect 20128 2932 20134 2984
rect 20898 2932 20904 2984
rect 20956 2972 20962 2984
rect 22281 2975 22339 2981
rect 22281 2972 22293 2975
rect 20956 2944 22293 2972
rect 20956 2932 20962 2944
rect 22281 2941 22293 2944
rect 22327 2941 22339 2975
rect 22281 2935 22339 2941
rect 23934 2932 23940 2984
rect 23992 2932 23998 2984
rect 25777 2975 25835 2981
rect 25777 2941 25789 2975
rect 25823 2972 25835 2975
rect 26970 2972 26976 2984
rect 25823 2944 26234 2972
rect 25823 2941 25835 2944
rect 25777 2935 25835 2941
rect 9968 2876 11652 2904
rect 11977 2907 12035 2913
rect 11977 2873 11989 2907
rect 12023 2904 12035 2907
rect 13722 2904 13728 2916
rect 12023 2876 13728 2904
rect 12023 2873 12035 2876
rect 11977 2867 12035 2873
rect 13722 2864 13728 2876
rect 13780 2864 13786 2916
rect 18969 2907 19027 2913
rect 18969 2873 18981 2907
rect 19015 2873 19027 2907
rect 26206 2904 26234 2944
rect 26436 2944 26976 2972
rect 26436 2904 26464 2944
rect 26970 2932 26976 2944
rect 27028 2932 27034 2984
rect 29086 2932 29092 2984
rect 29144 2932 29150 2984
rect 31404 2981 31432 3068
rect 31938 3000 31944 3052
rect 31996 3040 32002 3052
rect 32217 3043 32275 3049
rect 32217 3040 32229 3043
rect 31996 3012 32229 3040
rect 31996 3000 32002 3012
rect 32217 3009 32229 3012
rect 32263 3009 32275 3043
rect 32217 3003 32275 3009
rect 32769 3043 32827 3049
rect 32769 3009 32781 3043
rect 32815 3040 32827 3043
rect 33597 3043 33655 3049
rect 33597 3040 33609 3043
rect 32815 3012 33609 3040
rect 32815 3009 32827 3012
rect 32769 3003 32827 3009
rect 33597 3009 33609 3012
rect 33643 3009 33655 3043
rect 33597 3003 33655 3009
rect 33870 3000 33876 3052
rect 33928 3040 33934 3052
rect 35342 3040 35348 3052
rect 33928 3012 35348 3040
rect 33928 3000 33934 3012
rect 35342 3000 35348 3012
rect 35400 3000 35406 3052
rect 35618 3000 35624 3052
rect 35676 3040 35682 3052
rect 35805 3043 35863 3049
rect 35805 3040 35817 3043
rect 35676 3012 35817 3040
rect 35676 3000 35682 3012
rect 35805 3009 35817 3012
rect 35851 3009 35863 3043
rect 35805 3003 35863 3009
rect 31389 2975 31447 2981
rect 31389 2941 31401 2975
rect 31435 2941 31447 2975
rect 34057 2975 34115 2981
rect 34057 2972 34069 2975
rect 31389 2935 31447 2941
rect 33888 2944 34069 2972
rect 26206 2876 26464 2904
rect 26697 2907 26755 2913
rect 18969 2867 19027 2873
rect 26697 2873 26709 2907
rect 26743 2873 26755 2907
rect 26697 2867 26755 2873
rect 31573 2907 31631 2913
rect 31573 2873 31585 2907
rect 31619 2904 31631 2907
rect 33042 2904 33048 2916
rect 31619 2876 33048 2904
rect 31619 2873 31631 2876
rect 31573 2867 31631 2873
rect 1762 2796 1768 2848
rect 1820 2836 1826 2848
rect 2869 2839 2927 2845
rect 2869 2836 2881 2839
rect 1820 2808 2881 2836
rect 1820 2796 1826 2808
rect 2869 2805 2881 2808
rect 2915 2805 2927 2839
rect 2869 2799 2927 2805
rect 16669 2839 16727 2845
rect 16669 2805 16681 2839
rect 16715 2836 16727 2839
rect 16942 2836 16948 2848
rect 16715 2808 16948 2836
rect 16715 2805 16727 2808
rect 16669 2799 16727 2805
rect 16942 2796 16948 2808
rect 17000 2836 17006 2848
rect 18984 2836 19012 2867
rect 17000 2808 19012 2836
rect 26712 2836 26740 2867
rect 33042 2864 33048 2876
rect 33100 2864 33106 2916
rect 28166 2836 28172 2848
rect 26712 2808 28172 2836
rect 17000 2796 17006 2808
rect 28166 2796 28172 2808
rect 28224 2796 28230 2848
rect 31202 2796 31208 2848
rect 31260 2836 31266 2848
rect 33888 2836 33916 2944
rect 34057 2941 34069 2944
rect 34103 2941 34115 2975
rect 34057 2935 34115 2941
rect 34422 2932 34428 2984
rect 34480 2972 34486 2984
rect 35529 2975 35587 2981
rect 35529 2972 35541 2975
rect 34480 2944 35541 2972
rect 34480 2932 34486 2944
rect 35529 2941 35541 2944
rect 35575 2972 35587 2975
rect 36725 2975 36783 2981
rect 36725 2972 36737 2975
rect 35575 2944 36737 2972
rect 35575 2941 35587 2944
rect 35529 2935 35587 2941
rect 36725 2941 36737 2944
rect 36771 2941 36783 2975
rect 36725 2935 36783 2941
rect 34238 2864 34244 2916
rect 34296 2904 34302 2916
rect 35161 2907 35219 2913
rect 35161 2904 35173 2907
rect 34296 2876 35173 2904
rect 34296 2864 34302 2876
rect 35161 2873 35173 2876
rect 35207 2873 35219 2907
rect 35161 2867 35219 2873
rect 31260 2808 33916 2836
rect 31260 2796 31266 2808
rect 1104 2746 37812 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 37812 2746
rect 1104 2672 37812 2694
rect 12434 2592 12440 2644
rect 12492 2592 12498 2644
rect 15013 2635 15071 2641
rect 15013 2601 15025 2635
rect 15059 2632 15071 2635
rect 15470 2632 15476 2644
rect 15059 2604 15476 2632
rect 15059 2601 15071 2604
rect 15013 2595 15071 2601
rect 15470 2592 15476 2604
rect 15528 2592 15534 2644
rect 16482 2592 16488 2644
rect 16540 2632 16546 2644
rect 16669 2635 16727 2641
rect 16669 2632 16681 2635
rect 16540 2604 16681 2632
rect 16540 2592 16546 2604
rect 16669 2601 16681 2604
rect 16715 2601 16727 2635
rect 16669 2595 16727 2601
rect 19242 2592 19248 2644
rect 19300 2592 19306 2644
rect 19978 2632 19984 2644
rect 19904 2604 19984 2632
rect 9401 2567 9459 2573
rect 9401 2533 9413 2567
rect 9447 2564 9459 2567
rect 16850 2564 16856 2576
rect 9447 2536 16856 2564
rect 9447 2533 9459 2536
rect 9401 2527 9459 2533
rect 16850 2524 16856 2536
rect 16908 2524 16914 2576
rect 2409 2499 2467 2505
rect 2409 2465 2421 2499
rect 2455 2496 2467 2499
rect 2590 2496 2596 2508
rect 2455 2468 2596 2496
rect 2455 2465 2467 2468
rect 2409 2459 2467 2465
rect 2590 2456 2596 2468
rect 2648 2456 2654 2508
rect 5721 2499 5779 2505
rect 5721 2465 5733 2499
rect 5767 2496 5779 2499
rect 6086 2496 6092 2508
rect 5767 2468 6092 2496
rect 5767 2465 5779 2468
rect 5721 2459 5779 2465
rect 6086 2456 6092 2468
rect 6144 2456 6150 2508
rect 8297 2499 8355 2505
rect 8297 2465 8309 2499
rect 8343 2496 8355 2499
rect 9122 2496 9128 2508
rect 8343 2468 9128 2496
rect 8343 2465 8355 2468
rect 8297 2459 8355 2465
rect 9122 2456 9128 2468
rect 9180 2456 9186 2508
rect 10873 2499 10931 2505
rect 10873 2465 10885 2499
rect 10919 2496 10931 2499
rect 12066 2496 12072 2508
rect 10919 2468 12072 2496
rect 10919 2465 10931 2468
rect 10873 2459 10931 2465
rect 12066 2456 12072 2468
rect 12124 2456 12130 2508
rect 12526 2456 12532 2508
rect 12584 2456 12590 2508
rect 12618 2456 12624 2508
rect 12676 2456 12682 2508
rect 14461 2499 14519 2505
rect 14461 2465 14473 2499
rect 14507 2496 14519 2499
rect 14550 2496 14556 2508
rect 14507 2468 14556 2496
rect 14507 2465 14519 2468
rect 14461 2459 14519 2465
rect 14550 2456 14556 2468
rect 14608 2456 14614 2508
rect 17218 2456 17224 2508
rect 17276 2456 17282 2508
rect 18138 2456 18144 2508
rect 18196 2456 18202 2508
rect 19904 2505 19932 2604
rect 19978 2592 19984 2604
rect 20036 2592 20042 2644
rect 26142 2592 26148 2644
rect 26200 2592 26206 2644
rect 28445 2635 28503 2641
rect 28445 2601 28457 2635
rect 28491 2632 28503 2635
rect 28534 2632 28540 2644
rect 28491 2604 28540 2632
rect 28491 2601 28503 2604
rect 28445 2595 28503 2601
rect 28534 2592 28540 2604
rect 28592 2592 28598 2644
rect 28718 2592 28724 2644
rect 28776 2632 28782 2644
rect 31021 2635 31079 2641
rect 31021 2632 31033 2635
rect 28776 2604 31033 2632
rect 28776 2592 28782 2604
rect 31021 2601 31033 2604
rect 31067 2601 31079 2635
rect 31021 2595 31079 2601
rect 31846 2592 31852 2644
rect 31904 2632 31910 2644
rect 33137 2635 33195 2641
rect 33137 2632 33149 2635
rect 31904 2604 33149 2632
rect 31904 2592 31910 2604
rect 33137 2601 33149 2604
rect 33183 2601 33195 2635
rect 33137 2595 33195 2601
rect 33152 2564 33180 2595
rect 33594 2592 33600 2644
rect 33652 2592 33658 2644
rect 35894 2592 35900 2644
rect 35952 2632 35958 2644
rect 36173 2635 36231 2641
rect 36173 2632 36185 2635
rect 35952 2604 36185 2632
rect 35952 2592 35958 2604
rect 36173 2601 36185 2604
rect 36219 2601 36231 2635
rect 36173 2595 36231 2601
rect 37274 2592 37280 2644
rect 37332 2592 37338 2644
rect 34422 2564 34428 2576
rect 33152 2536 34428 2564
rect 34422 2524 34428 2536
rect 34480 2524 34486 2576
rect 34514 2524 34520 2576
rect 34572 2564 34578 2576
rect 34572 2536 36768 2564
rect 34572 2524 34578 2536
rect 19889 2499 19947 2505
rect 19889 2465 19901 2499
rect 19935 2465 19947 2499
rect 19889 2459 19947 2465
rect 19978 2456 19984 2508
rect 20036 2496 20042 2508
rect 20441 2499 20499 2505
rect 20441 2496 20453 2499
rect 20036 2468 20453 2496
rect 20036 2456 20042 2468
rect 20441 2465 20453 2468
rect 20487 2465 20499 2499
rect 20441 2459 20499 2465
rect 22186 2456 22192 2508
rect 22244 2456 22250 2508
rect 22830 2456 22836 2508
rect 22888 2496 22894 2508
rect 24857 2499 24915 2505
rect 24857 2496 24869 2499
rect 22888 2468 24869 2496
rect 22888 2456 22894 2468
rect 24857 2465 24869 2468
rect 24903 2465 24915 2499
rect 27433 2499 27491 2505
rect 27433 2496 27445 2499
rect 24857 2459 24915 2465
rect 26206 2468 27445 2496
rect 2682 2388 2688 2440
rect 2740 2388 2746 2440
rect 3326 2388 3332 2440
rect 3384 2388 3390 2440
rect 4706 2388 4712 2440
rect 4764 2388 4770 2440
rect 6181 2431 6239 2437
rect 6181 2397 6193 2431
rect 6227 2428 6239 2431
rect 6638 2428 6644 2440
rect 6227 2400 6644 2428
rect 6227 2397 6239 2400
rect 6181 2391 6239 2397
rect 6638 2388 6644 2400
rect 6696 2388 6702 2440
rect 8754 2388 8760 2440
rect 8812 2388 8818 2440
rect 9217 2431 9275 2437
rect 9217 2397 9229 2431
rect 9263 2397 9275 2431
rect 9217 2391 9275 2397
rect 9232 2360 9260 2391
rect 11146 2388 11152 2440
rect 11204 2388 11210 2440
rect 11885 2431 11943 2437
rect 11885 2397 11897 2431
rect 11931 2428 11943 2431
rect 12544 2428 12572 2456
rect 11931 2400 12572 2428
rect 11931 2397 11943 2400
rect 11885 2391 11943 2397
rect 12636 2360 12664 2456
rect 12713 2431 12771 2437
rect 12713 2397 12725 2431
rect 12759 2428 12771 2431
rect 12894 2428 12900 2440
rect 12759 2400 12900 2428
rect 12759 2397 12771 2400
rect 12713 2391 12771 2397
rect 12894 2388 12900 2400
rect 12952 2388 12958 2440
rect 15194 2388 15200 2440
rect 15252 2388 15258 2440
rect 17865 2431 17923 2437
rect 17865 2397 17877 2431
rect 17911 2428 17923 2431
rect 18046 2428 18052 2440
rect 17911 2400 18052 2428
rect 17911 2397 17923 2400
rect 17865 2391 17923 2397
rect 18046 2388 18052 2400
rect 18104 2388 18110 2440
rect 20070 2388 20076 2440
rect 20128 2388 20134 2440
rect 20714 2388 20720 2440
rect 20772 2428 20778 2440
rect 21913 2431 21971 2437
rect 21913 2428 21925 2431
rect 20772 2400 21925 2428
rect 20772 2388 20778 2400
rect 21913 2397 21925 2400
rect 21959 2397 21971 2431
rect 21913 2391 21971 2397
rect 23934 2388 23940 2440
rect 23992 2428 23998 2440
rect 24397 2431 24455 2437
rect 24397 2428 24409 2431
rect 23992 2400 24409 2428
rect 23992 2388 23998 2400
rect 24397 2397 24409 2400
rect 24443 2397 24455 2431
rect 24397 2391 24455 2397
rect 9232 2332 12664 2360
rect 13538 2320 13544 2372
rect 13596 2320 13602 2372
rect 16298 2320 16304 2372
rect 16356 2320 16362 2372
rect 24118 2320 24124 2372
rect 24176 2360 24182 2372
rect 26206 2360 26234 2468
rect 27433 2465 27445 2468
rect 27479 2465 27491 2499
rect 30009 2499 30067 2505
rect 30009 2496 30021 2499
rect 27433 2459 27491 2465
rect 27632 2468 30021 2496
rect 26694 2388 26700 2440
rect 26752 2388 26758 2440
rect 26970 2388 26976 2440
rect 27028 2388 27034 2440
rect 27154 2388 27160 2440
rect 27212 2428 27218 2440
rect 27632 2428 27660 2468
rect 30009 2465 30021 2468
rect 30055 2465 30067 2499
rect 30009 2459 30067 2465
rect 30282 2456 30288 2508
rect 30340 2496 30346 2508
rect 31573 2499 31631 2505
rect 31573 2496 31585 2499
rect 30340 2468 31585 2496
rect 30340 2456 30346 2468
rect 31573 2465 31585 2468
rect 31619 2465 31631 2499
rect 31573 2459 31631 2465
rect 32490 2456 32496 2508
rect 32548 2456 32554 2508
rect 33134 2456 33140 2508
rect 33192 2496 33198 2508
rect 36740 2505 36768 2536
rect 35161 2499 35219 2505
rect 35161 2496 35173 2499
rect 33192 2468 35173 2496
rect 33192 2456 33198 2468
rect 35161 2465 35173 2468
rect 35207 2465 35219 2499
rect 35161 2459 35219 2465
rect 36725 2499 36783 2505
rect 36725 2465 36737 2499
rect 36771 2465 36783 2499
rect 36725 2459 36783 2465
rect 27212 2400 27660 2428
rect 27212 2388 27218 2400
rect 27798 2388 27804 2440
rect 27856 2428 27862 2440
rect 28997 2431 29055 2437
rect 28997 2428 29009 2431
rect 27856 2400 29009 2428
rect 27856 2388 27862 2400
rect 28997 2397 29009 2400
rect 29043 2397 29055 2431
rect 28997 2391 29055 2397
rect 29086 2388 29092 2440
rect 29144 2428 29150 2440
rect 29549 2431 29607 2437
rect 29549 2428 29561 2431
rect 29144 2400 29561 2428
rect 29144 2388 29150 2400
rect 29549 2397 29561 2400
rect 29595 2397 29607 2431
rect 29549 2391 29607 2397
rect 31754 2388 31760 2440
rect 31812 2428 31818 2440
rect 32217 2431 32275 2437
rect 32217 2428 32229 2431
rect 31812 2400 32229 2428
rect 31812 2388 31818 2400
rect 32217 2397 32229 2400
rect 32263 2397 32275 2431
rect 32217 2391 32275 2397
rect 33226 2388 33232 2440
rect 33284 2428 33290 2440
rect 34149 2431 34207 2437
rect 34149 2428 34161 2431
rect 33284 2400 34161 2428
rect 33284 2388 33290 2400
rect 34149 2397 34161 2400
rect 34195 2397 34207 2431
rect 34149 2391 34207 2397
rect 34698 2388 34704 2440
rect 34756 2388 34762 2440
rect 37461 2431 37519 2437
rect 37461 2397 37473 2431
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 24176 2332 26234 2360
rect 37476 2360 37504 2391
rect 37918 2360 37924 2372
rect 37476 2332 37924 2360
rect 24176 2320 24182 2332
rect 37918 2320 37924 2332
rect 37976 2320 37982 2372
rect 1104 2202 37812 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 37812 2202
rect 1104 2128 37812 2150
rect 21634 1300 21640 1352
rect 21692 1340 21698 1352
rect 34514 1340 34520 1352
rect 21692 1312 34520 1340
rect 21692 1300 21698 1312
rect 34514 1300 34520 1312
rect 34572 1300 34578 1352
<< via1 >>
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 29368 36252 29420 36304
rect 2872 36227 2924 36236
rect 2872 36193 2881 36227
rect 2881 36193 2915 36227
rect 2915 36193 2924 36227
rect 2872 36184 2924 36193
rect 8116 36227 8168 36236
rect 8116 36193 8125 36227
rect 8125 36193 8159 36227
rect 8159 36193 8168 36227
rect 8116 36184 8168 36193
rect 13360 36227 13412 36236
rect 13360 36193 13369 36227
rect 13369 36193 13403 36227
rect 13403 36193 13412 36227
rect 13360 36184 13412 36193
rect 18604 36227 18656 36236
rect 18604 36193 18613 36227
rect 18613 36193 18647 36227
rect 18647 36193 18656 36227
rect 18604 36184 18656 36193
rect 20720 36227 20772 36236
rect 20720 36193 20729 36227
rect 20729 36193 20763 36227
rect 20763 36193 20772 36227
rect 20720 36184 20772 36193
rect 25872 36184 25924 36236
rect 32864 36252 32916 36304
rect 2780 36116 2832 36168
rect 3608 36159 3660 36168
rect 3608 36125 3617 36159
rect 3617 36125 3651 36159
rect 3651 36125 3660 36159
rect 3608 36116 3660 36125
rect 4528 36116 4580 36168
rect 6552 36116 6604 36168
rect 8760 36159 8812 36168
rect 8760 36125 8769 36159
rect 8769 36125 8803 36159
rect 8803 36125 8812 36159
rect 8760 36116 8812 36125
rect 9772 36159 9824 36168
rect 9772 36125 9781 36159
rect 9781 36125 9815 36159
rect 9815 36125 9824 36159
rect 9772 36116 9824 36125
rect 12164 36116 12216 36168
rect 12440 36159 12492 36168
rect 12440 36125 12449 36159
rect 12449 36125 12483 36159
rect 12483 36125 12492 36159
rect 12440 36116 12492 36125
rect 14188 36116 14240 36168
rect 14464 36159 14516 36168
rect 14464 36125 14473 36159
rect 14473 36125 14507 36159
rect 14507 36125 14516 36159
rect 14464 36116 14516 36125
rect 17592 36159 17644 36168
rect 17592 36125 17601 36159
rect 17601 36125 17635 36159
rect 17635 36125 17644 36159
rect 17592 36116 17644 36125
rect 6736 36048 6788 36100
rect 11980 36048 12032 36100
rect 17224 36048 17276 36100
rect 19340 36116 19392 36168
rect 20812 36116 20864 36168
rect 22284 36159 22336 36168
rect 22284 36125 22293 36159
rect 22293 36125 22327 36159
rect 22327 36125 22336 36159
rect 22284 36116 22336 36125
rect 24032 36116 24084 36168
rect 25964 36159 26016 36168
rect 25964 36125 25973 36159
rect 25973 36125 26007 36159
rect 26007 36125 26016 36159
rect 25964 36116 26016 36125
rect 35348 36184 35400 36236
rect 29092 36159 29144 36168
rect 29092 36125 29101 36159
rect 29101 36125 29135 36159
rect 29135 36125 29144 36159
rect 29092 36116 29144 36125
rect 22744 36091 22796 36100
rect 22744 36057 22753 36091
rect 22753 36057 22787 36091
rect 22787 36057 22796 36091
rect 22744 36048 22796 36057
rect 24860 36091 24912 36100
rect 24860 36057 24869 36091
rect 24869 36057 24903 36091
rect 24903 36057 24912 36091
rect 24860 36048 24912 36057
rect 31576 36159 31628 36168
rect 31576 36125 31585 36159
rect 31585 36125 31619 36159
rect 31619 36125 31628 36159
rect 31576 36116 31628 36125
rect 31668 36116 31720 36168
rect 34152 36159 34204 36168
rect 34152 36125 34161 36159
rect 34161 36125 34195 36159
rect 34195 36125 34204 36159
rect 34152 36116 34204 36125
rect 35900 36159 35952 36168
rect 35900 36125 35909 36159
rect 35909 36125 35943 36159
rect 35943 36125 35952 36159
rect 35900 36116 35952 36125
rect 33692 36048 33744 36100
rect 35532 36048 35584 36100
rect 2136 35980 2188 36032
rect 4712 36023 4764 36032
rect 4712 35989 4721 36023
rect 4721 35989 4755 36023
rect 4755 35989 4764 36023
rect 4712 35980 4764 35989
rect 9220 36023 9272 36032
rect 9220 35989 9229 36023
rect 9229 35989 9263 36023
rect 9263 35989 9272 36023
rect 9220 35980 9272 35989
rect 11796 36023 11848 36032
rect 11796 35989 11805 36023
rect 11805 35989 11839 36023
rect 11839 35989 11848 36023
rect 11796 35980 11848 35989
rect 15016 36023 15068 36032
rect 15016 35989 15025 36023
rect 15025 35989 15059 36023
rect 15059 35989 15068 36023
rect 15016 35980 15068 35989
rect 19248 36023 19300 36032
rect 19248 35989 19257 36023
rect 19257 35989 19291 36023
rect 19291 35989 19300 36023
rect 19248 35980 19300 35989
rect 19432 35980 19484 36032
rect 27068 35980 27120 36032
rect 29552 35980 29604 36032
rect 33600 36023 33652 36032
rect 33600 35989 33609 36023
rect 33609 35989 33643 36023
rect 33643 35989 33652 36023
rect 33600 35980 33652 35989
rect 36176 36023 36228 36032
rect 36176 35989 36185 36023
rect 36185 35989 36219 36023
rect 36219 35989 36228 36023
rect 36176 35980 36228 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 22284 35776 22336 35828
rect 3608 35708 3660 35760
rect 4620 35708 4672 35760
rect 8760 35708 8812 35760
rect 14188 35751 14240 35760
rect 14188 35717 14197 35751
rect 14197 35717 14231 35751
rect 14231 35717 14240 35751
rect 14188 35708 14240 35717
rect 19432 35751 19484 35760
rect 19432 35717 19441 35751
rect 19441 35717 19475 35751
rect 19475 35717 19484 35751
rect 19432 35708 19484 35717
rect 20812 35751 20864 35760
rect 20812 35717 20821 35751
rect 20821 35717 20855 35751
rect 20855 35717 20864 35751
rect 20812 35708 20864 35717
rect 31668 35708 31720 35760
rect 35900 35708 35952 35760
rect 3148 35640 3200 35692
rect 3700 35683 3752 35692
rect 3700 35649 3709 35683
rect 3709 35649 3743 35683
rect 3743 35649 3752 35683
rect 3700 35640 3752 35649
rect 5724 35640 5776 35692
rect 6736 35683 6788 35692
rect 6736 35649 6745 35683
rect 6745 35649 6779 35683
rect 6779 35649 6788 35683
rect 6736 35640 6788 35649
rect 8852 35640 8904 35692
rect 10140 35683 10192 35692
rect 10140 35649 10149 35683
rect 10149 35649 10183 35683
rect 10183 35649 10192 35683
rect 10140 35640 10192 35649
rect 11980 35683 12032 35692
rect 11980 35649 11989 35683
rect 11989 35649 12023 35683
rect 12023 35649 12032 35683
rect 11980 35640 12032 35649
rect 14648 35640 14700 35692
rect 15292 35683 15344 35692
rect 15292 35649 15301 35683
rect 15301 35649 15335 35683
rect 15335 35649 15344 35683
rect 15292 35640 15344 35649
rect 17224 35683 17276 35692
rect 17224 35649 17233 35683
rect 17233 35649 17267 35683
rect 17267 35649 17276 35683
rect 17224 35640 17276 35649
rect 19984 35683 20036 35692
rect 19984 35649 19993 35683
rect 19993 35649 20027 35683
rect 20027 35649 20036 35683
rect 19984 35640 20036 35649
rect 20352 35683 20404 35692
rect 20352 35649 20361 35683
rect 20361 35649 20395 35683
rect 20395 35649 20404 35683
rect 20352 35640 20404 35649
rect 22744 35683 22796 35692
rect 22744 35649 22753 35683
rect 22753 35649 22787 35683
rect 22787 35649 22796 35683
rect 22744 35640 22796 35649
rect 24860 35640 24912 35692
rect 27528 35683 27580 35692
rect 27528 35649 27537 35683
rect 27537 35649 27571 35683
rect 27571 35649 27580 35683
rect 27528 35640 27580 35649
rect 30472 35683 30524 35692
rect 30472 35649 30481 35683
rect 30481 35649 30515 35683
rect 30515 35649 30524 35683
rect 30472 35640 30524 35649
rect 3792 35572 3844 35624
rect 6368 35572 6420 35624
rect 9864 35572 9916 35624
rect 11612 35572 11664 35624
rect 15016 35572 15068 35624
rect 16856 35572 16908 35624
rect 21916 35615 21968 35624
rect 21916 35581 21925 35615
rect 21925 35581 21959 35615
rect 21959 35581 21968 35615
rect 21916 35572 21968 35581
rect 22100 35572 22152 35624
rect 23848 35572 23900 35624
rect 24768 35504 24820 35556
rect 27344 35572 27396 35624
rect 30840 35572 30892 35624
rect 33692 35683 33744 35692
rect 33692 35649 33701 35683
rect 33701 35649 33735 35683
rect 33735 35649 33744 35683
rect 33692 35640 33744 35649
rect 32496 35504 32548 35556
rect 36636 35547 36688 35556
rect 36636 35513 36645 35547
rect 36645 35513 36679 35547
rect 36679 35513 36688 35547
rect 36636 35504 36688 35513
rect 23388 35436 23440 35488
rect 29920 35436 29972 35488
rect 36360 35479 36412 35488
rect 36360 35445 36369 35479
rect 36369 35445 36403 35479
rect 36403 35445 36412 35479
rect 36360 35436 36412 35445
rect 36544 35479 36596 35488
rect 36544 35445 36553 35479
rect 36553 35445 36587 35479
rect 36587 35445 36596 35479
rect 36544 35436 36596 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 4620 35232 4672 35284
rect 9772 35232 9824 35284
rect 12440 35232 12492 35284
rect 14464 35232 14516 35284
rect 4804 35164 4856 35216
rect 17592 35232 17644 35284
rect 19340 35232 19392 35284
rect 31576 35232 31628 35284
rect 4620 35096 4672 35148
rect 11796 35096 11848 35148
rect 14188 35139 14240 35148
rect 14188 35105 14197 35139
rect 14197 35105 14231 35139
rect 14231 35105 14240 35139
rect 14188 35096 14240 35105
rect 19248 35096 19300 35148
rect 1952 35071 2004 35080
rect 1952 35037 1961 35071
rect 1961 35037 1995 35071
rect 1995 35037 2004 35071
rect 1952 35028 2004 35037
rect 9588 35028 9640 35080
rect 2044 34960 2096 35012
rect 2964 34960 3016 35012
rect 4896 34960 4948 35012
rect 6368 34960 6420 35012
rect 7656 34960 7708 35012
rect 8944 34960 8996 35012
rect 11244 34960 11296 35012
rect 13176 34960 13228 35012
rect 22928 35028 22980 35080
rect 29920 35028 29972 35080
rect 33324 35232 33376 35284
rect 33416 35164 33468 35216
rect 36544 35232 36596 35284
rect 34520 35164 34572 35216
rect 36452 35164 36504 35216
rect 1124 34892 1176 34944
rect 3056 34892 3108 34944
rect 3884 34892 3936 34944
rect 5908 34935 5960 34944
rect 5908 34901 5917 34935
rect 5917 34901 5951 34935
rect 5951 34901 5960 34935
rect 5908 34892 5960 34901
rect 7380 34935 7432 34944
rect 7380 34901 7389 34935
rect 7389 34901 7423 34935
rect 7423 34901 7432 34935
rect 7380 34892 7432 34901
rect 11336 34892 11388 34944
rect 12072 34935 12124 34944
rect 12072 34901 12081 34935
rect 12081 34901 12115 34935
rect 12115 34901 12124 34935
rect 12072 34892 12124 34901
rect 13544 34892 13596 34944
rect 14740 34935 14792 34944
rect 14740 34901 14749 34935
rect 14749 34901 14783 34935
rect 14783 34901 14792 34935
rect 14740 34892 14792 34901
rect 16764 35003 16816 35012
rect 16764 34969 16773 35003
rect 16773 34969 16807 35003
rect 16807 34969 16816 35003
rect 16764 34960 16816 34969
rect 18972 34960 19024 35012
rect 20168 34960 20220 35012
rect 22100 34960 22152 35012
rect 23940 34960 23992 35012
rect 26148 34960 26200 35012
rect 27436 34960 27488 35012
rect 28540 34960 28592 35012
rect 30104 35003 30156 35012
rect 30104 34969 30138 35003
rect 30138 34969 30156 35003
rect 30104 34960 30156 34969
rect 31392 34960 31444 35012
rect 34520 35071 34572 35080
rect 34520 35037 34529 35071
rect 34529 35037 34563 35071
rect 34563 35037 34572 35071
rect 34520 35028 34572 35037
rect 34796 35071 34848 35080
rect 34796 35037 34805 35071
rect 34805 35037 34839 35071
rect 34839 35037 34848 35071
rect 34796 35028 34848 35037
rect 34704 34960 34756 35012
rect 35624 34960 35676 35012
rect 16856 34935 16908 34944
rect 16856 34901 16865 34935
rect 16865 34901 16899 34935
rect 16899 34901 16908 34935
rect 16856 34892 16908 34901
rect 18420 34935 18472 34944
rect 18420 34901 18429 34935
rect 18429 34901 18463 34935
rect 18463 34901 18472 34935
rect 18420 34892 18472 34901
rect 21180 34935 21232 34944
rect 21180 34901 21189 34935
rect 21189 34901 21223 34935
rect 21223 34901 21232 34935
rect 21180 34892 21232 34901
rect 24216 34935 24268 34944
rect 24216 34901 24225 34935
rect 24225 34901 24259 34935
rect 24259 34901 24268 34935
rect 24216 34892 24268 34901
rect 24860 34935 24912 34944
rect 24860 34901 24869 34935
rect 24869 34901 24903 34935
rect 24903 34901 24912 34935
rect 24860 34892 24912 34901
rect 27896 34935 27948 34944
rect 27896 34901 27905 34935
rect 27905 34901 27939 34935
rect 27939 34901 27948 34935
rect 27896 34892 27948 34901
rect 31208 34935 31260 34944
rect 31208 34901 31217 34935
rect 31217 34901 31251 34935
rect 31251 34901 31260 34935
rect 31208 34892 31260 34901
rect 32128 34892 32180 34944
rect 34152 34892 34204 34944
rect 36268 35028 36320 35080
rect 36084 35003 36136 35012
rect 36084 34969 36093 35003
rect 36093 34969 36127 35003
rect 36127 34969 36136 35003
rect 36084 34960 36136 34969
rect 36912 34935 36964 34944
rect 36912 34901 36921 34935
rect 36921 34901 36955 34935
rect 36955 34901 36964 34935
rect 36912 34892 36964 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 2044 34688 2096 34740
rect 2780 34731 2832 34740
rect 2780 34697 2789 34731
rect 2789 34697 2823 34731
rect 2823 34697 2832 34731
rect 2780 34688 2832 34697
rect 2688 34620 2740 34672
rect 5724 34688 5776 34740
rect 5908 34688 5960 34740
rect 1952 34552 2004 34604
rect 2136 34595 2188 34604
rect 2136 34561 2145 34595
rect 2145 34561 2179 34595
rect 2179 34561 2188 34595
rect 2136 34552 2188 34561
rect 3884 34595 3936 34604
rect 3884 34561 3902 34595
rect 3902 34561 3936 34595
rect 3884 34552 3936 34561
rect 6000 34595 6052 34604
rect 6000 34561 6009 34595
rect 6009 34561 6043 34595
rect 6043 34561 6052 34595
rect 6000 34552 6052 34561
rect 7380 34688 7432 34740
rect 8852 34688 8904 34740
rect 8944 34731 8996 34740
rect 8944 34697 8953 34731
rect 8953 34697 8987 34731
rect 8987 34697 8996 34731
rect 8944 34688 8996 34697
rect 11060 34688 11112 34740
rect 11244 34688 11296 34740
rect 12164 34731 12216 34740
rect 12164 34697 12173 34731
rect 12173 34697 12207 34731
rect 12207 34697 12216 34731
rect 12164 34688 12216 34697
rect 14740 34688 14792 34740
rect 15292 34688 15344 34740
rect 11336 34620 11388 34672
rect 13544 34620 13596 34672
rect 10140 34595 10192 34604
rect 10140 34561 10149 34595
rect 10149 34561 10183 34595
rect 10183 34561 10192 34595
rect 10140 34552 10192 34561
rect 10600 34595 10652 34604
rect 10600 34561 10609 34595
rect 10609 34561 10643 34595
rect 10643 34561 10652 34595
rect 10600 34552 10652 34561
rect 2964 34484 3016 34536
rect 8208 34527 8260 34536
rect 8208 34493 8217 34527
rect 8217 34493 8251 34527
rect 8251 34493 8260 34527
rect 8208 34484 8260 34493
rect 9588 34484 9640 34536
rect 2596 34416 2648 34468
rect 9220 34416 9272 34468
rect 11060 34416 11112 34468
rect 12072 34552 12124 34604
rect 14556 34552 14608 34604
rect 16856 34688 16908 34740
rect 17776 34731 17828 34740
rect 17776 34697 17785 34731
rect 17785 34697 17819 34731
rect 17819 34697 17828 34731
rect 17776 34688 17828 34697
rect 18972 34731 19024 34740
rect 18972 34697 18981 34731
rect 18981 34697 19015 34731
rect 19015 34697 19024 34731
rect 18972 34688 19024 34697
rect 19984 34688 20036 34740
rect 20168 34688 20220 34740
rect 23940 34688 23992 34740
rect 24032 34731 24084 34740
rect 24032 34697 24041 34731
rect 24041 34697 24075 34731
rect 24075 34697 24084 34731
rect 24032 34688 24084 34697
rect 24216 34688 24268 34740
rect 24768 34731 24820 34740
rect 24768 34697 24777 34731
rect 24777 34697 24811 34731
rect 24811 34697 24820 34731
rect 24768 34688 24820 34697
rect 24860 34688 24912 34740
rect 7012 34391 7064 34400
rect 7012 34357 7021 34391
rect 7021 34357 7055 34391
rect 7055 34357 7064 34391
rect 7012 34348 7064 34357
rect 8024 34391 8076 34400
rect 8024 34357 8033 34391
rect 8033 34357 8067 34391
rect 8067 34357 8076 34391
rect 8024 34348 8076 34357
rect 16856 34527 16908 34536
rect 16856 34493 16865 34527
rect 16865 34493 16899 34527
rect 16899 34493 16908 34527
rect 16856 34484 16908 34493
rect 18512 34527 18564 34536
rect 18512 34493 18521 34527
rect 18521 34493 18555 34527
rect 18555 34493 18564 34527
rect 18512 34484 18564 34493
rect 18420 34416 18472 34468
rect 22376 34620 22428 34672
rect 21180 34552 21232 34604
rect 21916 34552 21968 34604
rect 23388 34595 23440 34604
rect 23388 34561 23397 34595
rect 23397 34561 23431 34595
rect 23431 34561 23440 34595
rect 23388 34552 23440 34561
rect 26148 34688 26200 34740
rect 27528 34688 27580 34740
rect 27896 34688 27948 34740
rect 28540 34731 28592 34740
rect 28540 34697 28549 34731
rect 28549 34697 28583 34731
rect 28583 34697 28592 34731
rect 28540 34688 28592 34697
rect 29092 34688 29144 34740
rect 25412 34484 25464 34536
rect 27068 34595 27120 34604
rect 27068 34561 27077 34595
rect 27077 34561 27111 34595
rect 27111 34561 27120 34595
rect 27068 34552 27120 34561
rect 31668 34552 31720 34604
rect 31944 34595 31996 34604
rect 31944 34561 31953 34595
rect 31953 34561 31987 34595
rect 31987 34561 31996 34595
rect 31944 34552 31996 34561
rect 26608 34484 26660 34536
rect 26700 34527 26752 34536
rect 26700 34493 26709 34527
rect 26709 34493 26743 34527
rect 26743 34493 26752 34527
rect 26700 34484 26752 34493
rect 25964 34416 26016 34468
rect 29644 34484 29696 34536
rect 31392 34484 31444 34536
rect 34612 34688 34664 34740
rect 33324 34620 33376 34672
rect 34520 34620 34572 34672
rect 35348 34620 35400 34672
rect 32956 34552 33008 34604
rect 34060 34595 34112 34604
rect 34060 34561 34069 34595
rect 34069 34561 34103 34595
rect 34103 34561 34112 34595
rect 34060 34552 34112 34561
rect 36728 34552 36780 34604
rect 34336 34527 34388 34536
rect 34336 34493 34345 34527
rect 34345 34493 34379 34527
rect 34379 34493 34388 34527
rect 34336 34484 34388 34493
rect 34520 34484 34572 34536
rect 12072 34348 12124 34400
rect 13268 34391 13320 34400
rect 13268 34357 13277 34391
rect 13277 34357 13311 34391
rect 13311 34357 13320 34391
rect 13268 34348 13320 34357
rect 30932 34348 30984 34400
rect 34152 34348 34204 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 3700 34144 3752 34196
rect 6000 34144 6052 34196
rect 6552 34144 6604 34196
rect 7656 34187 7708 34196
rect 7656 34153 7665 34187
rect 7665 34153 7699 34187
rect 7699 34153 7708 34187
rect 7656 34144 7708 34153
rect 8208 34144 8260 34196
rect 10600 34187 10652 34196
rect 10600 34153 10609 34187
rect 10609 34153 10643 34187
rect 10643 34153 10652 34187
rect 10600 34144 10652 34153
rect 12072 34187 12124 34196
rect 12072 34153 12081 34187
rect 12081 34153 12115 34187
rect 12115 34153 12124 34187
rect 12072 34144 12124 34153
rect 2596 34008 2648 34060
rect 4252 34051 4304 34060
rect 4252 34017 4261 34051
rect 4261 34017 4295 34051
rect 4295 34017 4304 34051
rect 4252 34008 4304 34017
rect 4804 34008 4856 34060
rect 5264 34051 5316 34060
rect 5264 34017 5273 34051
rect 5273 34017 5307 34051
rect 5307 34017 5316 34051
rect 5264 34008 5316 34017
rect 7012 34008 7064 34060
rect 8024 34051 8076 34060
rect 8024 34017 8033 34051
rect 8033 34017 8067 34051
rect 8067 34017 8076 34051
rect 8024 34008 8076 34017
rect 9220 34008 9272 34060
rect 13176 34187 13228 34196
rect 13176 34153 13185 34187
rect 13185 34153 13219 34187
rect 13219 34153 13228 34187
rect 13176 34144 13228 34153
rect 14188 34144 14240 34196
rect 14740 34144 14792 34196
rect 22100 34144 22152 34196
rect 22928 34144 22980 34196
rect 25412 34187 25464 34196
rect 25412 34153 25421 34187
rect 25421 34153 25455 34187
rect 25455 34153 25464 34187
rect 25412 34144 25464 34153
rect 25964 34144 26016 34196
rect 27436 34187 27488 34196
rect 27436 34153 27445 34187
rect 27445 34153 27479 34187
rect 27479 34153 27488 34187
rect 27436 34144 27488 34153
rect 30104 34187 30156 34196
rect 30104 34153 30113 34187
rect 30113 34153 30147 34187
rect 30147 34153 30156 34187
rect 30104 34144 30156 34153
rect 13912 34076 13964 34128
rect 23388 34076 23440 34128
rect 13268 34051 13320 34060
rect 13268 34017 13277 34051
rect 13277 34017 13311 34051
rect 13311 34017 13320 34051
rect 13268 34008 13320 34017
rect 15016 34008 15068 34060
rect 22376 34051 22428 34060
rect 22376 34017 22385 34051
rect 22385 34017 22419 34051
rect 22419 34017 22428 34051
rect 22376 34008 22428 34017
rect 26608 34051 26660 34060
rect 26608 34017 26617 34051
rect 26617 34017 26651 34051
rect 26651 34017 26660 34051
rect 26608 34008 26660 34017
rect 30012 34119 30064 34128
rect 30012 34085 30021 34119
rect 30021 34085 30055 34119
rect 30055 34085 30064 34119
rect 30012 34076 30064 34085
rect 28724 34051 28776 34060
rect 28724 34017 28733 34051
rect 28733 34017 28767 34051
rect 28767 34017 28776 34051
rect 28724 34008 28776 34017
rect 29644 34051 29696 34060
rect 29644 34017 29653 34051
rect 29653 34017 29687 34051
rect 29687 34017 29696 34051
rect 32404 34144 32456 34196
rect 35256 34144 35308 34196
rect 35440 34144 35492 34196
rect 29644 34008 29696 34017
rect 3240 33940 3292 33992
rect 3792 33983 3844 33992
rect 3792 33949 3801 33983
rect 3801 33949 3835 33983
rect 3835 33949 3844 33983
rect 3792 33940 3844 33949
rect 4896 33940 4948 33992
rect 6828 33940 6880 33992
rect 28080 33983 28132 33992
rect 28080 33949 28089 33983
rect 28089 33949 28123 33983
rect 28123 33949 28132 33983
rect 28080 33940 28132 33949
rect 30472 33940 30524 33992
rect 33416 34008 33468 34060
rect 35716 34076 35768 34128
rect 35808 34008 35860 34060
rect 36176 34076 36228 34128
rect 36360 34076 36412 34128
rect 31760 33983 31812 33992
rect 31760 33949 31769 33983
rect 31769 33949 31803 33983
rect 31803 33949 31812 33983
rect 31760 33940 31812 33949
rect 33232 33983 33284 33992
rect 33232 33949 33241 33983
rect 33241 33949 33275 33983
rect 33275 33949 33284 33983
rect 33232 33940 33284 33949
rect 34612 33940 34664 33992
rect 2872 33804 2924 33856
rect 17316 33804 17368 33856
rect 18512 33804 18564 33856
rect 26700 33804 26752 33856
rect 27988 33804 28040 33856
rect 29184 33804 29236 33856
rect 30656 33804 30708 33856
rect 33600 33915 33652 33924
rect 33600 33881 33609 33915
rect 33609 33881 33643 33915
rect 33643 33881 33652 33915
rect 33600 33872 33652 33881
rect 34428 33804 34480 33856
rect 35716 33872 35768 33924
rect 36544 33915 36596 33924
rect 36544 33881 36553 33915
rect 36553 33881 36587 33915
rect 36587 33881 36596 33915
rect 36544 33872 36596 33881
rect 34704 33804 34756 33856
rect 35532 33804 35584 33856
rect 36268 33804 36320 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 5264 33600 5316 33652
rect 6368 33643 6420 33652
rect 6368 33609 6377 33643
rect 6377 33609 6411 33643
rect 6411 33609 6420 33643
rect 6368 33600 6420 33609
rect 6828 33600 6880 33652
rect 12072 33600 12124 33652
rect 2504 33464 2556 33516
rect 2872 33507 2924 33516
rect 2872 33473 2881 33507
rect 2881 33473 2915 33507
rect 2915 33473 2924 33507
rect 2872 33464 2924 33473
rect 4712 33507 4764 33516
rect 4712 33473 4721 33507
rect 4721 33473 4755 33507
rect 4755 33473 4764 33507
rect 4712 33464 4764 33473
rect 2596 33396 2648 33448
rect 3332 33439 3384 33448
rect 3332 33405 3341 33439
rect 3341 33405 3375 33439
rect 3375 33405 3384 33439
rect 3332 33396 3384 33405
rect 6000 33439 6052 33448
rect 6000 33405 6009 33439
rect 6009 33405 6043 33439
rect 6043 33405 6052 33439
rect 6000 33396 6052 33405
rect 13912 33600 13964 33652
rect 14556 33600 14608 33652
rect 14648 33464 14700 33516
rect 16856 33600 16908 33652
rect 17316 33600 17368 33652
rect 28724 33600 28776 33652
rect 29644 33600 29696 33652
rect 31760 33600 31812 33652
rect 27988 33575 28040 33584
rect 27988 33541 27997 33575
rect 27997 33541 28031 33575
rect 28031 33541 28040 33575
rect 27988 33532 28040 33541
rect 33140 33600 33192 33652
rect 31944 33532 31996 33584
rect 28080 33464 28132 33516
rect 29552 33507 29604 33516
rect 29552 33473 29561 33507
rect 29561 33473 29595 33507
rect 29595 33473 29604 33507
rect 29552 33464 29604 33473
rect 30932 33464 30984 33516
rect 31208 33464 31260 33516
rect 32404 33507 32456 33516
rect 32404 33473 32413 33507
rect 32413 33473 32447 33507
rect 32447 33473 32456 33507
rect 32404 33464 32456 33473
rect 32588 33507 32640 33516
rect 32588 33473 32597 33507
rect 32597 33473 32631 33507
rect 32631 33473 32640 33507
rect 32588 33464 32640 33473
rect 6552 33371 6604 33380
rect 6552 33337 6561 33371
rect 6561 33337 6595 33371
rect 6595 33337 6604 33371
rect 6552 33328 6604 33337
rect 14740 33371 14792 33380
rect 14740 33337 14749 33371
rect 14749 33337 14783 33371
rect 14783 33337 14792 33371
rect 14740 33328 14792 33337
rect 30656 33439 30708 33448
rect 30656 33405 30665 33439
rect 30665 33405 30699 33439
rect 30699 33405 30708 33439
rect 30656 33396 30708 33405
rect 35532 33600 35584 33652
rect 35716 33600 35768 33652
rect 35900 33600 35952 33652
rect 36176 33600 36228 33652
rect 36912 33532 36964 33584
rect 33968 33464 34020 33516
rect 35348 33507 35400 33516
rect 35348 33473 35357 33507
rect 35357 33473 35391 33507
rect 35391 33473 35400 33507
rect 35348 33464 35400 33473
rect 4712 33260 4764 33312
rect 34152 33260 34204 33312
rect 34704 33260 34756 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 32496 33099 32548 33108
rect 32496 33065 32505 33099
rect 32505 33065 32539 33099
rect 32539 33065 32548 33099
rect 32496 33056 32548 33065
rect 32956 33056 33008 33108
rect 1584 32963 1636 32972
rect 1584 32929 1593 32963
rect 1593 32929 1627 32963
rect 1627 32929 1636 32963
rect 1584 32920 1636 32929
rect 29184 32920 29236 32972
rect 32404 32988 32456 33040
rect 32772 32988 32824 33040
rect 33324 32988 33376 33040
rect 34244 32963 34296 32972
rect 34244 32929 34253 32963
rect 34253 32929 34287 32963
rect 34287 32929 34296 32963
rect 34244 32920 34296 32929
rect 2596 32895 2648 32904
rect 2596 32861 2605 32895
rect 2605 32861 2639 32895
rect 2639 32861 2648 32895
rect 2596 32852 2648 32861
rect 3792 32852 3844 32904
rect 6276 32852 6328 32904
rect 4528 32827 4580 32836
rect 4528 32793 4537 32827
rect 4537 32793 4571 32827
rect 4571 32793 4580 32827
rect 4528 32784 4580 32793
rect 3516 32759 3568 32768
rect 3516 32725 3525 32759
rect 3525 32725 3559 32759
rect 3559 32725 3568 32759
rect 3516 32716 3568 32725
rect 30288 32759 30340 32768
rect 30288 32725 30297 32759
rect 30297 32725 30331 32759
rect 30331 32725 30340 32759
rect 30288 32716 30340 32725
rect 32036 32852 32088 32904
rect 32312 32852 32364 32904
rect 33600 32852 33652 32904
rect 36084 33056 36136 33108
rect 36360 33056 36412 33108
rect 31944 32784 31996 32836
rect 34244 32784 34296 32836
rect 36176 32852 36228 32904
rect 36268 32895 36320 32904
rect 36268 32861 36277 32895
rect 36277 32861 36311 32895
rect 36311 32861 36320 32895
rect 36268 32852 36320 32861
rect 34520 32716 34572 32768
rect 35532 32784 35584 32836
rect 37188 32827 37240 32836
rect 37188 32793 37197 32827
rect 37197 32793 37231 32827
rect 37231 32793 37240 32827
rect 37188 32784 37240 32793
rect 35440 32716 35492 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 4528 32512 4580 32564
rect 6000 32512 6052 32564
rect 33232 32512 33284 32564
rect 3056 32487 3108 32496
rect 3056 32453 3065 32487
rect 3065 32453 3099 32487
rect 3099 32453 3108 32487
rect 3056 32444 3108 32453
rect 2596 32419 2648 32428
rect 2596 32385 2605 32419
rect 2605 32385 2639 32419
rect 2639 32385 2648 32419
rect 2596 32376 2648 32385
rect 34244 32444 34296 32496
rect 36544 32512 36596 32564
rect 4620 32376 4672 32428
rect 34336 32376 34388 32428
rect 36084 32444 36136 32496
rect 36360 32444 36412 32496
rect 36820 32444 36872 32496
rect 35808 32419 35860 32428
rect 35808 32385 35817 32419
rect 35817 32385 35851 32419
rect 35851 32385 35860 32419
rect 35808 32376 35860 32385
rect 1584 32351 1636 32360
rect 1584 32317 1593 32351
rect 1593 32317 1627 32351
rect 1627 32317 1636 32351
rect 1584 32308 1636 32317
rect 30656 32351 30708 32360
rect 30656 32317 30665 32351
rect 30665 32317 30699 32351
rect 30699 32317 30708 32351
rect 30656 32308 30708 32317
rect 30288 32240 30340 32292
rect 33692 32351 33744 32360
rect 33692 32317 33701 32351
rect 33701 32317 33735 32351
rect 33735 32317 33744 32351
rect 33692 32308 33744 32317
rect 35716 32308 35768 32360
rect 36636 32240 36688 32292
rect 33968 32172 34020 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 2596 31968 2648 32020
rect 30288 31968 30340 32020
rect 30656 31968 30708 32020
rect 32588 31968 32640 32020
rect 33324 31968 33376 32020
rect 32128 31875 32180 31884
rect 32128 31841 32137 31875
rect 32137 31841 32171 31875
rect 32171 31841 32180 31875
rect 32128 31832 32180 31841
rect 2780 31764 2832 31816
rect 2964 31807 3016 31816
rect 2964 31773 2973 31807
rect 2973 31773 3007 31807
rect 3007 31773 3016 31807
rect 2964 31764 3016 31773
rect 8116 31807 8168 31816
rect 8116 31773 8125 31807
rect 8125 31773 8159 31807
rect 8159 31773 8168 31807
rect 8116 31764 8168 31773
rect 10876 31764 10928 31816
rect 32772 31764 32824 31816
rect 34796 31968 34848 32020
rect 35440 31968 35492 32020
rect 36176 31968 36228 32020
rect 36728 31900 36780 31952
rect 37004 31943 37056 31952
rect 37004 31909 37013 31943
rect 37013 31909 37047 31943
rect 37047 31909 37056 31943
rect 37004 31900 37056 31909
rect 34612 31832 34664 31884
rect 35348 31832 35400 31884
rect 36820 31832 36872 31884
rect 34796 31807 34848 31816
rect 34796 31773 34805 31807
rect 34805 31773 34839 31807
rect 34839 31773 34848 31807
rect 34796 31764 34848 31773
rect 35532 31764 35584 31816
rect 4436 31671 4488 31680
rect 4436 31637 4445 31671
rect 4445 31637 4479 31671
rect 4479 31637 4488 31671
rect 4436 31628 4488 31637
rect 34244 31628 34296 31680
rect 34612 31628 34664 31680
rect 35532 31628 35584 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 2780 31424 2832 31476
rect 35808 31424 35860 31476
rect 36820 31467 36872 31476
rect 36820 31433 36829 31467
rect 36829 31433 36863 31467
rect 36863 31433 36872 31467
rect 36820 31424 36872 31433
rect 2596 31331 2648 31340
rect 2596 31297 2605 31331
rect 2605 31297 2639 31331
rect 2639 31297 2648 31331
rect 2596 31288 2648 31297
rect 4436 31288 4488 31340
rect 4620 31288 4672 31340
rect 31944 31288 31996 31340
rect 35440 31331 35492 31340
rect 35440 31297 35449 31331
rect 35449 31297 35483 31331
rect 35483 31297 35492 31331
rect 35440 31288 35492 31297
rect 35532 31288 35584 31340
rect 1584 31263 1636 31272
rect 1584 31229 1593 31263
rect 1593 31229 1627 31263
rect 1627 31229 1636 31263
rect 1584 31220 1636 31229
rect 2872 31263 2924 31272
rect 2872 31229 2881 31263
rect 2881 31229 2915 31263
rect 2915 31229 2924 31263
rect 2872 31220 2924 31229
rect 33508 31263 33560 31272
rect 33508 31229 33517 31263
rect 33517 31229 33551 31263
rect 33551 31229 33560 31263
rect 33508 31220 33560 31229
rect 36268 31399 36320 31408
rect 36268 31365 36277 31399
rect 36277 31365 36311 31399
rect 36311 31365 36320 31399
rect 36268 31356 36320 31365
rect 33416 31195 33468 31204
rect 33416 31161 33425 31195
rect 33425 31161 33459 31195
rect 33459 31161 33468 31195
rect 37004 31220 37056 31272
rect 33416 31152 33468 31161
rect 4068 31084 4120 31136
rect 37832 31152 37884 31204
rect 36452 31084 36504 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 2596 30880 2648 30932
rect 2872 30923 2924 30932
rect 2872 30889 2881 30923
rect 2881 30889 2915 30923
rect 2915 30889 2924 30923
rect 2872 30880 2924 30889
rect 3240 30880 3292 30932
rect 33416 30880 33468 30932
rect 34060 30880 34112 30932
rect 4620 30855 4672 30864
rect 4620 30821 4629 30855
rect 4629 30821 4663 30855
rect 4663 30821 4672 30855
rect 4620 30812 4672 30821
rect 4896 30744 4948 30796
rect 32404 30744 32456 30796
rect 34796 30812 34848 30864
rect 34704 30744 34756 30796
rect 3056 30676 3108 30728
rect 3424 30719 3476 30728
rect 3424 30685 3433 30719
rect 3433 30685 3467 30719
rect 3467 30685 3476 30719
rect 3424 30676 3476 30685
rect 4712 30676 4764 30728
rect 35256 30676 35308 30728
rect 35992 30719 36044 30728
rect 35992 30685 36001 30719
rect 36001 30685 36035 30719
rect 36035 30685 36044 30719
rect 35992 30676 36044 30685
rect 36268 30719 36320 30728
rect 36268 30685 36277 30719
rect 36277 30685 36311 30719
rect 36311 30685 36320 30719
rect 36268 30676 36320 30685
rect 34796 30651 34848 30660
rect 34796 30617 34805 30651
rect 34805 30617 34839 30651
rect 34839 30617 34848 30651
rect 34796 30608 34848 30617
rect 37188 30651 37240 30660
rect 37188 30617 37197 30651
rect 37197 30617 37231 30651
rect 37231 30617 37240 30651
rect 37188 30608 37240 30617
rect 4620 30540 4672 30592
rect 35532 30540 35584 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 3056 30336 3108 30388
rect 35992 30336 36044 30388
rect 2688 30200 2740 30252
rect 3240 30200 3292 30252
rect 34520 30268 34572 30320
rect 35532 30268 35584 30320
rect 33140 30200 33192 30252
rect 35256 30243 35308 30252
rect 35256 30209 35265 30243
rect 35265 30209 35299 30243
rect 35299 30209 35308 30243
rect 35256 30200 35308 30209
rect 35348 30200 35400 30252
rect 4068 30175 4120 30184
rect 4068 30141 4077 30175
rect 4077 30141 4111 30175
rect 4111 30141 4120 30175
rect 4068 30132 4120 30141
rect 2964 29996 3016 30048
rect 34704 30039 34756 30048
rect 34704 30005 34713 30039
rect 34713 30005 34747 30039
rect 34747 30005 34756 30039
rect 34704 29996 34756 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 3424 29792 3476 29844
rect 3792 29835 3844 29844
rect 3792 29801 3801 29835
rect 3801 29801 3835 29835
rect 3835 29801 3844 29835
rect 3792 29792 3844 29801
rect 6276 29835 6328 29844
rect 6276 29801 6285 29835
rect 6285 29801 6319 29835
rect 6319 29801 6328 29835
rect 6276 29792 6328 29801
rect 10876 29835 10928 29844
rect 10876 29801 10885 29835
rect 10885 29801 10919 29835
rect 10919 29801 10928 29835
rect 10876 29792 10928 29801
rect 34704 29792 34756 29844
rect 34796 29792 34848 29844
rect 35716 29792 35768 29844
rect 6920 29699 6972 29708
rect 6920 29665 6929 29699
rect 6929 29665 6963 29699
rect 6963 29665 6972 29699
rect 6920 29656 6972 29665
rect 8116 29656 8168 29708
rect 36268 29656 36320 29708
rect 2688 29588 2740 29640
rect 3792 29588 3844 29640
rect 4620 29588 4672 29640
rect 13452 29588 13504 29640
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 3240 29248 3292 29300
rect 32772 29291 32824 29300
rect 32772 29257 32781 29291
rect 32781 29257 32815 29291
rect 32815 29257 32824 29291
rect 32772 29248 32824 29257
rect 34704 29248 34756 29300
rect 4896 29180 4948 29232
rect 2780 29112 2832 29164
rect 4068 29112 4120 29164
rect 30380 29155 30432 29164
rect 1584 29087 1636 29096
rect 1584 29053 1593 29087
rect 1593 29053 1627 29087
rect 1627 29053 1636 29087
rect 1584 29044 1636 29053
rect 4160 29087 4212 29096
rect 4160 29053 4169 29087
rect 4169 29053 4203 29087
rect 4203 29053 4212 29087
rect 4160 29044 4212 29053
rect 4620 28976 4672 29028
rect 20444 29087 20496 29096
rect 20444 29053 20453 29087
rect 20453 29053 20487 29087
rect 20487 29053 20496 29087
rect 20444 29044 20496 29053
rect 30380 29121 30389 29155
rect 30389 29121 30423 29155
rect 30423 29121 30432 29155
rect 30380 29112 30432 29121
rect 34612 29112 34664 29164
rect 32128 29087 32180 29096
rect 32128 29053 32137 29087
rect 32137 29053 32171 29087
rect 32171 29053 32180 29087
rect 32128 29044 32180 29053
rect 28448 29019 28500 29028
rect 28448 28985 28457 29019
rect 28457 28985 28491 29019
rect 28491 28985 28500 29019
rect 28448 28976 28500 28985
rect 29920 28976 29972 29028
rect 36084 29112 36136 29164
rect 34796 28976 34848 29028
rect 36912 29087 36964 29096
rect 36912 29053 36921 29087
rect 36921 29053 36955 29087
rect 36955 29053 36964 29087
rect 36912 29044 36964 29053
rect 36820 28976 36872 29028
rect 3884 28908 3936 28960
rect 4896 28951 4948 28960
rect 4896 28917 4905 28951
rect 4905 28917 4939 28951
rect 4939 28917 4948 28951
rect 4896 28908 4948 28917
rect 19248 28908 19300 28960
rect 35532 28908 35584 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 4068 28704 4120 28756
rect 20352 28704 20404 28756
rect 30380 28704 30432 28756
rect 1952 28543 2004 28552
rect 1952 28509 1961 28543
rect 1961 28509 1995 28543
rect 1995 28509 2004 28543
rect 1952 28500 2004 28509
rect 2688 28500 2740 28552
rect 3884 28543 3936 28552
rect 3884 28509 3893 28543
rect 3893 28509 3927 28543
rect 3927 28509 3936 28543
rect 3884 28500 3936 28509
rect 4896 28500 4948 28552
rect 19248 28543 19300 28552
rect 19248 28509 19257 28543
rect 19257 28509 19291 28543
rect 19291 28509 19300 28543
rect 19248 28500 19300 28509
rect 35348 28704 35400 28756
rect 36820 28747 36872 28756
rect 36820 28713 36829 28747
rect 36829 28713 36863 28747
rect 36863 28713 36872 28747
rect 36820 28704 36872 28713
rect 35164 28500 35216 28552
rect 35532 28500 35584 28552
rect 4436 28407 4488 28416
rect 4436 28373 4445 28407
rect 4445 28373 4479 28407
rect 4479 28373 4488 28407
rect 4436 28364 4488 28373
rect 35532 28364 35584 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 4436 28160 4488 28212
rect 35532 28160 35584 28212
rect 2780 28092 2832 28144
rect 2596 28067 2648 28076
rect 2596 28033 2605 28067
rect 2605 28033 2639 28067
rect 2639 28033 2648 28067
rect 2596 28024 2648 28033
rect 34796 28024 34848 28076
rect 36084 28092 36136 28144
rect 1584 27999 1636 28008
rect 1584 27965 1593 27999
rect 1593 27965 1627 27999
rect 1627 27965 1636 27999
rect 1584 27956 1636 27965
rect 35164 27956 35216 28008
rect 35440 27956 35492 28008
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 2504 27548 2556 27600
rect 3884 27548 3936 27600
rect 35440 27548 35492 27600
rect 2596 27480 2648 27532
rect 4988 27523 5040 27532
rect 4988 27489 4997 27523
rect 4997 27489 5031 27523
rect 5031 27489 5040 27523
rect 4988 27480 5040 27489
rect 34520 27523 34572 27532
rect 34520 27489 34529 27523
rect 34529 27489 34563 27523
rect 34563 27489 34572 27523
rect 34520 27480 34572 27489
rect 35808 27480 35860 27532
rect 4344 27412 4396 27464
rect 4620 27412 4672 27464
rect 35992 27455 36044 27464
rect 35992 27421 36001 27455
rect 36001 27421 36035 27455
rect 36035 27421 36044 27455
rect 35992 27412 36044 27421
rect 36268 27455 36320 27464
rect 36268 27421 36277 27455
rect 36277 27421 36311 27455
rect 36311 27421 36320 27455
rect 36268 27412 36320 27421
rect 3240 27344 3292 27396
rect 35532 27344 35584 27396
rect 37280 27387 37332 27396
rect 37280 27353 37289 27387
rect 37289 27353 37323 27387
rect 37323 27353 37332 27387
rect 37280 27344 37332 27353
rect 35440 27276 35492 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 3148 27072 3200 27124
rect 3792 27072 3844 27124
rect 4344 27072 4396 27124
rect 4620 27072 4672 27124
rect 13452 27115 13504 27124
rect 13452 27081 13461 27115
rect 13461 27081 13495 27115
rect 13495 27081 13504 27115
rect 13452 27072 13504 27081
rect 4988 27004 5040 27056
rect 1952 26979 2004 26988
rect 1952 26945 1961 26979
rect 1961 26945 1995 26979
rect 1995 26945 2004 26979
rect 1952 26936 2004 26945
rect 3332 26936 3384 26988
rect 3516 26936 3568 26988
rect 3976 26979 4028 26988
rect 3976 26945 3985 26979
rect 3985 26945 4019 26979
rect 4019 26945 4028 26979
rect 3976 26936 4028 26945
rect 9588 27004 9640 27056
rect 4068 26868 4120 26920
rect 4896 26911 4948 26920
rect 4896 26877 4905 26911
rect 4905 26877 4939 26911
rect 4939 26877 4948 26911
rect 4896 26868 4948 26877
rect 8300 26868 8352 26920
rect 35440 27072 35492 27124
rect 35532 27072 35584 27124
rect 35992 27072 36044 27124
rect 19248 27004 19300 27056
rect 35348 26936 35400 26988
rect 17316 26732 17368 26784
rect 17868 26775 17920 26784
rect 17868 26741 17877 26775
rect 17877 26741 17911 26775
rect 17911 26741 17920 26775
rect 17868 26732 17920 26741
rect 34704 26775 34756 26784
rect 34704 26741 34713 26775
rect 34713 26741 34747 26775
rect 34747 26741 34756 26775
rect 34704 26732 34756 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 3332 26528 3384 26580
rect 4896 26528 4948 26580
rect 33508 26528 33560 26580
rect 36268 26528 36320 26580
rect 1952 26435 2004 26444
rect 1952 26401 1961 26435
rect 1961 26401 1995 26435
rect 1995 26401 2004 26435
rect 1952 26392 2004 26401
rect 34704 26392 34756 26444
rect 3240 26324 3292 26376
rect 4804 26324 4856 26376
rect 6920 26324 6972 26376
rect 29000 26324 29052 26376
rect 8392 26256 8444 26308
rect 17316 26299 17368 26308
rect 17316 26265 17325 26299
rect 17325 26265 17359 26299
rect 17359 26265 17368 26299
rect 17316 26256 17368 26265
rect 34520 26188 34572 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 8300 26027 8352 26036
rect 8300 25993 8309 26027
rect 8309 25993 8343 26027
rect 8343 25993 8352 26027
rect 8300 25984 8352 25993
rect 20352 26027 20404 26036
rect 20352 25993 20361 26027
rect 20361 25993 20395 26027
rect 20395 25993 20404 26027
rect 20352 25984 20404 25993
rect 2780 25848 2832 25900
rect 8392 25848 8444 25900
rect 940 25780 992 25832
rect 3700 25780 3752 25832
rect 4804 25823 4856 25832
rect 4804 25789 4813 25823
rect 4813 25789 4847 25823
rect 4847 25789 4856 25823
rect 4804 25780 4856 25789
rect 4620 25712 4672 25764
rect 4988 25755 5040 25764
rect 4988 25721 4997 25755
rect 4997 25721 5031 25755
rect 5031 25721 5040 25755
rect 4988 25712 5040 25721
rect 35900 25891 35952 25900
rect 35900 25857 35909 25891
rect 35909 25857 35943 25891
rect 35943 25857 35952 25891
rect 35900 25848 35952 25857
rect 19432 25780 19484 25832
rect 34520 25780 34572 25832
rect 35624 25823 35676 25832
rect 35624 25789 35633 25823
rect 35633 25789 35667 25823
rect 35667 25789 35676 25823
rect 35624 25780 35676 25789
rect 37464 25780 37516 25832
rect 20260 25712 20312 25764
rect 28448 25712 28500 25764
rect 34704 25755 34756 25764
rect 34704 25721 34713 25755
rect 34713 25721 34747 25755
rect 34747 25721 34756 25755
rect 34704 25712 34756 25721
rect 34796 25712 34848 25764
rect 3792 25644 3844 25696
rect 4712 25644 4764 25696
rect 4896 25687 4948 25696
rect 4896 25653 4905 25687
rect 4905 25653 4939 25687
rect 4939 25653 4948 25687
rect 4896 25644 4948 25653
rect 35348 25644 35400 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 3700 25440 3752 25492
rect 4896 25440 4948 25492
rect 32128 25440 32180 25492
rect 35348 25440 35400 25492
rect 35624 25440 35676 25492
rect 1952 25279 2004 25288
rect 1952 25245 1961 25279
rect 1961 25245 1995 25279
rect 1995 25245 2004 25279
rect 1952 25236 2004 25245
rect 3792 25279 3844 25288
rect 3792 25245 3801 25279
rect 3801 25245 3835 25279
rect 3835 25245 3844 25279
rect 3792 25236 3844 25245
rect 4160 25236 4212 25288
rect 29644 25236 29696 25288
rect 35164 25236 35216 25288
rect 35440 25279 35492 25288
rect 35440 25245 35449 25279
rect 35449 25245 35483 25279
rect 35483 25245 35492 25279
rect 35440 25236 35492 25245
rect 4436 25143 4488 25152
rect 4436 25109 4445 25143
rect 4445 25109 4479 25143
rect 4479 25109 4488 25143
rect 4436 25100 4488 25109
rect 35348 25143 35400 25152
rect 35348 25109 35357 25143
rect 35357 25109 35391 25143
rect 35391 25109 35400 25143
rect 35348 25100 35400 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 35164 24896 35216 24948
rect 35532 24896 35584 24948
rect 2780 24828 2832 24880
rect 35900 24828 35952 24880
rect 2596 24803 2648 24812
rect 2596 24769 2605 24803
rect 2605 24769 2639 24803
rect 2639 24769 2648 24803
rect 2596 24760 2648 24769
rect 4436 24760 4488 24812
rect 34796 24760 34848 24812
rect 35348 24760 35400 24812
rect 940 24692 992 24744
rect 4620 24692 4672 24744
rect 4804 24735 4856 24744
rect 4804 24701 4813 24735
rect 4813 24701 4847 24735
rect 4847 24701 4856 24735
rect 4804 24692 4856 24701
rect 4160 24624 4212 24676
rect 3240 24556 3292 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 35532 24284 35584 24336
rect 2780 24148 2832 24200
rect 3792 24191 3844 24200
rect 3792 24157 3801 24191
rect 3801 24157 3835 24191
rect 3835 24157 3844 24191
rect 3792 24148 3844 24157
rect 4712 24148 4764 24200
rect 35992 24191 36044 24200
rect 35992 24157 36001 24191
rect 36001 24157 36035 24191
rect 36035 24157 36044 24191
rect 35992 24148 36044 24157
rect 36268 24191 36320 24200
rect 36268 24157 36277 24191
rect 36277 24157 36311 24191
rect 36311 24157 36320 24191
rect 36268 24148 36320 24157
rect 34520 24123 34572 24132
rect 34520 24089 34529 24123
rect 34529 24089 34563 24123
rect 34563 24089 34572 24123
rect 34520 24080 34572 24089
rect 36084 24080 36136 24132
rect 37280 24123 37332 24132
rect 37280 24089 37289 24123
rect 37289 24089 37323 24123
rect 37323 24089 37332 24123
rect 37280 24080 37332 24089
rect 2964 24012 3016 24064
rect 4436 24055 4488 24064
rect 4436 24021 4445 24055
rect 4445 24021 4479 24055
rect 4479 24021 4488 24055
rect 4436 24012 4488 24021
rect 35256 24055 35308 24064
rect 35256 24021 35265 24055
rect 35265 24021 35299 24055
rect 35299 24021 35308 24055
rect 35256 24012 35308 24021
rect 35348 24055 35400 24064
rect 35348 24021 35357 24055
rect 35357 24021 35391 24055
rect 35391 24021 35400 24055
rect 35348 24012 35400 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 3240 23808 3292 23860
rect 3792 23808 3844 23860
rect 4068 23851 4120 23860
rect 4068 23817 4077 23851
rect 4077 23817 4111 23851
rect 4111 23817 4120 23851
rect 4068 23808 4120 23817
rect 4436 23808 4488 23860
rect 35256 23808 35308 23860
rect 35348 23740 35400 23792
rect 35992 23808 36044 23860
rect 1952 23647 2004 23656
rect 1952 23613 1961 23647
rect 1961 23613 1995 23647
rect 1995 23613 2004 23647
rect 1952 23604 2004 23613
rect 3424 23647 3476 23656
rect 3424 23613 3433 23647
rect 3433 23613 3467 23647
rect 3467 23613 3476 23647
rect 3424 23604 3476 23613
rect 35440 23647 35492 23656
rect 35440 23613 35449 23647
rect 35449 23613 35483 23647
rect 35483 23613 35492 23647
rect 35440 23604 35492 23613
rect 2688 23468 2740 23520
rect 4068 23468 4120 23520
rect 35624 23468 35676 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 2596 23128 2648 23180
rect 4068 23264 4120 23316
rect 29000 23307 29052 23316
rect 29000 23273 29009 23307
rect 29009 23273 29043 23307
rect 29043 23273 29052 23307
rect 29000 23264 29052 23273
rect 36268 23128 36320 23180
rect 28356 23103 28408 23112
rect 28356 23069 28365 23103
rect 28365 23069 28399 23103
rect 28399 23069 28408 23103
rect 28356 23060 28408 23069
rect 35624 23060 35676 23112
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 36084 22763 36136 22772
rect 36084 22729 36093 22763
rect 36093 22729 36127 22763
rect 36127 22729 36136 22763
rect 36084 22720 36136 22729
rect 2596 22627 2648 22636
rect 2596 22593 2605 22627
rect 2605 22593 2639 22627
rect 2639 22593 2648 22627
rect 2596 22584 2648 22593
rect 1584 22559 1636 22568
rect 1584 22525 1593 22559
rect 1593 22525 1627 22559
rect 1627 22525 1636 22559
rect 1584 22516 1636 22525
rect 2964 22516 3016 22568
rect 4068 22559 4120 22568
rect 4068 22525 4077 22559
rect 4077 22525 4111 22559
rect 4111 22525 4120 22559
rect 4068 22516 4120 22525
rect 4620 22516 4672 22568
rect 36452 22559 36504 22568
rect 36452 22525 36461 22559
rect 36461 22525 36495 22559
rect 36495 22525 36504 22559
rect 36452 22516 36504 22525
rect 4160 22448 4212 22500
rect 2872 22423 2924 22432
rect 2872 22389 2881 22423
rect 2881 22389 2915 22423
rect 2915 22389 2924 22423
rect 2872 22380 2924 22389
rect 3608 22423 3660 22432
rect 3608 22389 3617 22423
rect 3617 22389 3651 22423
rect 3651 22389 3660 22423
rect 3608 22380 3660 22389
rect 37096 22423 37148 22432
rect 37096 22389 37105 22423
rect 37105 22389 37139 22423
rect 37139 22389 37148 22423
rect 37096 22380 37148 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 35624 22151 35676 22160
rect 35624 22117 35633 22151
rect 35633 22117 35667 22151
rect 35667 22117 35676 22151
rect 35624 22108 35676 22117
rect 36084 22040 36136 22092
rect 2780 21972 2832 22024
rect 3608 21972 3660 22024
rect 2964 21904 3016 21956
rect 19432 21972 19484 22024
rect 3792 21879 3844 21888
rect 3792 21845 3801 21879
rect 3801 21845 3835 21879
rect 3835 21845 3844 21879
rect 3792 21836 3844 21845
rect 4620 21836 4672 21888
rect 20352 21904 20404 21956
rect 24124 21972 24176 22024
rect 36544 21947 36596 21956
rect 36544 21913 36553 21947
rect 36553 21913 36587 21947
rect 36587 21913 36596 21947
rect 36544 21904 36596 21913
rect 28172 21836 28224 21888
rect 35532 21879 35584 21888
rect 35532 21845 35541 21879
rect 35541 21845 35575 21879
rect 35575 21845 35584 21879
rect 35532 21836 35584 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 3792 21632 3844 21684
rect 29644 21675 29696 21684
rect 29644 21641 29653 21675
rect 29653 21641 29687 21675
rect 29687 21641 29696 21675
rect 29644 21632 29696 21641
rect 29920 21675 29972 21684
rect 29920 21641 29929 21675
rect 29929 21641 29963 21675
rect 29963 21641 29972 21675
rect 29920 21632 29972 21641
rect 2596 21564 2648 21616
rect 28172 21564 28224 21616
rect 2872 21539 2924 21548
rect 2872 21505 2881 21539
rect 2881 21505 2915 21539
rect 2915 21505 2924 21539
rect 2872 21496 2924 21505
rect 36544 21632 36596 21684
rect 37464 21564 37516 21616
rect 4068 21471 4120 21480
rect 4068 21437 4077 21471
rect 4077 21437 4111 21471
rect 4111 21437 4120 21471
rect 4068 21428 4120 21437
rect 4620 21428 4672 21480
rect 27528 21428 27580 21480
rect 3976 21360 4028 21412
rect 3608 21335 3660 21344
rect 3608 21301 3617 21335
rect 3617 21301 3651 21335
rect 3651 21301 3660 21335
rect 3608 21292 3660 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 4620 21063 4672 21072
rect 4620 21029 4629 21063
rect 4629 21029 4663 21063
rect 4663 21029 4672 21063
rect 4620 21020 4672 21029
rect 4068 20952 4120 21004
rect 35440 20995 35492 21004
rect 35440 20961 35449 20995
rect 35449 20961 35483 20995
rect 35483 20961 35492 20995
rect 35440 20952 35492 20961
rect 2872 20884 2924 20936
rect 4344 20927 4396 20936
rect 4344 20893 4353 20927
rect 4353 20893 4387 20927
rect 4387 20893 4396 20927
rect 4344 20884 4396 20893
rect 35532 20884 35584 20936
rect 2596 20816 2648 20868
rect 36452 20816 36504 20868
rect 3516 20791 3568 20800
rect 3516 20757 3525 20791
rect 3525 20757 3559 20791
rect 3559 20757 3568 20791
rect 3516 20748 3568 20757
rect 4528 20791 4580 20800
rect 4528 20757 4537 20791
rect 4537 20757 4571 20791
rect 4571 20757 4580 20791
rect 4528 20748 4580 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 2872 20544 2924 20596
rect 20352 20544 20404 20596
rect 2780 20476 2832 20528
rect 4528 20476 4580 20528
rect 1952 20383 2004 20392
rect 1952 20349 1961 20383
rect 1961 20349 1995 20383
rect 1995 20349 2004 20383
rect 1952 20340 2004 20349
rect 3516 20340 3568 20392
rect 4344 20340 4396 20392
rect 22008 20272 22060 20324
rect 36084 20383 36136 20392
rect 36084 20349 36093 20383
rect 36093 20349 36127 20383
rect 36127 20349 36136 20383
rect 36084 20340 36136 20349
rect 37096 20340 37148 20392
rect 35992 20272 36044 20324
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 28356 20000 28408 20052
rect 940 19864 992 19916
rect 3056 19864 3108 19916
rect 2596 19839 2648 19848
rect 2596 19805 2605 19839
rect 2605 19805 2639 19839
rect 2639 19805 2648 19839
rect 2596 19796 2648 19805
rect 24400 19839 24452 19848
rect 24400 19805 24409 19839
rect 24409 19805 24443 19839
rect 24443 19805 24452 19839
rect 24400 19796 24452 19805
rect 34612 19796 34664 19848
rect 35716 20000 35768 20052
rect 35992 19864 36044 19916
rect 36084 19864 36136 19916
rect 37280 19864 37332 19916
rect 24676 19771 24728 19780
rect 24676 19737 24710 19771
rect 24710 19737 24728 19771
rect 24676 19728 24728 19737
rect 3240 19660 3292 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 3148 19456 3200 19508
rect 3424 19456 3476 19508
rect 1860 19388 1912 19440
rect 17316 19456 17368 19508
rect 20260 19456 20312 19508
rect 2964 19320 3016 19372
rect 1952 19295 2004 19304
rect 1952 19261 1961 19295
rect 1961 19261 1995 19295
rect 1995 19261 2004 19295
rect 1952 19252 2004 19261
rect 3148 19252 3200 19304
rect 4068 19320 4120 19372
rect 21640 19363 21692 19372
rect 21640 19329 21649 19363
rect 21649 19329 21683 19363
rect 21683 19329 21692 19363
rect 21640 19320 21692 19329
rect 36084 19320 36136 19372
rect 22468 19252 22520 19304
rect 34796 19252 34848 19304
rect 36912 19295 36964 19304
rect 36912 19261 36921 19295
rect 36921 19261 36955 19295
rect 36955 19261 36964 19295
rect 36912 19252 36964 19261
rect 3516 19227 3568 19236
rect 3516 19193 3525 19227
rect 3525 19193 3559 19227
rect 3559 19193 3568 19227
rect 3516 19184 3568 19193
rect 2320 19116 2372 19168
rect 3424 19159 3476 19168
rect 3424 19125 3433 19159
rect 3433 19125 3467 19159
rect 3467 19125 3476 19159
rect 3424 19116 3476 19125
rect 26976 19159 27028 19168
rect 26976 19125 26985 19159
rect 26985 19125 27019 19159
rect 27019 19125 27028 19159
rect 26976 19116 27028 19125
rect 35624 19159 35676 19168
rect 35624 19125 35633 19159
rect 35633 19125 35667 19159
rect 35667 19125 35676 19159
rect 35624 19116 35676 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1860 18955 1912 18964
rect 1860 18921 1869 18955
rect 1869 18921 1903 18955
rect 1903 18921 1912 18955
rect 1860 18912 1912 18921
rect 2320 18708 2372 18760
rect 37096 18887 37148 18896
rect 37096 18853 37105 18887
rect 37105 18853 37139 18887
rect 37139 18853 37148 18887
rect 37096 18844 37148 18853
rect 3608 18708 3660 18760
rect 4344 18751 4396 18760
rect 4344 18717 4353 18751
rect 4353 18717 4387 18751
rect 4387 18717 4396 18751
rect 4344 18708 4396 18717
rect 4620 18708 4672 18760
rect 35348 18708 35400 18760
rect 1952 18615 2004 18624
rect 1952 18581 1961 18615
rect 1961 18581 1995 18615
rect 1995 18581 2004 18615
rect 1952 18572 2004 18581
rect 3332 18572 3384 18624
rect 34704 18615 34756 18624
rect 34704 18581 34713 18615
rect 34713 18581 34747 18615
rect 34747 18581 34756 18615
rect 34704 18572 34756 18581
rect 37004 18640 37056 18692
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 1952 18368 2004 18420
rect 4344 18368 4396 18420
rect 22468 18411 22520 18420
rect 22468 18377 22477 18411
rect 22477 18377 22511 18411
rect 22511 18377 22520 18411
rect 22468 18368 22520 18377
rect 24124 18411 24176 18420
rect 24124 18377 24133 18411
rect 24133 18377 24167 18411
rect 24167 18377 24176 18411
rect 24124 18368 24176 18377
rect 34704 18368 34756 18420
rect 34796 18368 34848 18420
rect 35992 18368 36044 18420
rect 37004 18368 37056 18420
rect 3424 18300 3476 18352
rect 34612 18300 34664 18352
rect 2320 18232 2372 18284
rect 2964 18232 3016 18284
rect 3792 18139 3844 18148
rect 3792 18105 3801 18139
rect 3801 18105 3835 18139
rect 3835 18105 3844 18139
rect 3792 18096 3844 18105
rect 2964 18028 3016 18080
rect 21824 18207 21876 18216
rect 21824 18173 21833 18207
rect 21833 18173 21867 18207
rect 21867 18173 21876 18207
rect 21824 18164 21876 18173
rect 26976 18232 27028 18284
rect 36084 18300 36136 18352
rect 35624 18232 35676 18284
rect 34796 18164 34848 18216
rect 23480 18096 23532 18148
rect 4712 18028 4764 18080
rect 35532 18028 35584 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 27528 17867 27580 17876
rect 27528 17833 27537 17867
rect 27537 17833 27571 17867
rect 27571 17833 27580 17867
rect 27528 17824 27580 17833
rect 1584 17731 1636 17740
rect 1584 17697 1593 17731
rect 1593 17697 1627 17731
rect 1627 17697 1636 17731
rect 1584 17688 1636 17697
rect 2964 17688 3016 17740
rect 2596 17663 2648 17672
rect 2596 17629 2605 17663
rect 2605 17629 2639 17663
rect 2639 17629 2648 17663
rect 2596 17620 2648 17629
rect 3332 17620 3384 17672
rect 27896 17756 27948 17808
rect 11888 17620 11940 17672
rect 3884 17484 3936 17536
rect 7564 17527 7616 17536
rect 7564 17493 7573 17527
rect 7573 17493 7607 17527
rect 7607 17493 7616 17527
rect 7564 17484 7616 17493
rect 21916 17484 21968 17536
rect 35256 17663 35308 17672
rect 35256 17629 35265 17663
rect 35265 17629 35299 17663
rect 35299 17629 35308 17663
rect 35256 17620 35308 17629
rect 35348 17620 35400 17672
rect 35532 17620 35584 17672
rect 30196 17484 30248 17536
rect 34520 17527 34572 17536
rect 34520 17493 34529 17527
rect 34529 17493 34563 17527
rect 34563 17493 34572 17527
rect 34520 17484 34572 17493
rect 34704 17527 34756 17536
rect 34704 17493 34713 17527
rect 34713 17493 34747 17527
rect 34747 17493 34756 17527
rect 34704 17484 34756 17493
rect 36820 17527 36872 17536
rect 36820 17493 36829 17527
rect 36829 17493 36863 17527
rect 36863 17493 36872 17527
rect 36820 17484 36872 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 2596 17280 2648 17332
rect 7564 17280 7616 17332
rect 34520 17280 34572 17332
rect 35256 17280 35308 17332
rect 36820 17280 36872 17332
rect 3700 17144 3752 17196
rect 4620 17144 4672 17196
rect 4896 17119 4948 17128
rect 4896 17085 4905 17119
rect 4905 17085 4939 17119
rect 4939 17085 4948 17119
rect 4896 17076 4948 17085
rect 36268 17119 36320 17128
rect 36268 17085 36277 17119
rect 36277 17085 36311 17119
rect 36311 17085 36320 17119
rect 36268 17076 36320 17085
rect 2872 16983 2924 16992
rect 2872 16949 2881 16983
rect 2881 16949 2915 16983
rect 2915 16949 2924 16983
rect 2872 16940 2924 16949
rect 4620 16940 4672 16992
rect 20904 16983 20956 16992
rect 20904 16949 20913 16983
rect 20913 16949 20947 16983
rect 20947 16949 20956 16983
rect 20904 16940 20956 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 2872 16736 2924 16788
rect 23480 16736 23532 16788
rect 34612 16736 34664 16788
rect 20904 16668 20956 16720
rect 21456 16668 21508 16720
rect 21916 16711 21968 16720
rect 21916 16677 21925 16711
rect 21925 16677 21959 16711
rect 21959 16677 21968 16711
rect 21916 16668 21968 16677
rect 3516 16600 3568 16652
rect 14280 16600 14332 16652
rect 34704 16668 34756 16720
rect 37188 16643 37240 16652
rect 37188 16609 37197 16643
rect 37197 16609 37231 16643
rect 37231 16609 37240 16643
rect 37188 16600 37240 16609
rect 1584 16575 1636 16584
rect 1584 16541 1593 16575
rect 1593 16541 1627 16575
rect 1627 16541 1636 16575
rect 1584 16532 1636 16541
rect 2596 16575 2648 16584
rect 2596 16541 2605 16575
rect 2605 16541 2639 16575
rect 2639 16541 2648 16575
rect 2596 16532 2648 16541
rect 3884 16532 3936 16584
rect 4252 16464 4304 16516
rect 13268 16464 13320 16516
rect 2872 16439 2924 16448
rect 2872 16405 2881 16439
rect 2881 16405 2915 16439
rect 2915 16405 2924 16439
rect 2872 16396 2924 16405
rect 3240 16396 3292 16448
rect 6552 16396 6604 16448
rect 20444 16396 20496 16448
rect 20720 16396 20772 16448
rect 24676 16532 24728 16584
rect 35992 16575 36044 16584
rect 35992 16541 36001 16575
rect 36001 16541 36035 16575
rect 36035 16541 36044 16575
rect 35992 16532 36044 16541
rect 36268 16575 36320 16584
rect 36268 16541 36277 16575
rect 36277 16541 36311 16575
rect 36311 16541 36320 16575
rect 36268 16532 36320 16541
rect 22284 16439 22336 16448
rect 22284 16405 22293 16439
rect 22293 16405 22327 16439
rect 22327 16405 22336 16439
rect 22284 16396 22336 16405
rect 24400 16396 24452 16448
rect 35440 16396 35492 16448
rect 35532 16396 35584 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 2596 16192 2648 16244
rect 2872 16192 2924 16244
rect 4252 16235 4304 16244
rect 4252 16201 4261 16235
rect 4261 16201 4295 16235
rect 4295 16201 4304 16235
rect 4252 16192 4304 16201
rect 13268 16235 13320 16244
rect 13268 16201 13277 16235
rect 13277 16201 13311 16235
rect 13311 16201 13320 16235
rect 13268 16192 13320 16201
rect 4068 16124 4120 16176
rect 4712 16124 4764 16176
rect 12808 16167 12860 16176
rect 12808 16133 12817 16167
rect 12817 16133 12851 16167
rect 12851 16133 12860 16167
rect 16120 16192 16172 16244
rect 17868 16192 17920 16244
rect 20720 16192 20772 16244
rect 21824 16192 21876 16244
rect 22284 16192 22336 16244
rect 35440 16192 35492 16244
rect 35992 16192 36044 16244
rect 12808 16124 12860 16133
rect 4620 16056 4672 16108
rect 20444 16099 20496 16108
rect 20444 16065 20478 16099
rect 20478 16065 20496 16099
rect 20444 16056 20496 16065
rect 21916 16056 21968 16108
rect 35532 16124 35584 16176
rect 35348 16056 35400 16108
rect 4896 15920 4948 15972
rect 13084 15963 13136 15972
rect 13084 15929 13093 15963
rect 13093 15929 13127 15963
rect 13127 15929 13136 15963
rect 13084 15920 13136 15929
rect 25320 15920 25372 15972
rect 23204 15895 23256 15904
rect 23204 15861 23213 15895
rect 23213 15861 23247 15895
rect 23247 15861 23256 15895
rect 23204 15852 23256 15861
rect 24400 15852 24452 15904
rect 34704 15895 34756 15904
rect 34704 15861 34713 15895
rect 34713 15861 34747 15895
rect 34747 15861 34756 15895
rect 34704 15852 34756 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 3240 15648 3292 15700
rect 3700 15648 3752 15700
rect 2872 15580 2924 15632
rect 11888 15623 11940 15632
rect 11888 15589 11897 15623
rect 11897 15589 11931 15623
rect 11931 15589 11940 15623
rect 11888 15580 11940 15589
rect 2596 15376 2648 15428
rect 2688 15308 2740 15360
rect 4068 15351 4120 15360
rect 4068 15317 4077 15351
rect 4077 15317 4111 15351
rect 4111 15317 4120 15351
rect 4068 15308 4120 15317
rect 12808 15648 12860 15700
rect 21916 15691 21968 15700
rect 21916 15657 21925 15691
rect 21925 15657 21959 15691
rect 21959 15657 21968 15691
rect 21916 15648 21968 15657
rect 24860 15580 24912 15632
rect 21456 15555 21508 15564
rect 21456 15521 21465 15555
rect 21465 15521 21499 15555
rect 21499 15521 21508 15555
rect 21456 15512 21508 15521
rect 34704 15512 34756 15564
rect 22008 15487 22060 15496
rect 22008 15453 22017 15487
rect 22017 15453 22051 15487
rect 22051 15453 22060 15487
rect 22008 15444 22060 15453
rect 22928 15444 22980 15496
rect 36544 15419 36596 15428
rect 36544 15385 36553 15419
rect 36553 15385 36587 15419
rect 36587 15385 36596 15419
rect 36544 15376 36596 15385
rect 13820 15308 13872 15360
rect 23388 15308 23440 15360
rect 34520 15308 34572 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 21456 15104 21508 15156
rect 1584 15079 1636 15088
rect 1584 15045 1593 15079
rect 1593 15045 1627 15079
rect 1627 15045 1636 15079
rect 1584 15036 1636 15045
rect 36912 15079 36964 15088
rect 36912 15045 36921 15079
rect 36921 15045 36955 15079
rect 36955 15045 36964 15079
rect 36912 15036 36964 15045
rect 2596 15011 2648 15020
rect 2596 14977 2605 15011
rect 2605 14977 2639 15011
rect 2639 14977 2648 15011
rect 2596 14968 2648 14977
rect 36544 14968 36596 15020
rect 1952 14900 2004 14952
rect 3976 14900 4028 14952
rect 3884 14832 3936 14884
rect 34428 14943 34480 14952
rect 34428 14909 34437 14943
rect 34437 14909 34471 14943
rect 34471 14909 34480 14943
rect 34428 14900 34480 14909
rect 35440 14900 35492 14952
rect 34704 14875 34756 14884
rect 34704 14841 34713 14875
rect 34713 14841 34747 14875
rect 34747 14841 34756 14875
rect 34704 14832 34756 14841
rect 3608 14807 3660 14816
rect 3608 14773 3617 14807
rect 3617 14773 3651 14807
rect 3651 14773 3660 14807
rect 3608 14764 3660 14773
rect 4068 14764 4120 14816
rect 35532 14764 35584 14816
rect 35716 14764 35768 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 1952 14603 2004 14612
rect 1952 14569 1961 14603
rect 1961 14569 1995 14603
rect 1995 14569 2004 14603
rect 1952 14560 2004 14569
rect 3608 14560 3660 14612
rect 3976 14560 4028 14612
rect 35440 14560 35492 14612
rect 3516 14424 3568 14476
rect 35348 14424 35400 14476
rect 34796 14399 34848 14408
rect 34796 14365 34805 14399
rect 34805 14365 34839 14399
rect 34839 14365 34848 14399
rect 34796 14356 34848 14365
rect 35532 14356 35584 14408
rect 3792 14263 3844 14272
rect 3792 14229 3801 14263
rect 3801 14229 3835 14263
rect 3835 14229 3844 14263
rect 3792 14220 3844 14229
rect 35808 14220 35860 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 34796 14016 34848 14068
rect 35808 14016 35860 14068
rect 25320 13923 25372 13932
rect 25320 13889 25329 13923
rect 25329 13889 25363 13923
rect 25363 13889 25372 13923
rect 25320 13880 25372 13889
rect 35716 13880 35768 13932
rect 2596 13812 2648 13864
rect 4068 13855 4120 13864
rect 4068 13821 4077 13855
rect 4077 13821 4111 13855
rect 4111 13821 4120 13855
rect 4068 13812 4120 13821
rect 29460 13812 29512 13864
rect 36268 13855 36320 13864
rect 36268 13821 36277 13855
rect 36277 13821 36311 13855
rect 36311 13821 36320 13855
rect 36268 13812 36320 13821
rect 3792 13787 3844 13796
rect 3792 13753 3801 13787
rect 3801 13753 3835 13787
rect 3835 13753 3844 13787
rect 3792 13744 3844 13753
rect 2964 13676 3016 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 2872 13515 2924 13524
rect 2872 13481 2881 13515
rect 2881 13481 2915 13515
rect 2915 13481 2924 13515
rect 2872 13472 2924 13481
rect 35440 13404 35492 13456
rect 940 13336 992 13388
rect 3424 13379 3476 13388
rect 3424 13345 3433 13379
rect 3433 13345 3467 13379
rect 3467 13345 3476 13379
rect 3424 13336 3476 13345
rect 6552 13379 6604 13388
rect 6552 13345 6561 13379
rect 6561 13345 6595 13379
rect 6595 13345 6604 13379
rect 6552 13336 6604 13345
rect 23204 13379 23256 13388
rect 23204 13345 23213 13379
rect 23213 13345 23247 13379
rect 23247 13345 23256 13379
rect 23204 13336 23256 13345
rect 37280 13336 37332 13388
rect 2596 13311 2648 13320
rect 2596 13277 2605 13311
rect 2605 13277 2639 13311
rect 2639 13277 2648 13311
rect 2596 13268 2648 13277
rect 3792 13311 3844 13320
rect 3792 13277 3801 13311
rect 3801 13277 3835 13311
rect 3835 13277 3844 13311
rect 3792 13268 3844 13277
rect 11060 13311 11112 13320
rect 11060 13277 11069 13311
rect 11069 13277 11103 13311
rect 11103 13277 11112 13311
rect 11060 13268 11112 13277
rect 13084 13268 13136 13320
rect 24860 13268 24912 13320
rect 28908 13268 28960 13320
rect 35992 13311 36044 13320
rect 35992 13277 36001 13311
rect 36001 13277 36035 13311
rect 36035 13277 36044 13311
rect 35992 13268 36044 13277
rect 36268 13311 36320 13320
rect 36268 13277 36277 13311
rect 36277 13277 36311 13311
rect 36311 13277 36320 13311
rect 36268 13268 36320 13277
rect 4436 13175 4488 13184
rect 4436 13141 4445 13175
rect 4445 13141 4479 13175
rect 4479 13141 4488 13175
rect 4436 13132 4488 13141
rect 7196 13175 7248 13184
rect 7196 13141 7205 13175
rect 7205 13141 7239 13175
rect 7239 13141 7248 13175
rect 7196 13132 7248 13141
rect 10416 13175 10468 13184
rect 10416 13141 10425 13175
rect 10425 13141 10459 13175
rect 10459 13141 10468 13175
rect 10416 13132 10468 13141
rect 23756 13175 23808 13184
rect 23756 13141 23765 13175
rect 23765 13141 23799 13175
rect 23799 13141 23808 13175
rect 23756 13132 23808 13141
rect 25964 13175 26016 13184
rect 25964 13141 25973 13175
rect 25973 13141 26007 13175
rect 26007 13141 26016 13175
rect 25964 13132 26016 13141
rect 34520 13175 34572 13184
rect 34520 13141 34529 13175
rect 34529 13141 34563 13175
rect 34563 13141 34572 13175
rect 34520 13132 34572 13141
rect 35532 13200 35584 13252
rect 35440 13132 35492 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 3792 12928 3844 12980
rect 4436 12928 4488 12980
rect 35440 12928 35492 12980
rect 35532 12928 35584 12980
rect 35992 12928 36044 12980
rect 1952 12835 2004 12844
rect 1952 12801 1961 12835
rect 1961 12801 1995 12835
rect 1995 12801 2004 12835
rect 1952 12792 2004 12801
rect 2964 12792 3016 12844
rect 3516 12792 3568 12844
rect 13820 12860 13872 12912
rect 14280 12792 14332 12844
rect 35348 12792 35400 12844
rect 3424 12631 3476 12640
rect 3424 12597 3433 12631
rect 3433 12597 3467 12631
rect 3467 12597 3476 12631
rect 3424 12588 3476 12597
rect 17224 12588 17276 12640
rect 34704 12631 34756 12640
rect 34704 12597 34713 12631
rect 34713 12597 34747 12631
rect 34747 12597 34756 12631
rect 34704 12588 34756 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 3424 12291 3476 12300
rect 3424 12257 3433 12291
rect 3433 12257 3467 12291
rect 3467 12257 3476 12291
rect 3424 12248 3476 12257
rect 34704 12248 34756 12300
rect 36544 12155 36596 12164
rect 36544 12121 36553 12155
rect 36553 12121 36587 12155
rect 36587 12121 36596 12155
rect 36544 12112 36596 12121
rect 2596 12044 2648 12096
rect 34520 12044 34572 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 36544 11840 36596 11892
rect 940 11772 992 11824
rect 2596 11747 2648 11756
rect 2596 11713 2605 11747
rect 2605 11713 2639 11747
rect 2639 11713 2648 11747
rect 2596 11704 2648 11713
rect 3700 11704 3752 11756
rect 37464 11772 37516 11824
rect 34520 11636 34572 11688
rect 35440 11636 35492 11688
rect 34704 11611 34756 11620
rect 34704 11577 34713 11611
rect 34713 11577 34747 11611
rect 34747 11577 34756 11611
rect 34704 11568 34756 11577
rect 2872 11543 2924 11552
rect 2872 11509 2881 11543
rect 2881 11509 2915 11543
rect 2915 11509 2924 11543
rect 2872 11500 2924 11509
rect 3424 11500 3476 11552
rect 3608 11543 3660 11552
rect 3608 11509 3617 11543
rect 3617 11509 3651 11543
rect 3651 11509 3660 11543
rect 3608 11500 3660 11509
rect 4068 11500 4120 11552
rect 35532 11500 35584 11552
rect 35624 11543 35676 11552
rect 35624 11509 35633 11543
rect 35633 11509 35667 11543
rect 35667 11509 35676 11543
rect 35624 11500 35676 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 1952 11203 2004 11212
rect 1952 11169 1961 11203
rect 1961 11169 1995 11203
rect 1995 11169 2004 11203
rect 1952 11160 2004 11169
rect 3608 11296 3660 11348
rect 35440 11296 35492 11348
rect 35348 11160 35400 11212
rect 34796 11135 34848 11144
rect 34796 11101 34805 11135
rect 34805 11101 34839 11135
rect 34839 11101 34848 11135
rect 34796 11092 34848 11101
rect 35532 11092 35584 11144
rect 3516 10956 3568 11008
rect 36820 10999 36872 11008
rect 36820 10965 36829 10999
rect 36829 10965 36863 10999
rect 36863 10965 36872 10999
rect 36820 10956 36872 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 28908 10795 28960 10804
rect 28908 10761 28917 10795
rect 28917 10761 28951 10795
rect 28951 10761 28960 10795
rect 28908 10752 28960 10761
rect 34796 10752 34848 10804
rect 17224 10659 17276 10668
rect 17224 10625 17233 10659
rect 17233 10625 17267 10659
rect 17267 10625 17276 10659
rect 17224 10616 17276 10625
rect 27896 10659 27948 10668
rect 27896 10625 27905 10659
rect 27905 10625 27939 10659
rect 27939 10625 27948 10659
rect 27896 10616 27948 10625
rect 28540 10616 28592 10668
rect 29460 10659 29512 10668
rect 29460 10625 29469 10659
rect 29469 10625 29503 10659
rect 29503 10625 29512 10659
rect 29460 10616 29512 10625
rect 35624 10616 35676 10668
rect 36820 10616 36872 10668
rect 36084 10591 36136 10600
rect 36084 10557 36093 10591
rect 36093 10557 36127 10591
rect 36127 10557 36136 10591
rect 36084 10548 36136 10557
rect 2596 10412 2648 10464
rect 2872 10412 2924 10464
rect 3608 10455 3660 10464
rect 3608 10421 3617 10455
rect 3617 10421 3651 10455
rect 3651 10421 3660 10455
rect 3608 10412 3660 10421
rect 4068 10412 4120 10464
rect 19340 10412 19392 10464
rect 27344 10455 27396 10464
rect 27344 10421 27353 10455
rect 27353 10421 27387 10455
rect 27387 10421 27396 10455
rect 27344 10412 27396 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 2872 10251 2924 10260
rect 2872 10217 2881 10251
rect 2881 10217 2915 10251
rect 2915 10217 2924 10251
rect 2872 10208 2924 10217
rect 11060 10208 11112 10260
rect 22928 10251 22980 10260
rect 22928 10217 22937 10251
rect 22937 10217 22971 10251
rect 22971 10217 22980 10251
rect 22928 10208 22980 10217
rect 35440 10140 35492 10192
rect 940 10072 992 10124
rect 7196 10072 7248 10124
rect 23756 10072 23808 10124
rect 35532 10072 35584 10124
rect 36084 10072 36136 10124
rect 37280 10072 37332 10124
rect 2596 10047 2648 10056
rect 2596 10013 2605 10047
rect 2605 10013 2639 10047
rect 2639 10013 2648 10047
rect 2596 10004 2648 10013
rect 3516 10047 3568 10056
rect 3516 10013 3525 10047
rect 3525 10013 3559 10047
rect 3559 10013 3568 10047
rect 3516 10004 3568 10013
rect 3792 10047 3844 10056
rect 3792 10013 3801 10047
rect 3801 10013 3835 10047
rect 3835 10013 3844 10047
rect 3792 10004 3844 10013
rect 16856 10004 16908 10056
rect 20904 10004 20956 10056
rect 35348 10004 35400 10056
rect 35992 10047 36044 10056
rect 35992 10013 36001 10047
rect 36001 10013 36035 10047
rect 36035 10013 36044 10047
rect 35992 10004 36044 10013
rect 4436 9911 4488 9920
rect 4436 9877 4445 9911
rect 4445 9877 4479 9911
rect 4479 9877 4488 9911
rect 4436 9868 4488 9877
rect 17132 9911 17184 9920
rect 17132 9877 17141 9911
rect 17141 9877 17175 9911
rect 17175 9877 17184 9911
rect 17132 9868 17184 9877
rect 31024 9911 31076 9920
rect 31024 9877 31033 9911
rect 31033 9877 31067 9911
rect 31067 9877 31076 9911
rect 34520 9979 34572 9988
rect 34520 9945 34529 9979
rect 34529 9945 34563 9979
rect 34563 9945 34572 9979
rect 34520 9936 34572 9945
rect 35808 9936 35860 9988
rect 31024 9868 31076 9877
rect 35440 9868 35492 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 3792 9664 3844 9716
rect 8668 9664 8720 9716
rect 17132 9664 17184 9716
rect 3608 9596 3660 9648
rect 1952 9571 2004 9580
rect 1952 9537 1961 9571
rect 1961 9537 1995 9571
rect 1995 9537 2004 9571
rect 1952 9528 2004 9537
rect 4436 9528 4488 9580
rect 35440 9664 35492 9716
rect 35992 9664 36044 9716
rect 35532 9596 35584 9648
rect 35348 9528 35400 9580
rect 3424 9367 3476 9376
rect 3424 9333 3433 9367
rect 3433 9333 3467 9367
rect 3467 9333 3476 9367
rect 3424 9324 3476 9333
rect 34704 9367 34756 9376
rect 34704 9333 34713 9367
rect 34713 9333 34747 9367
rect 34747 9333 34756 9367
rect 34704 9324 34756 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 3424 9120 3476 9172
rect 34704 9120 34756 9172
rect 36544 8891 36596 8900
rect 36544 8857 36553 8891
rect 36553 8857 36587 8891
rect 36587 8857 36596 8891
rect 36544 8848 36596 8857
rect 2596 8780 2648 8832
rect 34520 8780 34572 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 3424 8576 3476 8628
rect 34704 8576 34756 8628
rect 36544 8576 36596 8628
rect 940 8508 992 8560
rect 2596 8483 2648 8492
rect 2596 8449 2605 8483
rect 2605 8449 2639 8483
rect 2639 8449 2648 8483
rect 2596 8440 2648 8449
rect 34520 8372 34572 8424
rect 4068 8304 4120 8356
rect 37464 8508 37516 8560
rect 35440 8372 35492 8424
rect 2780 8236 2832 8288
rect 5448 8236 5500 8288
rect 35532 8236 35584 8288
rect 35624 8279 35676 8288
rect 35624 8245 35633 8279
rect 35633 8245 35667 8279
rect 35667 8245 35676 8279
rect 35624 8236 35676 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 12072 8032 12124 8084
rect 14280 8032 14332 8084
rect 35440 8032 35492 8084
rect 1952 7939 2004 7948
rect 1952 7905 1961 7939
rect 1961 7905 1995 7939
rect 1995 7905 2004 7939
rect 1952 7896 2004 7905
rect 19340 7896 19392 7948
rect 35348 7896 35400 7948
rect 2780 7828 2832 7880
rect 34704 7828 34756 7880
rect 34796 7871 34848 7880
rect 34796 7837 34805 7871
rect 34805 7837 34839 7871
rect 34839 7837 34848 7871
rect 34796 7828 34848 7837
rect 35532 7828 35584 7880
rect 10416 7803 10468 7812
rect 10416 7769 10425 7803
rect 10425 7769 10459 7803
rect 10459 7769 10468 7803
rect 10416 7760 10468 7769
rect 20260 7760 20312 7812
rect 20628 7760 20680 7812
rect 37280 7803 37332 7812
rect 37280 7769 37289 7803
rect 37289 7769 37323 7803
rect 37323 7769 37332 7803
rect 37280 7760 37332 7769
rect 4436 7735 4488 7744
rect 4436 7701 4445 7735
rect 4445 7701 4479 7735
rect 4479 7701 4488 7735
rect 4436 7692 4488 7701
rect 19248 7735 19300 7744
rect 19248 7701 19257 7735
rect 19257 7701 19291 7735
rect 19291 7701 19300 7735
rect 19248 7692 19300 7701
rect 33692 7692 33744 7744
rect 36820 7735 36872 7744
rect 36820 7701 36829 7735
rect 36829 7701 36863 7735
rect 36863 7701 36872 7735
rect 36820 7692 36872 7701
rect 36912 7692 36964 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 4712 7420 4764 7472
rect 10416 7488 10468 7540
rect 20628 7488 20680 7540
rect 34796 7488 34848 7540
rect 31024 7420 31076 7472
rect 1952 7352 2004 7404
rect 3332 7395 3384 7404
rect 3332 7361 3341 7395
rect 3341 7361 3375 7395
rect 3375 7361 3384 7395
rect 36820 7488 36872 7540
rect 3332 7352 3384 7361
rect 35624 7352 35676 7404
rect 4988 7327 5040 7336
rect 4988 7293 4997 7327
rect 4997 7293 5031 7327
rect 5031 7293 5040 7327
rect 4988 7284 5040 7293
rect 5448 7284 5500 7336
rect 33508 7327 33560 7336
rect 33508 7293 33517 7327
rect 33517 7293 33551 7327
rect 33551 7293 33560 7327
rect 33508 7284 33560 7293
rect 34336 7284 34388 7336
rect 36176 7327 36228 7336
rect 36176 7293 36185 7327
rect 36185 7293 36219 7327
rect 36219 7293 36228 7327
rect 36176 7284 36228 7293
rect 4804 7216 4856 7268
rect 3424 7148 3476 7200
rect 3700 7191 3752 7200
rect 3700 7157 3709 7191
rect 3709 7157 3743 7191
rect 3743 7157 3752 7191
rect 3700 7148 3752 7157
rect 3792 7148 3844 7200
rect 5172 7191 5224 7200
rect 5172 7157 5181 7191
rect 5181 7157 5215 7191
rect 5215 7157 5224 7191
rect 5172 7148 5224 7157
rect 24400 7148 24452 7200
rect 29552 7148 29604 7200
rect 33968 7148 34020 7200
rect 34244 7191 34296 7200
rect 34244 7157 34253 7191
rect 34253 7157 34287 7191
rect 34287 7157 34296 7191
rect 34244 7148 34296 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 3332 6851 3384 6860
rect 3332 6817 3341 6851
rect 3341 6817 3375 6851
rect 3375 6817 3384 6851
rect 3332 6808 3384 6817
rect 4804 6944 4856 6996
rect 4988 6876 5040 6928
rect 35440 6876 35492 6928
rect 4620 6808 4672 6860
rect 33692 6808 33744 6860
rect 34244 6808 34296 6860
rect 37188 6851 37240 6860
rect 37188 6817 37197 6851
rect 37197 6817 37231 6851
rect 37231 6817 37240 6851
rect 37188 6808 37240 6817
rect 5172 6740 5224 6792
rect 35992 6783 36044 6792
rect 35992 6749 36001 6783
rect 36001 6749 36035 6783
rect 36035 6749 36044 6783
rect 35992 6740 36044 6749
rect 36176 6783 36228 6792
rect 36176 6749 36185 6783
rect 36185 6749 36219 6783
rect 36219 6749 36228 6783
rect 36176 6740 36228 6749
rect 2780 6604 2832 6656
rect 4712 6672 4764 6724
rect 5448 6604 5500 6656
rect 32404 6647 32456 6656
rect 32404 6613 32413 6647
rect 32413 6613 32447 6647
rect 32447 6613 32456 6647
rect 32404 6604 32456 6613
rect 33048 6604 33100 6656
rect 34152 6604 34204 6656
rect 34520 6604 34572 6656
rect 35256 6647 35308 6656
rect 35256 6613 35265 6647
rect 35265 6613 35299 6647
rect 35299 6613 35308 6647
rect 35256 6604 35308 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 4988 6400 5040 6452
rect 33508 6400 33560 6452
rect 35256 6400 35308 6452
rect 35992 6400 36044 6452
rect 1584 6375 1636 6384
rect 1584 6341 1593 6375
rect 1593 6341 1627 6375
rect 1627 6341 1636 6375
rect 1584 6332 1636 6341
rect 2596 6307 2648 6316
rect 2596 6273 2605 6307
rect 2605 6273 2639 6307
rect 2639 6273 2648 6307
rect 2596 6264 2648 6273
rect 3424 6307 3476 6316
rect 3424 6273 3433 6307
rect 3433 6273 3467 6307
rect 3467 6273 3476 6307
rect 3424 6264 3476 6273
rect 34060 6264 34112 6316
rect 3608 6239 3660 6248
rect 3608 6205 3617 6239
rect 3617 6205 3651 6239
rect 3651 6205 3660 6239
rect 3608 6196 3660 6205
rect 18512 6239 18564 6248
rect 18512 6205 18521 6239
rect 18521 6205 18555 6239
rect 18555 6205 18564 6239
rect 18512 6196 18564 6205
rect 19248 6196 19300 6248
rect 34152 6196 34204 6248
rect 34520 6239 34572 6248
rect 34520 6205 34529 6239
rect 34529 6205 34563 6239
rect 34563 6205 34572 6239
rect 34520 6196 34572 6205
rect 34704 6239 34756 6248
rect 34704 6205 34713 6239
rect 34713 6205 34747 6239
rect 34747 6205 34756 6239
rect 34704 6196 34756 6205
rect 35256 6307 35308 6316
rect 35256 6273 35265 6307
rect 35265 6273 35299 6307
rect 35299 6273 35308 6307
rect 35256 6264 35308 6273
rect 35348 6264 35400 6316
rect 2872 6103 2924 6112
rect 2872 6069 2881 6103
rect 2881 6069 2915 6103
rect 2915 6069 2924 6103
rect 2872 6060 2924 6069
rect 14004 6103 14056 6112
rect 14004 6069 14013 6103
rect 14013 6069 14047 6103
rect 14047 6069 14056 6103
rect 14004 6060 14056 6069
rect 20720 6060 20772 6112
rect 33876 6103 33928 6112
rect 33876 6069 33885 6103
rect 33885 6069 33919 6103
rect 33919 6069 33928 6103
rect 33876 6060 33928 6069
rect 36176 6060 36228 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 2596 5856 2648 5908
rect 3608 5856 3660 5908
rect 30196 5899 30248 5908
rect 30196 5865 30205 5899
rect 30205 5865 30239 5899
rect 30239 5865 30248 5899
rect 30196 5856 30248 5865
rect 33876 5856 33928 5908
rect 13544 5831 13596 5840
rect 13544 5797 13553 5831
rect 13553 5797 13587 5831
rect 13587 5797 13596 5831
rect 13544 5788 13596 5797
rect 14464 5831 14516 5840
rect 14464 5797 14473 5831
rect 14473 5797 14507 5831
rect 14507 5797 14516 5831
rect 14464 5788 14516 5797
rect 16488 5788 16540 5840
rect 34152 5788 34204 5840
rect 2780 5720 2832 5772
rect 3700 5652 3752 5704
rect 10876 5652 10928 5704
rect 10968 5695 11020 5704
rect 10968 5661 10977 5695
rect 10977 5661 11011 5695
rect 11011 5661 11020 5695
rect 10968 5652 11020 5661
rect 11888 5720 11940 5772
rect 32404 5720 32456 5772
rect 9312 5584 9364 5636
rect 12164 5652 12216 5704
rect 13084 5695 13136 5704
rect 13084 5661 13093 5695
rect 13093 5661 13127 5695
rect 13127 5661 13136 5695
rect 13084 5652 13136 5661
rect 14004 5584 14056 5636
rect 15752 5584 15804 5636
rect 31392 5584 31444 5636
rect 33876 5652 33928 5704
rect 33968 5652 34020 5704
rect 34244 5720 34296 5772
rect 34612 5652 34664 5704
rect 35716 5652 35768 5704
rect 34428 5584 34480 5636
rect 9956 5516 10008 5568
rect 10876 5516 10928 5568
rect 11244 5516 11296 5568
rect 11980 5516 12032 5568
rect 14372 5516 14424 5568
rect 15200 5559 15252 5568
rect 15200 5525 15209 5559
rect 15209 5525 15243 5559
rect 15243 5525 15252 5559
rect 15200 5516 15252 5525
rect 29092 5559 29144 5568
rect 29092 5525 29101 5559
rect 29101 5525 29135 5559
rect 29135 5525 29144 5559
rect 29092 5516 29144 5525
rect 29552 5516 29604 5568
rect 32220 5516 32272 5568
rect 35624 5584 35676 5636
rect 35900 5627 35952 5636
rect 35900 5593 35909 5627
rect 35909 5593 35943 5627
rect 35943 5593 35952 5627
rect 35900 5584 35952 5593
rect 36544 5627 36596 5636
rect 36544 5593 36553 5627
rect 36553 5593 36587 5627
rect 36587 5593 36596 5627
rect 36544 5584 36596 5593
rect 34888 5516 34940 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 3516 5355 3568 5364
rect 3516 5321 3525 5355
rect 3525 5321 3559 5355
rect 3559 5321 3568 5355
rect 3516 5312 3568 5321
rect 3792 5244 3844 5296
rect 2872 5219 2924 5228
rect 2872 5185 2881 5219
rect 2881 5185 2915 5219
rect 2915 5185 2924 5219
rect 2872 5176 2924 5185
rect 9956 5108 10008 5160
rect 11244 5151 11296 5160
rect 11244 5117 11253 5151
rect 11253 5117 11287 5151
rect 11287 5117 11296 5151
rect 11244 5108 11296 5117
rect 13084 5312 13136 5364
rect 14464 5312 14516 5364
rect 14924 5355 14976 5364
rect 14924 5321 14933 5355
rect 14933 5321 14967 5355
rect 14967 5321 14976 5355
rect 14924 5312 14976 5321
rect 15752 5312 15804 5364
rect 16120 5287 16172 5296
rect 16120 5253 16129 5287
rect 16129 5253 16163 5287
rect 16163 5253 16172 5287
rect 16120 5244 16172 5253
rect 13084 5151 13136 5160
rect 13084 5117 13093 5151
rect 13093 5117 13127 5151
rect 13127 5117 13136 5151
rect 13084 5108 13136 5117
rect 13728 5151 13780 5160
rect 13728 5117 13737 5151
rect 13737 5117 13771 5151
rect 13771 5117 13780 5151
rect 13728 5108 13780 5117
rect 14464 5151 14516 5160
rect 14464 5117 14473 5151
rect 14473 5117 14507 5151
rect 14507 5117 14516 5151
rect 14464 5108 14516 5117
rect 15476 5151 15528 5160
rect 15476 5117 15485 5151
rect 15485 5117 15519 5151
rect 15519 5117 15528 5151
rect 15476 5108 15528 5117
rect 25964 5176 26016 5228
rect 31392 5219 31444 5228
rect 31392 5185 31401 5219
rect 31401 5185 31435 5219
rect 31435 5185 31444 5219
rect 31392 5176 31444 5185
rect 34244 5244 34296 5296
rect 35900 5312 35952 5364
rect 34520 5244 34572 5296
rect 34612 5244 34664 5296
rect 12256 5040 12308 5092
rect 18512 5040 18564 5092
rect 2596 4972 2648 5024
rect 9772 4972 9824 5024
rect 9956 5015 10008 5024
rect 9956 4981 9965 5015
rect 9965 4981 9999 5015
rect 9999 4981 10008 5015
rect 9956 4972 10008 4981
rect 10600 5015 10652 5024
rect 10600 4981 10609 5015
rect 10609 4981 10643 5015
rect 10643 4981 10652 5015
rect 10600 4972 10652 4981
rect 10692 5015 10744 5024
rect 10692 4981 10701 5015
rect 10701 4981 10735 5015
rect 10735 4981 10744 5015
rect 10692 4972 10744 4981
rect 12624 4972 12676 5024
rect 17684 4972 17736 5024
rect 27160 5151 27212 5160
rect 27160 5117 27169 5151
rect 27169 5117 27203 5151
rect 27203 5117 27212 5151
rect 27160 5108 27212 5117
rect 28172 5151 28224 5160
rect 28172 5117 28181 5151
rect 28181 5117 28215 5151
rect 28215 5117 28224 5151
rect 28172 5108 28224 5117
rect 29460 5151 29512 5160
rect 29460 5117 29469 5151
rect 29469 5117 29503 5151
rect 29503 5117 29512 5151
rect 29460 5108 29512 5117
rect 29552 5108 29604 5160
rect 30196 5108 30248 5160
rect 30656 5108 30708 5160
rect 29368 5040 29420 5092
rect 31852 5040 31904 5092
rect 32772 5151 32824 5160
rect 32772 5117 32781 5151
rect 32781 5117 32815 5151
rect 32815 5117 32824 5151
rect 32772 5108 32824 5117
rect 34796 5108 34848 5160
rect 32404 5040 32456 5092
rect 19340 4972 19392 5024
rect 26240 4972 26292 5024
rect 27804 5015 27856 5024
rect 27804 4981 27813 5015
rect 27813 4981 27847 5015
rect 27847 4981 27856 5015
rect 27804 4972 27856 4981
rect 30288 5015 30340 5024
rect 30288 4981 30297 5015
rect 30297 4981 30331 5015
rect 30331 4981 30340 5015
rect 30288 4972 30340 4981
rect 31760 4972 31812 5024
rect 31944 5015 31996 5024
rect 31944 4981 31953 5015
rect 31953 4981 31987 5015
rect 31987 4981 31996 5015
rect 31944 4972 31996 4981
rect 32220 4972 32272 5024
rect 32680 5015 32732 5024
rect 32680 4981 32689 5015
rect 32689 4981 32723 5015
rect 32723 4981 32732 5015
rect 32680 4972 32732 4981
rect 36084 5151 36136 5160
rect 36084 5117 36093 5151
rect 36093 5117 36127 5151
rect 36127 5117 36136 5151
rect 36084 5108 36136 5117
rect 37096 4972 37148 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 10968 4768 11020 4820
rect 13084 4768 13136 4820
rect 29460 4768 29512 4820
rect 33876 4768 33928 4820
rect 36084 4768 36136 4820
rect 9772 4743 9824 4752
rect 9772 4709 9781 4743
rect 9781 4709 9815 4743
rect 9815 4709 9824 4743
rect 9772 4700 9824 4709
rect 940 4632 992 4684
rect 19248 4700 19300 4752
rect 26148 4743 26200 4752
rect 26148 4709 26157 4743
rect 26157 4709 26191 4743
rect 26191 4709 26200 4743
rect 26148 4700 26200 4709
rect 31392 4700 31444 4752
rect 12072 4675 12124 4684
rect 12072 4641 12081 4675
rect 12081 4641 12115 4675
rect 12115 4641 12124 4675
rect 12072 4632 12124 4641
rect 13544 4632 13596 4684
rect 14924 4632 14976 4684
rect 16672 4675 16724 4684
rect 16672 4641 16681 4675
rect 16681 4641 16715 4675
rect 16715 4641 16724 4675
rect 16672 4632 16724 4641
rect 2596 4607 2648 4616
rect 2596 4573 2605 4607
rect 2605 4573 2639 4607
rect 2639 4573 2648 4607
rect 2596 4564 2648 4573
rect 10600 4564 10652 4616
rect 12440 4564 12492 4616
rect 13176 4607 13228 4616
rect 13176 4573 13185 4607
rect 13185 4573 13219 4607
rect 13219 4573 13228 4607
rect 13176 4564 13228 4573
rect 13820 4607 13872 4616
rect 13820 4573 13829 4607
rect 13829 4573 13863 4607
rect 13863 4573 13872 4607
rect 13820 4564 13872 4573
rect 16488 4607 16540 4616
rect 16488 4573 16497 4607
rect 16497 4573 16531 4607
rect 16531 4573 16540 4607
rect 16488 4564 16540 4573
rect 18236 4607 18288 4616
rect 18236 4573 18245 4607
rect 18245 4573 18279 4607
rect 18279 4573 18288 4607
rect 18236 4564 18288 4573
rect 5448 4496 5500 4548
rect 9956 4496 10008 4548
rect 27712 4632 27764 4684
rect 29460 4632 29512 4684
rect 30196 4632 30248 4684
rect 31116 4675 31168 4684
rect 31116 4641 31125 4675
rect 31125 4641 31159 4675
rect 31159 4641 31168 4675
rect 31116 4632 31168 4641
rect 26332 4607 26384 4616
rect 26332 4573 26341 4607
rect 26341 4573 26375 4607
rect 26375 4573 26384 4607
rect 26332 4564 26384 4573
rect 28632 4607 28684 4616
rect 28632 4573 28641 4607
rect 28641 4573 28675 4607
rect 28675 4573 28684 4607
rect 28632 4564 28684 4573
rect 28724 4564 28776 4616
rect 33876 4632 33928 4684
rect 34060 4675 34112 4684
rect 34060 4641 34069 4675
rect 34069 4641 34103 4675
rect 34103 4641 34112 4675
rect 34060 4632 34112 4641
rect 33508 4564 33560 4616
rect 34796 4564 34848 4616
rect 35808 4632 35860 4684
rect 37648 4632 37700 4684
rect 11060 4428 11112 4480
rect 12532 4471 12584 4480
rect 12532 4437 12541 4471
rect 12541 4437 12575 4471
rect 12575 4437 12584 4471
rect 12532 4428 12584 4437
rect 14096 4471 14148 4480
rect 14096 4437 14105 4471
rect 14105 4437 14139 4471
rect 14139 4437 14148 4471
rect 14096 4428 14148 4437
rect 15660 4471 15712 4480
rect 15660 4437 15669 4471
rect 15669 4437 15703 4471
rect 15703 4437 15712 4471
rect 15660 4428 15712 4437
rect 15844 4471 15896 4480
rect 15844 4437 15853 4471
rect 15853 4437 15887 4471
rect 15887 4437 15896 4471
rect 15844 4428 15896 4437
rect 17224 4471 17276 4480
rect 17224 4437 17233 4471
rect 17233 4437 17267 4471
rect 17267 4437 17276 4471
rect 17224 4428 17276 4437
rect 17316 4428 17368 4480
rect 18788 4428 18840 4480
rect 19340 4428 19392 4480
rect 33692 4496 33744 4548
rect 36544 4564 36596 4616
rect 37096 4564 37148 4616
rect 26240 4428 26292 4480
rect 26700 4428 26752 4480
rect 27068 4471 27120 4480
rect 27068 4437 27077 4471
rect 27077 4437 27111 4471
rect 27111 4437 27120 4471
rect 27068 4428 27120 4437
rect 28448 4471 28500 4480
rect 28448 4437 28457 4471
rect 28457 4437 28491 4471
rect 28491 4437 28500 4471
rect 28448 4428 28500 4437
rect 30104 4471 30156 4480
rect 30104 4437 30113 4471
rect 30113 4437 30147 4471
rect 30147 4437 30156 4471
rect 30104 4428 30156 4437
rect 34520 4428 34572 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 12072 4224 12124 4276
rect 13176 4224 13228 4276
rect 26976 4224 27028 4276
rect 28632 4224 28684 4276
rect 31116 4224 31168 4276
rect 37004 4224 37056 4276
rect 2964 4088 3016 4140
rect 9312 4131 9364 4140
rect 9312 4097 9321 4131
rect 9321 4097 9355 4131
rect 9355 4097 9364 4131
rect 9312 4088 9364 4097
rect 10140 4131 10192 4140
rect 10140 4097 10149 4131
rect 10149 4097 10183 4131
rect 10183 4097 10192 4131
rect 10140 4088 10192 4097
rect 11888 4088 11940 4140
rect 14372 4131 14424 4140
rect 14372 4097 14390 4131
rect 14390 4097 14424 4131
rect 26240 4156 26292 4208
rect 14648 4131 14700 4140
rect 14372 4088 14424 4097
rect 14648 4097 14657 4131
rect 14657 4097 14691 4131
rect 14691 4097 14700 4131
rect 14648 4088 14700 4097
rect 15292 4131 15344 4140
rect 15292 4097 15301 4131
rect 15301 4097 15335 4131
rect 15335 4097 15344 4131
rect 15292 4088 15344 4097
rect 10600 4063 10652 4072
rect 10600 4029 10609 4063
rect 10609 4029 10643 4063
rect 10643 4029 10652 4063
rect 10600 4020 10652 4029
rect 13636 4020 13688 4072
rect 15016 4020 15068 4072
rect 16948 4063 17000 4072
rect 16948 4029 16957 4063
rect 16957 4029 16991 4063
rect 16991 4029 17000 4063
rect 16948 4020 17000 4029
rect 18052 4063 18104 4072
rect 18052 4029 18061 4063
rect 18061 4029 18095 4063
rect 18095 4029 18104 4063
rect 18052 4020 18104 4029
rect 19156 4063 19208 4072
rect 19156 4029 19165 4063
rect 19165 4029 19199 4063
rect 19199 4029 19208 4063
rect 19156 4020 19208 4029
rect 25320 4020 25372 4072
rect 2596 3884 2648 3936
rect 32772 4156 32824 4208
rect 26976 4131 27028 4140
rect 26976 4097 26985 4131
rect 26985 4097 27019 4131
rect 27019 4097 27028 4131
rect 26976 4088 27028 4097
rect 28724 4088 28776 4140
rect 30472 4131 30524 4140
rect 30472 4097 30481 4131
rect 30481 4097 30515 4131
rect 30515 4097 30524 4131
rect 30472 4088 30524 4097
rect 32496 4088 32548 4140
rect 34152 4156 34204 4208
rect 34796 4156 34848 4208
rect 34244 4088 34296 4140
rect 34520 4088 34572 4140
rect 35440 4088 35492 4140
rect 35900 4131 35952 4140
rect 35900 4097 35909 4131
rect 35909 4097 35943 4131
rect 35943 4097 35952 4131
rect 35900 4088 35952 4097
rect 36636 4131 36688 4140
rect 36636 4097 36645 4131
rect 36645 4097 36679 4131
rect 36679 4097 36688 4131
rect 36636 4088 36688 4097
rect 27528 4063 27580 4072
rect 27528 4029 27537 4063
rect 27537 4029 27571 4063
rect 27571 4029 27580 4063
rect 27528 4020 27580 4029
rect 28632 4020 28684 4072
rect 29736 4020 29788 4072
rect 32128 4063 32180 4072
rect 32128 4029 32137 4063
rect 32137 4029 32171 4063
rect 32171 4029 32180 4063
rect 32128 4020 32180 4029
rect 14464 3884 14516 3936
rect 19984 3884 20036 3936
rect 24860 3927 24912 3936
rect 24860 3893 24869 3927
rect 24869 3893 24903 3927
rect 24903 3893 24912 3927
rect 24860 3884 24912 3893
rect 26884 3884 26936 3936
rect 30656 3952 30708 4004
rect 33140 3884 33192 3936
rect 34428 3884 34480 3936
rect 34612 3884 34664 3936
rect 36912 3884 36964 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 12164 3723 12216 3732
rect 12164 3689 12173 3723
rect 12173 3689 12207 3723
rect 12207 3689 12216 3723
rect 12164 3680 12216 3689
rect 13820 3680 13872 3732
rect 14648 3680 14700 3732
rect 940 3544 992 3596
rect 2596 3519 2648 3528
rect 2596 3485 2605 3519
rect 2605 3485 2639 3519
rect 2639 3485 2648 3519
rect 2596 3476 2648 3485
rect 10324 3612 10376 3664
rect 10140 3587 10192 3596
rect 10140 3553 10149 3587
rect 10149 3553 10183 3587
rect 10183 3553 10192 3587
rect 10140 3544 10192 3553
rect 12072 3544 12124 3596
rect 16672 3680 16724 3732
rect 18236 3680 18288 3732
rect 26332 3680 26384 3732
rect 26976 3680 27028 3732
rect 29552 3680 29604 3732
rect 32128 3680 32180 3732
rect 29460 3612 29512 3664
rect 8668 3519 8720 3528
rect 8668 3485 8677 3519
rect 8677 3485 8711 3519
rect 8711 3485 8720 3519
rect 8668 3476 8720 3485
rect 10692 3476 10744 3528
rect 15200 3476 15252 3528
rect 19248 3587 19300 3596
rect 19248 3553 19257 3587
rect 19257 3553 19291 3587
rect 19291 3553 19300 3587
rect 19248 3544 19300 3553
rect 17408 3519 17460 3528
rect 17408 3485 17417 3519
rect 17417 3485 17451 3519
rect 17451 3485 17460 3519
rect 17408 3476 17460 3485
rect 6644 3451 6696 3460
rect 6644 3417 6653 3451
rect 6653 3417 6687 3451
rect 6687 3417 6696 3451
rect 6644 3408 6696 3417
rect 8300 3451 8352 3460
rect 8300 3417 8309 3451
rect 8309 3417 8343 3451
rect 8343 3417 8352 3451
rect 8300 3408 8352 3417
rect 11060 3451 11112 3460
rect 11060 3417 11094 3451
rect 11094 3417 11112 3451
rect 11060 3408 11112 3417
rect 12072 3408 12124 3460
rect 17960 3408 18012 3460
rect 18788 3408 18840 3460
rect 14556 3383 14608 3392
rect 14556 3349 14565 3383
rect 14565 3349 14599 3383
rect 14599 3349 14608 3383
rect 14556 3340 14608 3349
rect 19432 3340 19484 3392
rect 24860 3408 24912 3460
rect 27528 3544 27580 3596
rect 32772 3680 32824 3732
rect 34336 3680 34388 3732
rect 34520 3680 34572 3732
rect 34612 3680 34664 3732
rect 26884 3519 26936 3528
rect 26884 3485 26893 3519
rect 26893 3485 26927 3519
rect 26927 3485 26936 3519
rect 26884 3476 26936 3485
rect 27068 3476 27120 3528
rect 29092 3476 29144 3528
rect 29552 3519 29604 3528
rect 29552 3485 29561 3519
rect 29561 3485 29595 3519
rect 29595 3485 29604 3519
rect 29552 3476 29604 3485
rect 34428 3587 34480 3596
rect 34428 3553 34437 3587
rect 34437 3553 34471 3587
rect 34471 3553 34480 3587
rect 34428 3544 34480 3553
rect 26792 3408 26844 3460
rect 30104 3408 30156 3460
rect 34152 3476 34204 3528
rect 35716 3612 35768 3664
rect 37096 3723 37148 3732
rect 37096 3689 37105 3723
rect 37105 3689 37139 3723
rect 37139 3689 37148 3723
rect 37096 3680 37148 3689
rect 36176 3476 36228 3528
rect 31392 3408 31444 3460
rect 32680 3408 32732 3460
rect 31024 3340 31076 3392
rect 33692 3340 33744 3392
rect 34520 3340 34572 3392
rect 34796 3340 34848 3392
rect 36268 3408 36320 3460
rect 36912 3408 36964 3460
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 8300 3136 8352 3188
rect 12072 3179 12124 3188
rect 12072 3145 12081 3179
rect 12081 3145 12115 3179
rect 12115 3145 12124 3179
rect 12072 3136 12124 3145
rect 2596 3043 2648 3052
rect 2596 3009 2605 3043
rect 2605 3009 2639 3043
rect 2639 3009 2648 3043
rect 2596 3000 2648 3009
rect 9956 3000 10008 3052
rect 11980 3000 12032 3052
rect 12256 3000 12308 3052
rect 14096 3000 14148 3052
rect 15844 3136 15896 3188
rect 17408 3136 17460 3188
rect 17960 3136 18012 3188
rect 19156 3136 19208 3188
rect 19432 3136 19484 3188
rect 26240 3136 26292 3188
rect 26792 3179 26844 3188
rect 26792 3145 26801 3179
rect 26801 3145 26835 3179
rect 26835 3145 26844 3179
rect 26792 3136 26844 3145
rect 27160 3136 27212 3188
rect 29552 3179 29604 3188
rect 29552 3145 29561 3179
rect 29561 3145 29595 3179
rect 29595 3145 29604 3179
rect 29552 3136 29604 3145
rect 30472 3136 30524 3188
rect 31024 3179 31076 3188
rect 31024 3145 31033 3179
rect 31033 3145 31067 3179
rect 31067 3145 31076 3179
rect 31024 3136 31076 3145
rect 34244 3136 34296 3188
rect 15292 3111 15344 3120
rect 15292 3077 15301 3111
rect 15301 3077 15335 3111
rect 15335 3077 15344 3111
rect 15292 3068 15344 3077
rect 15660 3000 15712 3052
rect 17316 3043 17368 3052
rect 17316 3009 17325 3043
rect 17325 3009 17359 3043
rect 17359 3009 17368 3043
rect 17316 3000 17368 3009
rect 17684 3111 17736 3120
rect 17684 3077 17718 3111
rect 17718 3077 17736 3111
rect 17684 3068 17736 3077
rect 20628 3111 20680 3120
rect 1584 2975 1636 2984
rect 1584 2941 1593 2975
rect 1593 2941 1627 2975
rect 1627 2941 1636 2975
rect 1584 2932 1636 2941
rect 7656 2975 7708 2984
rect 7656 2941 7665 2975
rect 7665 2941 7699 2975
rect 7699 2941 7708 2975
rect 7656 2932 7708 2941
rect 8760 2932 8812 2984
rect 11152 2932 11204 2984
rect 12900 2975 12952 2984
rect 12900 2941 12909 2975
rect 12909 2941 12943 2975
rect 12943 2941 12952 2975
rect 12900 2932 12952 2941
rect 15200 2932 15252 2984
rect 19340 2975 19392 2984
rect 19340 2941 19349 2975
rect 19349 2941 19383 2975
rect 19383 2941 19392 2975
rect 20628 3077 20637 3111
rect 20637 3077 20671 3111
rect 20671 3077 20680 3111
rect 20628 3068 20680 3077
rect 27712 3068 27764 3120
rect 22192 3000 22244 3052
rect 23388 3043 23440 3052
rect 23388 3009 23397 3043
rect 23397 3009 23431 3043
rect 23431 3009 23440 3043
rect 23388 3000 23440 3009
rect 27344 3000 27396 3052
rect 31392 3068 31444 3120
rect 31852 3111 31904 3120
rect 31852 3077 31861 3111
rect 31861 3077 31895 3111
rect 31895 3077 31904 3111
rect 31852 3068 31904 3077
rect 33508 3068 33560 3120
rect 28448 3000 28500 3052
rect 29368 3000 29420 3052
rect 19340 2932 19392 2941
rect 20076 2975 20128 2984
rect 20076 2941 20085 2975
rect 20085 2941 20119 2975
rect 20119 2941 20128 2975
rect 20076 2932 20128 2941
rect 20904 2932 20956 2984
rect 23940 2975 23992 2984
rect 23940 2941 23949 2975
rect 23949 2941 23983 2975
rect 23983 2941 23992 2975
rect 23940 2932 23992 2941
rect 13728 2864 13780 2916
rect 26976 2932 27028 2984
rect 29092 2975 29144 2984
rect 29092 2941 29101 2975
rect 29101 2941 29135 2975
rect 29135 2941 29144 2975
rect 29092 2932 29144 2941
rect 31944 3000 31996 3052
rect 33876 3000 33928 3052
rect 35348 3000 35400 3052
rect 35624 3000 35676 3052
rect 1768 2796 1820 2848
rect 16948 2796 17000 2848
rect 33048 2864 33100 2916
rect 28172 2796 28224 2848
rect 31208 2796 31260 2848
rect 34428 2932 34480 2984
rect 34244 2864 34296 2916
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 12440 2635 12492 2644
rect 12440 2601 12449 2635
rect 12449 2601 12483 2635
rect 12483 2601 12492 2635
rect 12440 2592 12492 2601
rect 15476 2592 15528 2644
rect 16488 2592 16540 2644
rect 19248 2635 19300 2644
rect 19248 2601 19257 2635
rect 19257 2601 19291 2635
rect 19291 2601 19300 2635
rect 19248 2592 19300 2601
rect 16856 2524 16908 2576
rect 2596 2456 2648 2508
rect 6092 2456 6144 2508
rect 9128 2456 9180 2508
rect 12072 2456 12124 2508
rect 12532 2456 12584 2508
rect 12624 2456 12676 2508
rect 14556 2456 14608 2508
rect 17224 2499 17276 2508
rect 17224 2465 17233 2499
rect 17233 2465 17267 2499
rect 17267 2465 17276 2499
rect 17224 2456 17276 2465
rect 18144 2499 18196 2508
rect 18144 2465 18153 2499
rect 18153 2465 18187 2499
rect 18187 2465 18196 2499
rect 18144 2456 18196 2465
rect 19984 2592 20036 2644
rect 26148 2635 26200 2644
rect 26148 2601 26157 2635
rect 26157 2601 26191 2635
rect 26191 2601 26200 2635
rect 26148 2592 26200 2601
rect 28540 2592 28592 2644
rect 28724 2592 28776 2644
rect 31852 2592 31904 2644
rect 33600 2635 33652 2644
rect 33600 2601 33609 2635
rect 33609 2601 33643 2635
rect 33643 2601 33652 2635
rect 33600 2592 33652 2601
rect 35900 2592 35952 2644
rect 37280 2635 37332 2644
rect 37280 2601 37289 2635
rect 37289 2601 37323 2635
rect 37323 2601 37332 2635
rect 37280 2592 37332 2601
rect 34428 2524 34480 2576
rect 34520 2524 34572 2576
rect 19984 2456 20036 2508
rect 22192 2499 22244 2508
rect 22192 2465 22201 2499
rect 22201 2465 22235 2499
rect 22235 2465 22244 2499
rect 22192 2456 22244 2465
rect 22836 2456 22888 2508
rect 2688 2431 2740 2440
rect 2688 2397 2697 2431
rect 2697 2397 2731 2431
rect 2731 2397 2740 2431
rect 2688 2388 2740 2397
rect 3332 2431 3384 2440
rect 3332 2397 3341 2431
rect 3341 2397 3375 2431
rect 3375 2397 3384 2431
rect 3332 2388 3384 2397
rect 4712 2431 4764 2440
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 4712 2388 4764 2397
rect 6644 2388 6696 2440
rect 8760 2431 8812 2440
rect 8760 2397 8769 2431
rect 8769 2397 8803 2431
rect 8803 2397 8812 2431
rect 8760 2388 8812 2397
rect 11152 2431 11204 2440
rect 11152 2397 11161 2431
rect 11161 2397 11195 2431
rect 11195 2397 11204 2431
rect 11152 2388 11204 2397
rect 12900 2388 12952 2440
rect 15200 2431 15252 2440
rect 15200 2397 15209 2431
rect 15209 2397 15243 2431
rect 15243 2397 15252 2431
rect 15200 2388 15252 2397
rect 18052 2388 18104 2440
rect 20076 2431 20128 2440
rect 20076 2397 20085 2431
rect 20085 2397 20119 2431
rect 20119 2397 20128 2431
rect 20076 2388 20128 2397
rect 20720 2388 20772 2440
rect 23940 2388 23992 2440
rect 13544 2363 13596 2372
rect 13544 2329 13553 2363
rect 13553 2329 13587 2363
rect 13587 2329 13596 2363
rect 13544 2320 13596 2329
rect 16304 2363 16356 2372
rect 16304 2329 16313 2363
rect 16313 2329 16347 2363
rect 16347 2329 16356 2363
rect 16304 2320 16356 2329
rect 24124 2320 24176 2372
rect 26700 2431 26752 2440
rect 26700 2397 26709 2431
rect 26709 2397 26743 2431
rect 26743 2397 26752 2431
rect 26700 2388 26752 2397
rect 26976 2431 27028 2440
rect 26976 2397 26985 2431
rect 26985 2397 27019 2431
rect 27019 2397 27028 2431
rect 26976 2388 27028 2397
rect 27160 2388 27212 2440
rect 30288 2456 30340 2508
rect 32496 2499 32548 2508
rect 32496 2465 32505 2499
rect 32505 2465 32539 2499
rect 32539 2465 32548 2499
rect 32496 2456 32548 2465
rect 33140 2456 33192 2508
rect 27804 2388 27856 2440
rect 29092 2388 29144 2440
rect 31760 2388 31812 2440
rect 33232 2388 33284 2440
rect 34704 2431 34756 2440
rect 34704 2397 34713 2431
rect 34713 2397 34747 2431
rect 34747 2397 34756 2431
rect 34704 2388 34756 2397
rect 37924 2320 37976 2372
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 21640 1300 21692 1352
rect 34520 1300 34572 1352
<< metal2 >>
rect 1122 38200 1178 39000
rect 2870 38200 2926 39000
rect 4618 38200 4674 39000
rect 6366 38200 6422 39000
rect 8114 38200 8170 39000
rect 9862 38200 9918 39000
rect 11610 38200 11666 39000
rect 13358 38200 13414 39000
rect 15106 38200 15162 39000
rect 16854 38200 16910 39000
rect 18602 38200 18658 39000
rect 20350 38298 20406 39000
rect 20350 38270 20668 38298
rect 20350 38200 20406 38270
rect 1136 34950 1164 38200
rect 2884 36242 2912 38200
rect 3330 36544 3386 36553
rect 3330 36479 3386 36488
rect 2872 36236 2924 36242
rect 2872 36178 2924 36184
rect 2780 36168 2832 36174
rect 2780 36110 2832 36116
rect 2136 36032 2188 36038
rect 2136 35974 2188 35980
rect 1952 35080 2004 35086
rect 1952 35022 2004 35028
rect 1124 34944 1176 34950
rect 1124 34886 1176 34892
rect 1964 34610 1992 35022
rect 2044 35012 2096 35018
rect 2044 34954 2096 34960
rect 2056 34746 2084 34954
rect 2044 34740 2096 34746
rect 2044 34682 2096 34688
rect 2148 34610 2176 35974
rect 2792 34746 2820 36110
rect 3148 35692 3200 35698
rect 3148 35634 3200 35640
rect 2964 35012 3016 35018
rect 2964 34954 3016 34960
rect 2780 34740 2832 34746
rect 2780 34682 2832 34688
rect 2688 34672 2740 34678
rect 2688 34614 2740 34620
rect 1952 34604 2004 34610
rect 1952 34546 2004 34552
rect 2136 34604 2188 34610
rect 2136 34546 2188 34552
rect 2596 34468 2648 34474
rect 2596 34410 2648 34416
rect 2608 34066 2636 34410
rect 2596 34060 2648 34066
rect 2596 34002 2648 34008
rect 2504 33516 2556 33522
rect 2504 33458 2556 33464
rect 1582 33280 1638 33289
rect 1582 33215 1638 33224
rect 1596 32978 1624 33215
rect 1584 32972 1636 32978
rect 1584 32914 1636 32920
rect 1584 32360 1636 32366
rect 1584 32302 1636 32308
rect 1596 31657 1624 32302
rect 1582 31648 1638 31657
rect 1582 31583 1638 31592
rect 1584 31272 1636 31278
rect 1584 31214 1636 31220
rect 1596 30297 1624 31214
rect 1582 30288 1638 30297
rect 1582 30223 1638 30232
rect 1584 29096 1636 29102
rect 1584 29038 1636 29044
rect 1596 28393 1624 29038
rect 1952 28552 2004 28558
rect 1952 28494 2004 28500
rect 1582 28384 1638 28393
rect 1582 28319 1638 28328
rect 1584 28008 1636 28014
rect 1584 27950 1636 27956
rect 1596 27033 1624 27950
rect 1582 27024 1638 27033
rect 1964 26994 1992 28494
rect 2516 27606 2544 33458
rect 2596 33448 2648 33454
rect 2596 33390 2648 33396
rect 2608 32910 2636 33390
rect 2596 32904 2648 32910
rect 2596 32846 2648 32852
rect 2596 32428 2648 32434
rect 2596 32370 2648 32376
rect 2608 32026 2636 32370
rect 2596 32020 2648 32026
rect 2596 31962 2648 31968
rect 2596 31340 2648 31346
rect 2596 31282 2648 31288
rect 2608 30938 2636 31282
rect 2596 30932 2648 30938
rect 2596 30874 2648 30880
rect 2700 30258 2728 34614
rect 2976 34542 3004 34954
rect 3056 34944 3108 34950
rect 3056 34886 3108 34892
rect 2964 34536 3016 34542
rect 2964 34478 3016 34484
rect 2872 33856 2924 33862
rect 2872 33798 2924 33804
rect 2884 33522 2912 33798
rect 2872 33516 2924 33522
rect 2872 33458 2924 33464
rect 3068 32502 3096 34886
rect 3056 32496 3108 32502
rect 3056 32438 3108 32444
rect 2780 31816 2832 31822
rect 2780 31758 2832 31764
rect 2964 31816 3016 31822
rect 2964 31758 3016 31764
rect 2792 31482 2820 31758
rect 2780 31476 2832 31482
rect 2780 31418 2832 31424
rect 2872 31272 2924 31278
rect 2872 31214 2924 31220
rect 2884 30938 2912 31214
rect 2872 30932 2924 30938
rect 2872 30874 2924 30880
rect 2688 30252 2740 30258
rect 2688 30194 2740 30200
rect 2700 29646 2728 30194
rect 2976 30054 3004 31758
rect 3056 30728 3108 30734
rect 3056 30670 3108 30676
rect 3068 30394 3096 30670
rect 3056 30388 3108 30394
rect 3056 30330 3108 30336
rect 2964 30048 3016 30054
rect 2964 29990 3016 29996
rect 2688 29640 2740 29646
rect 2688 29582 2740 29588
rect 2700 28558 2728 29582
rect 2780 29164 2832 29170
rect 2780 29106 2832 29112
rect 2688 28552 2740 28558
rect 2688 28494 2740 28500
rect 2792 28150 2820 29106
rect 2780 28144 2832 28150
rect 2780 28086 2832 28092
rect 2596 28076 2648 28082
rect 2596 28018 2648 28024
rect 2504 27600 2556 27606
rect 2504 27542 2556 27548
rect 2608 27538 2636 28018
rect 2596 27532 2648 27538
rect 2596 27474 2648 27480
rect 3160 27130 3188 35634
rect 3240 33992 3292 33998
rect 3240 33934 3292 33940
rect 3252 30938 3280 33934
rect 3344 33454 3372 36479
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 3608 36168 3660 36174
rect 3608 36110 3660 36116
rect 4528 36168 4580 36174
rect 4528 36110 4580 36116
rect 3620 35766 3648 36110
rect 3608 35760 3660 35766
rect 3608 35702 3660 35708
rect 3700 35692 3752 35698
rect 3700 35634 3752 35640
rect 3712 34202 3740 35634
rect 3792 35624 3844 35630
rect 3792 35566 3844 35572
rect 4540 35578 4568 36110
rect 4632 35766 4660 38200
rect 4712 36032 4764 36038
rect 4712 35974 4764 35980
rect 4620 35760 4672 35766
rect 4620 35702 4672 35708
rect 3700 34196 3752 34202
rect 3700 34138 3752 34144
rect 3804 33998 3832 35566
rect 4540 35550 4660 35578
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4632 35290 4660 35550
rect 4620 35284 4672 35290
rect 4620 35226 4672 35232
rect 4620 35148 4672 35154
rect 4620 35090 4672 35096
rect 3884 34944 3936 34950
rect 3884 34886 3936 34892
rect 4066 34912 4122 34921
rect 3896 34610 3924 34886
rect 4066 34847 4122 34856
rect 3884 34604 3936 34610
rect 3884 34546 3936 34552
rect 4080 34082 4108 34847
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4080 34054 4200 34082
rect 4172 34048 4200 34054
rect 4252 34060 4304 34066
rect 4172 34020 4252 34048
rect 4252 34002 4304 34008
rect 3792 33992 3844 33998
rect 3792 33934 3844 33940
rect 3332 33448 3384 33454
rect 3332 33390 3384 33396
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 3792 32904 3844 32910
rect 3792 32846 3844 32852
rect 3516 32768 3568 32774
rect 3516 32710 3568 32716
rect 3240 30932 3292 30938
rect 3240 30874 3292 30880
rect 3424 30728 3476 30734
rect 3424 30670 3476 30676
rect 3240 30252 3292 30258
rect 3240 30194 3292 30200
rect 3252 29306 3280 30194
rect 3436 29850 3464 30670
rect 3424 29844 3476 29850
rect 3424 29786 3476 29792
rect 3240 29300 3292 29306
rect 3240 29242 3292 29248
rect 3240 27396 3292 27402
rect 3240 27338 3292 27344
rect 3148 27124 3200 27130
rect 3148 27066 3200 27072
rect 1582 26959 1638 26968
rect 1952 26988 2004 26994
rect 1952 26930 2004 26936
rect 1964 26450 1992 26930
rect 1952 26444 2004 26450
rect 1952 26386 2004 26392
rect 940 25832 992 25838
rect 940 25774 992 25780
rect 952 25129 980 25774
rect 1964 25294 1992 26386
rect 3252 26382 3280 27338
rect 3528 26994 3556 32710
rect 3804 29850 3832 32846
rect 4528 32836 4580 32842
rect 4528 32778 4580 32784
rect 4540 32570 4568 32778
rect 4528 32564 4580 32570
rect 4528 32506 4580 32512
rect 4632 32434 4660 35090
rect 4724 33522 4752 35974
rect 5724 35692 5776 35698
rect 5724 35634 5776 35640
rect 4804 35216 4856 35222
rect 4804 35158 4856 35164
rect 4816 34066 4844 35158
rect 4896 35012 4948 35018
rect 4896 34954 4948 34960
rect 4804 34060 4856 34066
rect 4804 34002 4856 34008
rect 4908 33998 4936 34954
rect 5736 34746 5764 35634
rect 6380 35630 6408 38200
rect 8128 36242 8156 38200
rect 8116 36236 8168 36242
rect 8116 36178 8168 36184
rect 6552 36168 6604 36174
rect 6552 36110 6604 36116
rect 8760 36168 8812 36174
rect 8760 36110 8812 36116
rect 9772 36168 9824 36174
rect 9772 36110 9824 36116
rect 6368 35624 6420 35630
rect 6368 35566 6420 35572
rect 6368 35012 6420 35018
rect 6368 34954 6420 34960
rect 5908 34944 5960 34950
rect 5908 34886 5960 34892
rect 5920 34746 5948 34886
rect 5724 34740 5776 34746
rect 5724 34682 5776 34688
rect 5908 34740 5960 34746
rect 5908 34682 5960 34688
rect 6000 34604 6052 34610
rect 6000 34546 6052 34552
rect 6012 34202 6040 34546
rect 6000 34196 6052 34202
rect 6000 34138 6052 34144
rect 5264 34060 5316 34066
rect 5264 34002 5316 34008
rect 4896 33992 4948 33998
rect 4896 33934 4948 33940
rect 4712 33516 4764 33522
rect 4712 33458 4764 33464
rect 4712 33312 4764 33318
rect 4712 33254 4764 33260
rect 4620 32428 4672 32434
rect 4620 32370 4672 32376
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4436 31680 4488 31686
rect 4436 31622 4488 31628
rect 4448 31346 4476 31622
rect 4436 31340 4488 31346
rect 4436 31282 4488 31288
rect 4620 31340 4672 31346
rect 4620 31282 4672 31288
rect 4068 31136 4120 31142
rect 4068 31078 4120 31084
rect 4080 30190 4108 31078
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4632 30870 4660 31282
rect 4620 30864 4672 30870
rect 4620 30806 4672 30812
rect 4724 30734 4752 33254
rect 4908 30802 4936 33934
rect 5276 33658 5304 34002
rect 6380 33658 6408 34954
rect 6564 34202 6592 36110
rect 6736 36100 6788 36106
rect 6736 36042 6788 36048
rect 6748 35698 6776 36042
rect 8772 35766 8800 36110
rect 9220 36032 9272 36038
rect 9220 35974 9272 35980
rect 8760 35760 8812 35766
rect 8760 35702 8812 35708
rect 6736 35692 6788 35698
rect 6736 35634 6788 35640
rect 8852 35692 8904 35698
rect 8852 35634 8904 35640
rect 7656 35012 7708 35018
rect 7656 34954 7708 34960
rect 7380 34944 7432 34950
rect 7380 34886 7432 34892
rect 7392 34746 7420 34886
rect 7380 34740 7432 34746
rect 7380 34682 7432 34688
rect 7012 34400 7064 34406
rect 7012 34342 7064 34348
rect 6552 34196 6604 34202
rect 6552 34138 6604 34144
rect 5264 33652 5316 33658
rect 5264 33594 5316 33600
rect 6368 33652 6420 33658
rect 6368 33594 6420 33600
rect 6000 33448 6052 33454
rect 6000 33390 6052 33396
rect 6012 32570 6040 33390
rect 6564 33386 6592 34138
rect 7024 34066 7052 34342
rect 7668 34202 7696 34954
rect 8864 34746 8892 35634
rect 8944 35012 8996 35018
rect 8944 34954 8996 34960
rect 8956 34746 8984 34954
rect 8852 34740 8904 34746
rect 8852 34682 8904 34688
rect 8944 34740 8996 34746
rect 8944 34682 8996 34688
rect 8208 34536 8260 34542
rect 8208 34478 8260 34484
rect 8024 34400 8076 34406
rect 8024 34342 8076 34348
rect 7656 34196 7708 34202
rect 7656 34138 7708 34144
rect 8036 34066 8064 34342
rect 8220 34202 8248 34478
rect 9232 34474 9260 35974
rect 9784 35290 9812 36110
rect 9876 35630 9904 38200
rect 10140 35692 10192 35698
rect 10140 35634 10192 35640
rect 9864 35624 9916 35630
rect 9864 35566 9916 35572
rect 9772 35284 9824 35290
rect 9772 35226 9824 35232
rect 9588 35080 9640 35086
rect 9588 35022 9640 35028
rect 9600 34542 9628 35022
rect 10152 34610 10180 35634
rect 11624 35630 11652 38200
rect 13372 36242 13400 38200
rect 13360 36236 13412 36242
rect 13360 36178 13412 36184
rect 12164 36168 12216 36174
rect 12164 36110 12216 36116
rect 12440 36168 12492 36174
rect 12440 36110 12492 36116
rect 14188 36168 14240 36174
rect 14188 36110 14240 36116
rect 14464 36168 14516 36174
rect 14464 36110 14516 36116
rect 11980 36100 12032 36106
rect 11980 36042 12032 36048
rect 11796 36032 11848 36038
rect 11796 35974 11848 35980
rect 11612 35624 11664 35630
rect 11612 35566 11664 35572
rect 11808 35154 11836 35974
rect 11992 35698 12020 36042
rect 11980 35692 12032 35698
rect 11980 35634 12032 35640
rect 11796 35148 11848 35154
rect 11796 35090 11848 35096
rect 11244 35012 11296 35018
rect 11244 34954 11296 34960
rect 11256 34746 11284 34954
rect 11336 34944 11388 34950
rect 11336 34886 11388 34892
rect 12072 34944 12124 34950
rect 12072 34886 12124 34892
rect 11060 34740 11112 34746
rect 11060 34682 11112 34688
rect 11244 34740 11296 34746
rect 11244 34682 11296 34688
rect 10140 34604 10192 34610
rect 10140 34546 10192 34552
rect 10600 34604 10652 34610
rect 10600 34546 10652 34552
rect 9588 34536 9640 34542
rect 9588 34478 9640 34484
rect 9220 34468 9272 34474
rect 9220 34410 9272 34416
rect 8208 34196 8260 34202
rect 8208 34138 8260 34144
rect 9232 34066 9260 34410
rect 7012 34060 7064 34066
rect 7012 34002 7064 34008
rect 8024 34060 8076 34066
rect 8024 34002 8076 34008
rect 9220 34060 9272 34066
rect 9220 34002 9272 34008
rect 6828 33992 6880 33998
rect 6828 33934 6880 33940
rect 6840 33658 6868 33934
rect 6828 33652 6880 33658
rect 6828 33594 6880 33600
rect 6552 33380 6604 33386
rect 6552 33322 6604 33328
rect 6276 32904 6328 32910
rect 6276 32846 6328 32852
rect 6000 32564 6052 32570
rect 6000 32506 6052 32512
rect 4896 30796 4948 30802
rect 4896 30738 4948 30744
rect 4712 30728 4764 30734
rect 4712 30670 4764 30676
rect 4620 30592 4672 30598
rect 4620 30534 4672 30540
rect 4068 30184 4120 30190
rect 4068 30126 4120 30132
rect 3792 29844 3844 29850
rect 3792 29786 3844 29792
rect 3792 29640 3844 29646
rect 3792 29582 3844 29588
rect 3804 27130 3832 29582
rect 4080 29170 4108 30126
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4632 29646 4660 30534
rect 4620 29640 4672 29646
rect 4620 29582 4672 29588
rect 4068 29164 4120 29170
rect 4068 29106 4120 29112
rect 4160 29096 4212 29102
rect 4080 29044 4160 29050
rect 4080 29038 4212 29044
rect 4080 29022 4200 29038
rect 4620 29028 4672 29034
rect 3884 28960 3936 28966
rect 3884 28902 3936 28908
rect 3896 28558 3924 28902
rect 4080 28762 4108 29022
rect 4620 28970 4672 28976
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4068 28756 4120 28762
rect 4068 28698 4120 28704
rect 3884 28552 3936 28558
rect 3884 28494 3936 28500
rect 3896 27606 3924 28494
rect 4436 28416 4488 28422
rect 4436 28358 4488 28364
rect 4448 28218 4476 28358
rect 4436 28212 4488 28218
rect 4436 28154 4488 28160
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 3884 27600 3936 27606
rect 3884 27542 3936 27548
rect 4632 27470 4660 28970
rect 4344 27464 4396 27470
rect 4344 27406 4396 27412
rect 4620 27464 4672 27470
rect 4620 27406 4672 27412
rect 4356 27130 4384 27406
rect 4632 27130 4660 27406
rect 3792 27124 3844 27130
rect 3792 27066 3844 27072
rect 4344 27124 4396 27130
rect 4344 27066 4396 27072
rect 4620 27124 4672 27130
rect 4620 27066 4672 27072
rect 3332 26988 3384 26994
rect 3332 26930 3384 26936
rect 3516 26988 3568 26994
rect 3516 26930 3568 26936
rect 3976 26988 4028 26994
rect 3976 26930 4028 26936
rect 3344 26586 3372 26930
rect 3332 26580 3384 26586
rect 3332 26522 3384 26528
rect 3240 26376 3292 26382
rect 3240 26318 3292 26324
rect 2780 25900 2832 25906
rect 2780 25842 2832 25848
rect 1952 25288 2004 25294
rect 1952 25230 2004 25236
rect 938 25120 994 25129
rect 938 25055 994 25064
rect 940 24744 992 24750
rect 940 24686 992 24692
rect 952 23497 980 24686
rect 1964 23662 1992 25230
rect 2792 24886 2820 25842
rect 3700 25832 3752 25838
rect 3700 25774 3752 25780
rect 3712 25498 3740 25774
rect 3792 25696 3844 25702
rect 3792 25638 3844 25644
rect 3700 25492 3752 25498
rect 3700 25434 3752 25440
rect 3804 25294 3832 25638
rect 3792 25288 3844 25294
rect 3792 25230 3844 25236
rect 2780 24880 2832 24886
rect 2780 24822 2832 24828
rect 2596 24812 2648 24818
rect 2596 24754 2648 24760
rect 1952 23656 2004 23662
rect 1952 23598 2004 23604
rect 938 23488 994 23497
rect 938 23423 994 23432
rect 2608 23186 2636 24754
rect 3240 24608 3292 24614
rect 3240 24550 3292 24556
rect 2780 24200 2832 24206
rect 2780 24142 2832 24148
rect 2688 23520 2740 23526
rect 2792 23474 2820 24142
rect 2964 24064 3016 24070
rect 2964 24006 3016 24012
rect 2740 23468 2820 23474
rect 2688 23462 2820 23468
rect 2700 23446 2820 23462
rect 2596 23180 2648 23186
rect 2596 23122 2648 23128
rect 2596 22636 2648 22642
rect 2596 22578 2648 22584
rect 1584 22568 1636 22574
rect 1584 22510 1636 22516
rect 1596 22001 1624 22510
rect 1582 21992 1638 22001
rect 1582 21927 1638 21936
rect 2608 21622 2636 22578
rect 2792 22030 2820 23446
rect 2976 22658 3004 24006
rect 3252 23866 3280 24550
rect 3792 24200 3844 24206
rect 3792 24142 3844 24148
rect 3804 23866 3832 24142
rect 3240 23860 3292 23866
rect 3240 23802 3292 23808
rect 3792 23860 3844 23866
rect 3792 23802 3844 23808
rect 3424 23656 3476 23662
rect 3424 23598 3476 23604
rect 2976 22630 3096 22658
rect 2964 22568 3016 22574
rect 2964 22510 3016 22516
rect 2872 22432 2924 22438
rect 2872 22374 2924 22380
rect 2780 22024 2832 22030
rect 2780 21966 2832 21972
rect 2596 21616 2648 21622
rect 2596 21558 2648 21564
rect 2596 20868 2648 20874
rect 2596 20810 2648 20816
rect 1952 20392 2004 20398
rect 1952 20334 2004 20340
rect 938 20224 994 20233
rect 938 20159 994 20168
rect 952 19922 980 20159
rect 940 19916 992 19922
rect 940 19858 992 19864
rect 1860 19440 1912 19446
rect 1860 19382 1912 19388
rect 1872 18970 1900 19382
rect 1964 19310 1992 20334
rect 2608 19854 2636 20810
rect 2792 20534 2820 21966
rect 2884 21554 2912 22374
rect 2976 21962 3004 22510
rect 2964 21956 3016 21962
rect 2964 21898 3016 21904
rect 2872 21548 2924 21554
rect 2872 21490 2924 21496
rect 2872 20936 2924 20942
rect 2872 20878 2924 20884
rect 2884 20602 2912 20878
rect 2872 20596 2924 20602
rect 2872 20538 2924 20544
rect 2780 20528 2832 20534
rect 2780 20470 2832 20476
rect 3068 19922 3096 22630
rect 3056 19916 3108 19922
rect 3056 19858 3108 19864
rect 2596 19848 2648 19854
rect 2596 19790 2648 19796
rect 3240 19712 3292 19718
rect 3240 19654 3292 19660
rect 3148 19508 3200 19514
rect 3148 19450 3200 19456
rect 2964 19372 3016 19378
rect 2964 19314 3016 19320
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 2320 19168 2372 19174
rect 2320 19110 2372 19116
rect 1860 18964 1912 18970
rect 1860 18906 1912 18912
rect 2332 18766 2360 19110
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 1952 18624 2004 18630
rect 1582 18592 1638 18601
rect 1952 18566 2004 18572
rect 1582 18527 1638 18536
rect 1596 17746 1624 18527
rect 1964 18426 1992 18566
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 2332 18290 2360 18702
rect 2976 18290 3004 19314
rect 3160 19310 3188 19450
rect 3148 19304 3200 19310
rect 3148 19246 3200 19252
rect 2320 18284 2372 18290
rect 2320 18226 2372 18232
rect 2964 18284 3016 18290
rect 2964 18226 3016 18232
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 2976 17746 3004 18022
rect 1584 17740 1636 17746
rect 1584 17682 1636 17688
rect 2964 17740 3016 17746
rect 2964 17682 3016 17688
rect 2596 17672 2648 17678
rect 2596 17614 2648 17620
rect 2608 17338 2636 17614
rect 2596 17332 2648 17338
rect 2596 17274 2648 17280
rect 2872 16992 2924 16998
rect 2872 16934 2924 16940
rect 2884 16794 2912 16934
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 1582 16688 1638 16697
rect 1582 16623 1638 16632
rect 1596 16590 1624 16623
rect 1584 16584 1636 16590
rect 1584 16526 1636 16532
rect 2596 16584 2648 16590
rect 3252 16574 3280 19654
rect 3436 19514 3464 23598
rect 3608 22432 3660 22438
rect 3608 22374 3660 22380
rect 3620 22030 3648 22374
rect 3608 22024 3660 22030
rect 3608 21966 3660 21972
rect 3792 21888 3844 21894
rect 3792 21830 3844 21836
rect 3804 21690 3832 21830
rect 3792 21684 3844 21690
rect 3792 21626 3844 21632
rect 3988 21418 4016 26930
rect 4068 26920 4120 26926
rect 4068 26862 4120 26868
rect 4080 23866 4108 26862
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4724 26234 4752 30670
rect 4908 29238 4936 30738
rect 6288 29850 6316 32846
rect 8116 31816 8168 31822
rect 8116 31758 8168 31764
rect 6276 29844 6328 29850
rect 6276 29786 6328 29792
rect 8128 29714 8156 31758
rect 6920 29708 6972 29714
rect 6920 29650 6972 29656
rect 8116 29708 8168 29714
rect 8116 29650 8168 29656
rect 4896 29232 4948 29238
rect 4948 29180 5028 29186
rect 4896 29174 5028 29180
rect 4908 29158 5028 29174
rect 4896 28960 4948 28966
rect 4896 28902 4948 28908
rect 4908 28558 4936 28902
rect 4896 28552 4948 28558
rect 4896 28494 4948 28500
rect 5000 27538 5028 29158
rect 4988 27532 5040 27538
rect 4988 27474 5040 27480
rect 5000 27146 5028 27474
rect 4816 27118 5028 27146
rect 4816 26382 4844 27118
rect 4988 27056 5040 27062
rect 4988 26998 5040 27004
rect 4896 26920 4948 26926
rect 4896 26862 4948 26868
rect 4908 26586 4936 26862
rect 4896 26580 4948 26586
rect 4896 26522 4948 26528
rect 4804 26376 4856 26382
rect 4804 26318 4856 26324
rect 4632 26206 4752 26234
rect 4632 25770 4660 26206
rect 4816 25838 4844 26318
rect 4804 25832 4856 25838
rect 4804 25774 4856 25780
rect 4620 25764 4672 25770
rect 4620 25706 4672 25712
rect 4712 25696 4764 25702
rect 4712 25638 4764 25644
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4160 25288 4212 25294
rect 4160 25230 4212 25236
rect 4172 24682 4200 25230
rect 4436 25152 4488 25158
rect 4436 25094 4488 25100
rect 4448 24818 4476 25094
rect 4436 24812 4488 24818
rect 4436 24754 4488 24760
rect 4620 24744 4672 24750
rect 4620 24686 4672 24692
rect 4160 24676 4212 24682
rect 4160 24618 4212 24624
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4436 24064 4488 24070
rect 4436 24006 4488 24012
rect 4448 23866 4476 24006
rect 4068 23860 4120 23866
rect 4068 23802 4120 23808
rect 4436 23860 4488 23866
rect 4436 23802 4488 23808
rect 4068 23520 4120 23526
rect 4068 23462 4120 23468
rect 4080 23322 4108 23462
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4068 23316 4120 23322
rect 4068 23258 4120 23264
rect 4080 23202 4108 23258
rect 4080 23174 4200 23202
rect 4068 22568 4120 22574
rect 4068 22510 4120 22516
rect 4080 21486 4108 22510
rect 4172 22506 4200 23174
rect 4632 22574 4660 24686
rect 4724 24206 4752 25638
rect 4816 24750 4844 25774
rect 5000 25770 5028 26998
rect 6932 26382 6960 29650
rect 9600 27062 9628 34478
rect 10612 34202 10640 34546
rect 11072 34474 11100 34682
rect 11348 34678 11376 34886
rect 11336 34672 11388 34678
rect 11336 34614 11388 34620
rect 12084 34610 12112 34886
rect 12176 34746 12204 36110
rect 12452 35290 12480 36110
rect 14200 35766 14228 36110
rect 14188 35760 14240 35766
rect 14188 35702 14240 35708
rect 14476 35290 14504 36110
rect 15016 36032 15068 36038
rect 15016 35974 15068 35980
rect 15028 35894 15056 35974
rect 14936 35866 15056 35894
rect 14648 35692 14700 35698
rect 14648 35634 14700 35640
rect 12440 35284 12492 35290
rect 12440 35226 12492 35232
rect 14464 35284 14516 35290
rect 14464 35226 14516 35232
rect 14188 35148 14240 35154
rect 14188 35090 14240 35096
rect 13176 35012 13228 35018
rect 13176 34954 13228 34960
rect 12164 34740 12216 34746
rect 12164 34682 12216 34688
rect 12072 34604 12124 34610
rect 12072 34546 12124 34552
rect 11060 34468 11112 34474
rect 11060 34410 11112 34416
rect 12072 34400 12124 34406
rect 12072 34342 12124 34348
rect 12084 34202 12112 34342
rect 13188 34202 13216 34954
rect 13544 34944 13596 34950
rect 13544 34886 13596 34892
rect 13556 34678 13584 34886
rect 13544 34672 13596 34678
rect 13544 34614 13596 34620
rect 13268 34400 13320 34406
rect 13268 34342 13320 34348
rect 10600 34196 10652 34202
rect 10600 34138 10652 34144
rect 12072 34196 12124 34202
rect 12072 34138 12124 34144
rect 13176 34196 13228 34202
rect 13176 34138 13228 34144
rect 12084 33658 12112 34138
rect 13280 34066 13308 34342
rect 14200 34202 14228 35090
rect 14556 34604 14608 34610
rect 14556 34546 14608 34552
rect 14188 34196 14240 34202
rect 14188 34138 14240 34144
rect 13912 34128 13964 34134
rect 13912 34070 13964 34076
rect 13268 34060 13320 34066
rect 13268 34002 13320 34008
rect 13924 33658 13952 34070
rect 14568 33658 14596 34546
rect 12072 33652 12124 33658
rect 12072 33594 12124 33600
rect 13912 33652 13964 33658
rect 13912 33594 13964 33600
rect 14556 33652 14608 33658
rect 14556 33594 14608 33600
rect 14660 33522 14688 35634
rect 14936 35442 14964 35866
rect 15016 35624 15068 35630
rect 15120 35612 15148 38200
rect 15292 35692 15344 35698
rect 15292 35634 15344 35640
rect 15068 35584 15148 35612
rect 15016 35566 15068 35572
rect 14936 35414 15056 35442
rect 14740 34944 14792 34950
rect 14740 34886 14792 34892
rect 14752 34746 14780 34886
rect 14740 34740 14792 34746
rect 14740 34682 14792 34688
rect 14740 34196 14792 34202
rect 14740 34138 14792 34144
rect 14648 33516 14700 33522
rect 14648 33458 14700 33464
rect 14752 33386 14780 34138
rect 15028 34066 15056 35414
rect 15304 34746 15332 35634
rect 16868 35630 16896 38200
rect 18616 36242 18644 38200
rect 20640 37210 20668 38270
rect 22098 38200 22154 39000
rect 23846 38200 23902 39000
rect 25594 38298 25650 39000
rect 25594 38270 25912 38298
rect 25594 38200 25650 38270
rect 20640 37182 20760 37210
rect 20732 36242 20760 37182
rect 18604 36236 18656 36242
rect 18604 36178 18656 36184
rect 20720 36236 20772 36242
rect 20720 36178 20772 36184
rect 17592 36168 17644 36174
rect 17592 36110 17644 36116
rect 19340 36168 19392 36174
rect 19340 36110 19392 36116
rect 20812 36168 20864 36174
rect 20812 36110 20864 36116
rect 17224 36100 17276 36106
rect 17224 36042 17276 36048
rect 17236 35698 17264 36042
rect 17604 35894 17632 36110
rect 19248 36032 19300 36038
rect 19248 35974 19300 35980
rect 17604 35866 17816 35894
rect 17224 35692 17276 35698
rect 17224 35634 17276 35640
rect 16856 35624 16908 35630
rect 16856 35566 16908 35572
rect 17788 35306 17816 35866
rect 17604 35290 17816 35306
rect 17592 35284 17816 35290
rect 17644 35278 17816 35284
rect 17592 35226 17644 35232
rect 16764 35012 16816 35018
rect 16764 34954 16816 34960
rect 15292 34740 15344 34746
rect 15292 34682 15344 34688
rect 16776 34524 16804 34954
rect 16856 34944 16908 34950
rect 16856 34886 16908 34892
rect 16868 34746 16896 34886
rect 17788 34746 17816 35278
rect 19260 35154 19288 35974
rect 19352 35290 19380 36110
rect 19432 36032 19484 36038
rect 19432 35974 19484 35980
rect 19444 35766 19472 35974
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 20824 35766 20852 36110
rect 19432 35760 19484 35766
rect 19432 35702 19484 35708
rect 20812 35760 20864 35766
rect 20812 35702 20864 35708
rect 19984 35692 20036 35698
rect 19984 35634 20036 35640
rect 20352 35692 20404 35698
rect 20352 35634 20404 35640
rect 19340 35284 19392 35290
rect 19340 35226 19392 35232
rect 19248 35148 19300 35154
rect 19248 35090 19300 35096
rect 18972 35012 19024 35018
rect 18972 34954 19024 34960
rect 18420 34944 18472 34950
rect 18420 34886 18472 34892
rect 16856 34740 16908 34746
rect 16856 34682 16908 34688
rect 17776 34740 17828 34746
rect 17776 34682 17828 34688
rect 16856 34536 16908 34542
rect 16776 34496 16856 34524
rect 16856 34478 16908 34484
rect 15016 34060 15068 34066
rect 15016 34002 15068 34008
rect 16868 33658 16896 34478
rect 18432 34474 18460 34886
rect 18984 34746 19012 34954
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19996 34746 20024 35634
rect 20168 35012 20220 35018
rect 20168 34954 20220 34960
rect 20180 34746 20208 34954
rect 18972 34740 19024 34746
rect 18972 34682 19024 34688
rect 19984 34740 20036 34746
rect 19984 34682 20036 34688
rect 20168 34740 20220 34746
rect 20168 34682 20220 34688
rect 18512 34536 18564 34542
rect 18512 34478 18564 34484
rect 18420 34468 18472 34474
rect 18420 34410 18472 34416
rect 18524 33862 18552 34478
rect 17316 33856 17368 33862
rect 17316 33798 17368 33804
rect 18512 33856 18564 33862
rect 18512 33798 18564 33804
rect 17328 33658 17356 33798
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 16856 33652 16908 33658
rect 16856 33594 16908 33600
rect 17316 33652 17368 33658
rect 17316 33594 17368 33600
rect 14740 33380 14792 33386
rect 14740 33322 14792 33328
rect 10876 31816 10928 31822
rect 10876 31758 10928 31764
rect 10888 29850 10916 31758
rect 10876 29844 10928 29850
rect 10876 29786 10928 29792
rect 13452 29640 13504 29646
rect 13452 29582 13504 29588
rect 13464 27130 13492 29582
rect 13452 27124 13504 27130
rect 13452 27066 13504 27072
rect 9588 27056 9640 27062
rect 9588 26998 9640 27004
rect 8300 26920 8352 26926
rect 8300 26862 8352 26868
rect 6920 26376 6972 26382
rect 6920 26318 6972 26324
rect 8312 26042 8340 26862
rect 17328 26790 17356 33594
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19248 28960 19300 28966
rect 19248 28902 19300 28908
rect 19260 28558 19288 28902
rect 20364 28762 20392 35634
rect 22112 35630 22140 38200
rect 22284 36168 22336 36174
rect 22284 36110 22336 36116
rect 22296 35834 22324 36110
rect 22744 36100 22796 36106
rect 22744 36042 22796 36048
rect 22284 35828 22336 35834
rect 22284 35770 22336 35776
rect 22756 35698 22784 36042
rect 22744 35692 22796 35698
rect 22744 35634 22796 35640
rect 23860 35630 23888 38200
rect 25884 36242 25912 38270
rect 27342 38200 27398 39000
rect 29090 38298 29146 39000
rect 29090 38270 29408 38298
rect 29090 38200 29146 38270
rect 25872 36236 25924 36242
rect 25872 36178 25924 36184
rect 24032 36168 24084 36174
rect 24032 36110 24084 36116
rect 25964 36168 26016 36174
rect 25964 36110 26016 36116
rect 21916 35624 21968 35630
rect 21916 35566 21968 35572
rect 22100 35624 22152 35630
rect 22100 35566 22152 35572
rect 23848 35624 23900 35630
rect 23848 35566 23900 35572
rect 21180 34944 21232 34950
rect 21180 34886 21232 34892
rect 21192 34610 21220 34886
rect 21928 34610 21956 35566
rect 23388 35488 23440 35494
rect 23388 35430 23440 35436
rect 22928 35080 22980 35086
rect 22928 35022 22980 35028
rect 22100 35012 22152 35018
rect 22100 34954 22152 34960
rect 21180 34604 21232 34610
rect 21180 34546 21232 34552
rect 21916 34604 21968 34610
rect 21916 34546 21968 34552
rect 22112 34202 22140 34954
rect 22376 34672 22428 34678
rect 22376 34614 22428 34620
rect 22100 34196 22152 34202
rect 22100 34138 22152 34144
rect 22388 34066 22416 34614
rect 22940 34202 22968 35022
rect 23400 34610 23428 35430
rect 23940 35012 23992 35018
rect 23940 34954 23992 34960
rect 23952 34746 23980 34954
rect 24044 34746 24072 36110
rect 24860 36100 24912 36106
rect 24860 36042 24912 36048
rect 24872 35698 24900 36042
rect 24860 35692 24912 35698
rect 24860 35634 24912 35640
rect 24768 35556 24820 35562
rect 24768 35498 24820 35504
rect 24216 34944 24268 34950
rect 24216 34886 24268 34892
rect 24228 34746 24256 34886
rect 24780 34746 24808 35498
rect 24860 34944 24912 34950
rect 24860 34886 24912 34892
rect 24872 34746 24900 34886
rect 23940 34740 23992 34746
rect 23940 34682 23992 34688
rect 24032 34740 24084 34746
rect 24032 34682 24084 34688
rect 24216 34740 24268 34746
rect 24216 34682 24268 34688
rect 24768 34740 24820 34746
rect 24768 34682 24820 34688
rect 24860 34740 24912 34746
rect 24860 34682 24912 34688
rect 23388 34604 23440 34610
rect 23388 34546 23440 34552
rect 22928 34196 22980 34202
rect 22928 34138 22980 34144
rect 23400 34134 23428 34546
rect 25412 34536 25464 34542
rect 25412 34478 25464 34484
rect 25424 34202 25452 34478
rect 25976 34474 26004 36110
rect 27068 36032 27120 36038
rect 27068 35974 27120 35980
rect 26148 35012 26200 35018
rect 26148 34954 26200 34960
rect 26160 34746 26188 34954
rect 26148 34740 26200 34746
rect 26148 34682 26200 34688
rect 27080 34610 27108 35974
rect 27356 35630 27384 38200
rect 29380 36310 29408 38270
rect 30838 38200 30894 39000
rect 32586 38298 32642 39000
rect 34334 38298 34390 39000
rect 36082 38298 36138 39000
rect 32586 38270 32904 38298
rect 32586 38200 32642 38270
rect 29368 36304 29420 36310
rect 29368 36246 29420 36252
rect 29092 36168 29144 36174
rect 29092 36110 29144 36116
rect 27528 35692 27580 35698
rect 27528 35634 27580 35640
rect 27344 35624 27396 35630
rect 27344 35566 27396 35572
rect 27436 35012 27488 35018
rect 27436 34954 27488 34960
rect 27068 34604 27120 34610
rect 27068 34546 27120 34552
rect 26608 34536 26660 34542
rect 26608 34478 26660 34484
rect 26700 34536 26752 34542
rect 26700 34478 26752 34484
rect 25964 34468 26016 34474
rect 25964 34410 26016 34416
rect 25976 34202 26004 34410
rect 25412 34196 25464 34202
rect 25412 34138 25464 34144
rect 25964 34196 26016 34202
rect 25964 34138 26016 34144
rect 23388 34128 23440 34134
rect 23388 34070 23440 34076
rect 26620 34066 26648 34478
rect 22376 34060 22428 34066
rect 22376 34002 22428 34008
rect 26608 34060 26660 34066
rect 26608 34002 26660 34008
rect 26712 33862 26740 34478
rect 27448 34202 27476 34954
rect 27540 34746 27568 35634
rect 28540 35012 28592 35018
rect 28540 34954 28592 34960
rect 27896 34944 27948 34950
rect 27896 34886 27948 34892
rect 27908 34746 27936 34886
rect 28552 34746 28580 34954
rect 29104 34746 29132 36110
rect 29552 36032 29604 36038
rect 29552 35974 29604 35980
rect 27528 34740 27580 34746
rect 27528 34682 27580 34688
rect 27896 34740 27948 34746
rect 27896 34682 27948 34688
rect 28540 34740 28592 34746
rect 28540 34682 28592 34688
rect 29092 34740 29144 34746
rect 29092 34682 29144 34688
rect 27436 34196 27488 34202
rect 27436 34138 27488 34144
rect 28724 34060 28776 34066
rect 28724 34002 28776 34008
rect 28080 33992 28132 33998
rect 28080 33934 28132 33940
rect 26700 33856 26752 33862
rect 26700 33798 26752 33804
rect 27988 33856 28040 33862
rect 27988 33798 28040 33804
rect 28000 33590 28028 33798
rect 27988 33584 28040 33590
rect 27988 33526 28040 33532
rect 28092 33522 28120 33934
rect 28736 33658 28764 34002
rect 29184 33856 29236 33862
rect 29184 33798 29236 33804
rect 28724 33652 28776 33658
rect 28724 33594 28776 33600
rect 28080 33516 28132 33522
rect 28080 33458 28132 33464
rect 29196 32978 29224 33798
rect 29564 33522 29592 35974
rect 30472 35692 30524 35698
rect 30472 35634 30524 35640
rect 29920 35488 29972 35494
rect 29920 35430 29972 35436
rect 29932 35086 29960 35430
rect 29920 35080 29972 35086
rect 29920 35022 29972 35028
rect 29644 34536 29696 34542
rect 29644 34478 29696 34484
rect 29656 34066 29684 34478
rect 29644 34060 29696 34066
rect 29644 34002 29696 34008
rect 29656 33658 29684 34002
rect 29644 33652 29696 33658
rect 29644 33594 29696 33600
rect 29552 33516 29604 33522
rect 29552 33458 29604 33464
rect 29184 32972 29236 32978
rect 29184 32914 29236 32920
rect 20444 29096 20496 29102
rect 20444 29038 20496 29044
rect 20352 28756 20404 28762
rect 20352 28698 20404 28704
rect 19248 28552 19300 28558
rect 19248 28494 19300 28500
rect 19260 27062 19288 28494
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19248 27056 19300 27062
rect 19248 26998 19300 27004
rect 17316 26784 17368 26790
rect 17316 26726 17368 26732
rect 17868 26784 17920 26790
rect 17868 26726 17920 26732
rect 17328 26314 17356 26726
rect 8392 26308 8444 26314
rect 8392 26250 8444 26256
rect 17316 26308 17368 26314
rect 17316 26250 17368 26256
rect 8300 26036 8352 26042
rect 8300 25978 8352 25984
rect 8404 25906 8432 26250
rect 8392 25900 8444 25906
rect 8392 25842 8444 25848
rect 4988 25764 5040 25770
rect 4988 25706 5040 25712
rect 4896 25696 4948 25702
rect 4896 25638 4948 25644
rect 4908 25498 4936 25638
rect 4896 25492 4948 25498
rect 4896 25434 4948 25440
rect 4804 24744 4856 24750
rect 4804 24686 4856 24692
rect 4712 24200 4764 24206
rect 4712 24142 4764 24148
rect 4620 22568 4672 22574
rect 4620 22510 4672 22516
rect 4160 22500 4212 22506
rect 4160 22442 4212 22448
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4620 21888 4672 21894
rect 4620 21830 4672 21836
rect 4632 21486 4660 21830
rect 4068 21480 4120 21486
rect 4068 21422 4120 21428
rect 4620 21480 4672 21486
rect 4620 21422 4672 21428
rect 3976 21412 4028 21418
rect 3976 21354 4028 21360
rect 3608 21344 3660 21350
rect 3608 21286 3660 21292
rect 3516 20800 3568 20806
rect 3516 20742 3568 20748
rect 3528 20398 3556 20742
rect 3516 20392 3568 20398
rect 3516 20334 3568 20340
rect 3424 19508 3476 19514
rect 3424 19450 3476 19456
rect 3528 19242 3556 20334
rect 3516 19236 3568 19242
rect 3516 19178 3568 19184
rect 3424 19168 3476 19174
rect 3424 19110 3476 19116
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 3344 17678 3372 18566
rect 3436 18358 3464 19110
rect 3620 18766 3648 21286
rect 4080 21010 4108 21422
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4632 21078 4660 21422
rect 4620 21072 4672 21078
rect 4620 21014 4672 21020
rect 4068 21004 4120 21010
rect 4068 20946 4120 20952
rect 4080 19378 4108 20946
rect 4344 20936 4396 20942
rect 4344 20878 4396 20884
rect 4356 20398 4384 20878
rect 4528 20800 4580 20806
rect 4528 20742 4580 20748
rect 4540 20534 4568 20742
rect 4528 20528 4580 20534
rect 4528 20470 4580 20476
rect 4344 20392 4396 20398
rect 4344 20334 4396 20340
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 17328 19514 17356 26250
rect 17316 19508 17368 19514
rect 17316 19450 17368 19456
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 3608 18760 3660 18766
rect 3608 18702 3660 18708
rect 4344 18760 4396 18766
rect 4344 18702 4396 18708
rect 4620 18760 4672 18766
rect 4620 18702 4672 18708
rect 4356 18426 4384 18702
rect 4344 18420 4396 18426
rect 4344 18362 4396 18368
rect 3424 18352 3476 18358
rect 3424 18294 3476 18300
rect 3792 18148 3844 18154
rect 3792 18090 3844 18096
rect 3332 17672 3384 17678
rect 3332 17614 3384 17620
rect 3804 17354 3832 18090
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 3884 17536 3936 17542
rect 3884 17478 3936 17484
rect 3620 17326 3832 17354
rect 3516 16652 3568 16658
rect 3516 16594 3568 16600
rect 3252 16546 3464 16574
rect 2596 16526 2648 16532
rect 2608 16250 2636 16526
rect 2872 16448 2924 16454
rect 2872 16390 2924 16396
rect 3240 16448 3292 16454
rect 3240 16390 3292 16396
rect 2884 16250 2912 16390
rect 2596 16244 2648 16250
rect 2596 16186 2648 16192
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 3252 15706 3280 16390
rect 3240 15700 3292 15706
rect 3240 15642 3292 15648
rect 2872 15632 2924 15638
rect 2872 15574 2924 15580
rect 2596 15428 2648 15434
rect 2596 15370 2648 15376
rect 1582 15328 1638 15337
rect 1582 15263 1638 15272
rect 1596 15094 1624 15263
rect 1584 15088 1636 15094
rect 1584 15030 1636 15036
rect 2608 15026 2636 15370
rect 2688 15360 2740 15366
rect 2688 15302 2740 15308
rect 2596 15020 2648 15026
rect 2596 14962 2648 14968
rect 1952 14952 2004 14958
rect 1952 14894 2004 14900
rect 1964 14618 1992 14894
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 2596 13864 2648 13870
rect 2596 13806 2648 13812
rect 938 13696 994 13705
rect 938 13631 994 13640
rect 952 13394 980 13631
rect 940 13388 992 13394
rect 940 13330 992 13336
rect 2608 13326 2636 13806
rect 2596 13320 2648 13326
rect 2596 13262 2648 13268
rect 1952 12844 2004 12850
rect 1952 12786 2004 12792
rect 938 12064 994 12073
rect 938 11999 994 12008
rect 952 11830 980 11999
rect 940 11824 992 11830
rect 940 11766 992 11772
rect 1964 11218 1992 12786
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2608 11762 2636 12038
rect 2596 11756 2648 11762
rect 2596 11698 2648 11704
rect 1952 11212 2004 11218
rect 1952 11154 2004 11160
rect 938 10432 994 10441
rect 938 10367 994 10376
rect 952 10130 980 10367
rect 940 10124 992 10130
rect 940 10066 992 10072
rect 1964 9586 1992 11154
rect 2596 10464 2648 10470
rect 2596 10406 2648 10412
rect 2608 10062 2636 10406
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 1952 9580 2004 9586
rect 1952 9522 2004 9528
rect 938 8800 994 8809
rect 938 8735 994 8744
rect 952 8566 980 8735
rect 940 8560 992 8566
rect 940 8502 992 8508
rect 1964 7954 1992 9522
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 2608 8498 2636 8774
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 1952 7948 2004 7954
rect 1952 7890 2004 7896
rect 1964 7410 1992 7890
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 1582 7032 1638 7041
rect 1582 6967 1638 6976
rect 1596 6390 1624 6967
rect 1584 6384 1636 6390
rect 1584 6326 1636 6332
rect 2596 6316 2648 6322
rect 2596 6258 2648 6264
rect 2608 5914 2636 6258
rect 2596 5908 2648 5914
rect 2596 5850 2648 5856
rect 938 5536 994 5545
rect 938 5471 994 5480
rect 952 4690 980 5471
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 940 4684 992 4690
rect 940 4626 992 4632
rect 2608 4622 2636 4966
rect 2596 4616 2648 4622
rect 2596 4558 2648 4564
rect 2596 3936 2648 3942
rect 938 3904 994 3913
rect 2596 3878 2648 3884
rect 938 3839 994 3848
rect 952 3602 980 3839
rect 940 3596 992 3602
rect 940 3538 992 3544
rect 2608 3534 2636 3878
rect 2596 3528 2648 3534
rect 2596 3470 2648 3476
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 1584 2984 1636 2990
rect 1584 2926 1636 2932
rect 1596 2689 1624 2926
rect 1768 2848 1820 2854
rect 1768 2790 1820 2796
rect 1582 2680 1638 2689
rect 1582 2615 1638 2624
rect 1780 800 1808 2790
rect 2608 2514 2636 2994
rect 2596 2508 2648 2514
rect 2596 2450 2648 2456
rect 2700 2446 2728 15302
rect 2884 13530 2912 15574
rect 2964 13728 3016 13734
rect 2964 13670 3016 13676
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2976 12850 3004 13670
rect 3436 13394 3464 16546
rect 3528 14482 3556 16594
rect 3620 14906 3648 17326
rect 3700 17196 3752 17202
rect 3700 17138 3752 17144
rect 3712 15706 3740 17138
rect 3896 16590 3924 17478
rect 4632 17202 4660 18702
rect 4712 18080 4764 18086
rect 4712 18022 4764 18028
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 4620 16992 4672 16998
rect 4620 16934 4672 16940
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 3700 15700 3752 15706
rect 3700 15642 3752 15648
rect 3620 14878 3740 14906
rect 3896 14890 3924 16526
rect 4252 16516 4304 16522
rect 4252 16458 4304 16464
rect 4264 16250 4292 16458
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 4068 16176 4120 16182
rect 4068 16118 4120 16124
rect 4080 15366 4108 16118
rect 4632 16114 4660 16934
rect 4724 16182 4752 18022
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 7564 17536 7616 17542
rect 7564 17478 7616 17484
rect 7576 17338 7604 17478
rect 7564 17332 7616 17338
rect 7564 17274 7616 17280
rect 4896 17128 4948 17134
rect 4896 17070 4948 17076
rect 4712 16176 4764 16182
rect 4712 16118 4764 16124
rect 4620 16108 4672 16114
rect 4620 16050 4672 16056
rect 4908 15978 4936 17070
rect 6552 16448 6604 16454
rect 6552 16390 6604 16396
rect 4896 15972 4948 15978
rect 4896 15914 4948 15920
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4068 15360 4120 15366
rect 4068 15302 4120 15308
rect 3976 14952 4028 14958
rect 3976 14894 4028 14900
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3620 14618 3648 14758
rect 3608 14612 3660 14618
rect 3608 14554 3660 14560
rect 3516 14476 3568 14482
rect 3516 14418 3568 14424
rect 3424 13388 3476 13394
rect 3424 13330 3476 13336
rect 3528 12850 3556 14418
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 3516 12844 3568 12850
rect 3516 12786 3568 12792
rect 3424 12640 3476 12646
rect 3424 12582 3476 12588
rect 3436 12306 3464 12582
rect 3424 12300 3476 12306
rect 3424 12242 3476 12248
rect 3436 11558 3464 12242
rect 3712 11762 3740 14878
rect 3884 14884 3936 14890
rect 3884 14826 3936 14832
rect 3988 14618 4016 14894
rect 4080 14822 4108 15302
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 3792 14272 3844 14278
rect 3792 14214 3844 14220
rect 3804 13802 3832 14214
rect 4080 13870 4108 14758
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 3792 13796 3844 13802
rect 3792 13738 3844 13744
rect 3792 13320 3844 13326
rect 3792 13262 3844 13268
rect 3804 12986 3832 13262
rect 3792 12980 3844 12986
rect 3792 12922 3844 12928
rect 3700 11756 3752 11762
rect 3700 11698 3752 11704
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 2884 10554 2912 11494
rect 3620 11354 3648 11494
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 3516 11008 3568 11014
rect 3516 10950 3568 10956
rect 2884 10526 3004 10554
rect 2872 10464 2924 10470
rect 2872 10406 2924 10412
rect 2884 10266 2912 10406
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 2792 7886 2820 8230
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2792 5778 2820 6598
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 2884 5234 2912 6054
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2976 4146 3004 10526
rect 3528 10062 3556 10950
rect 3608 10464 3660 10470
rect 3608 10406 3660 10412
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 3620 9654 3648 10406
rect 3608 9648 3660 9654
rect 3608 9590 3660 9596
rect 3712 9466 3740 11698
rect 4080 11558 4108 13806
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 6564 13394 6592 16390
rect 11900 15638 11928 17614
rect 14280 16652 14332 16658
rect 14280 16594 14332 16600
rect 13268 16516 13320 16522
rect 13268 16458 13320 16464
rect 13280 16250 13308 16458
rect 13268 16244 13320 16250
rect 13268 16186 13320 16192
rect 12808 16176 12860 16182
rect 12808 16118 12860 16124
rect 12820 15706 12848 16118
rect 13084 15972 13136 15978
rect 13084 15914 13136 15920
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 11888 15632 11940 15638
rect 11888 15574 11940 15580
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 13096 13326 13124 15914
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 4436 13184 4488 13190
rect 4436 13126 4488 13132
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 4448 12986 4476 13126
rect 4436 12980 4488 12986
rect 4436 12922 4488 12928
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 4080 10470 4108 11494
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 3804 9722 3832 9998
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 3528 9438 3740 9466
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3436 9178 3464 9318
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3436 8634 3464 9114
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3344 6866 3372 7346
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3332 6860 3384 6866
rect 3332 6802 3384 6808
rect 3436 6322 3464 7142
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3528 5370 3556 9438
rect 4080 8362 4108 10406
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 7208 10130 7236 13126
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 10428 10044 10456 13126
rect 11072 10266 11100 13262
rect 13832 12918 13860 15302
rect 13820 12912 13872 12918
rect 13820 12854 13872 12860
rect 14292 12850 14320 16594
rect 17880 16250 17908 26726
rect 20456 26234 20484 29038
rect 29932 29034 29960 35022
rect 30104 35012 30156 35018
rect 30104 34954 30156 34960
rect 30010 34504 30066 34513
rect 30010 34439 30066 34448
rect 30024 34134 30052 34439
rect 30116 34202 30144 34954
rect 30104 34196 30156 34202
rect 30104 34138 30156 34144
rect 30012 34128 30064 34134
rect 30012 34070 30064 34076
rect 30484 33998 30512 35634
rect 30852 35630 30880 38200
rect 32876 36310 32904 38270
rect 34256 38270 34390 38298
rect 32864 36304 32916 36310
rect 32864 36246 32916 36252
rect 31576 36168 31628 36174
rect 31576 36110 31628 36116
rect 31668 36168 31720 36174
rect 31668 36110 31720 36116
rect 34152 36168 34204 36174
rect 34152 36110 34204 36116
rect 30840 35624 30892 35630
rect 30840 35566 30892 35572
rect 31588 35290 31616 36110
rect 31680 35766 31708 36110
rect 33692 36100 33744 36106
rect 33692 36042 33744 36048
rect 33600 36032 33652 36038
rect 33600 35974 33652 35980
rect 31668 35760 31720 35766
rect 31668 35702 31720 35708
rect 33612 35714 33640 35974
rect 33704 35894 33732 36042
rect 33704 35866 33824 35894
rect 33612 35698 33732 35714
rect 33612 35692 33744 35698
rect 33612 35686 33692 35692
rect 33692 35634 33744 35640
rect 33796 35578 33824 35866
rect 32496 35556 32548 35562
rect 32496 35498 32548 35504
rect 33704 35550 33824 35578
rect 31576 35284 31628 35290
rect 31576 35226 31628 35232
rect 31392 35012 31444 35018
rect 31392 34954 31444 34960
rect 31208 34944 31260 34950
rect 31208 34886 31260 34892
rect 30932 34400 30984 34406
rect 30932 34342 30984 34348
rect 30472 33992 30524 33998
rect 30472 33934 30524 33940
rect 30656 33856 30708 33862
rect 30656 33798 30708 33804
rect 30668 33454 30696 33798
rect 30944 33522 30972 34342
rect 31220 33522 31248 34886
rect 31404 34542 31432 34954
rect 32128 34944 32180 34950
rect 32128 34886 32180 34892
rect 31668 34604 31720 34610
rect 31668 34546 31720 34552
rect 31944 34604 31996 34610
rect 31944 34546 31996 34552
rect 31392 34536 31444 34542
rect 31392 34478 31444 34484
rect 30932 33516 30984 33522
rect 30932 33458 30984 33464
rect 31208 33516 31260 33522
rect 31208 33458 31260 33464
rect 30656 33448 30708 33454
rect 30656 33390 30708 33396
rect 31680 33017 31708 34546
rect 31760 33992 31812 33998
rect 31760 33934 31812 33940
rect 31772 33658 31800 33934
rect 31760 33652 31812 33658
rect 31760 33594 31812 33600
rect 31956 33590 31984 34546
rect 32034 34504 32090 34513
rect 32034 34439 32090 34448
rect 31944 33584 31996 33590
rect 31944 33526 31996 33532
rect 31666 33008 31722 33017
rect 31666 32943 31722 32952
rect 32048 32910 32076 34439
rect 32036 32904 32088 32910
rect 32036 32846 32088 32852
rect 31944 32836 31996 32842
rect 31944 32778 31996 32784
rect 30288 32768 30340 32774
rect 30288 32710 30340 32716
rect 30300 32298 30328 32710
rect 30656 32360 30708 32366
rect 30656 32302 30708 32308
rect 30288 32292 30340 32298
rect 30288 32234 30340 32240
rect 30300 32026 30328 32234
rect 30668 32026 30696 32302
rect 30288 32020 30340 32026
rect 30288 31962 30340 31968
rect 30656 32020 30708 32026
rect 30656 31962 30708 31968
rect 31956 31346 31984 32778
rect 32140 31890 32168 34886
rect 32404 34196 32456 34202
rect 32404 34138 32456 34144
rect 32416 33522 32444 34138
rect 32404 33516 32456 33522
rect 32404 33458 32456 33464
rect 32416 33130 32444 33458
rect 32324 33102 32444 33130
rect 32508 33114 32536 35498
rect 33324 35284 33376 35290
rect 33324 35226 33376 35232
rect 33336 34678 33364 35226
rect 33416 35216 33468 35222
rect 33416 35158 33468 35164
rect 33324 34672 33376 34678
rect 33324 34614 33376 34620
rect 32956 34604 33008 34610
rect 32956 34546 33008 34552
rect 32588 33516 32640 33522
rect 32588 33458 32640 33464
rect 32496 33108 32548 33114
rect 32324 32910 32352 33102
rect 32496 33050 32548 33056
rect 32404 33040 32456 33046
rect 32404 32982 32456 32988
rect 32312 32904 32364 32910
rect 32312 32846 32364 32852
rect 32128 31884 32180 31890
rect 32128 31826 32180 31832
rect 31944 31340 31996 31346
rect 31944 31282 31996 31288
rect 32416 30802 32444 32982
rect 32600 32026 32628 33458
rect 32968 33114 32996 34546
rect 33428 34066 33456 35158
rect 33416 34060 33468 34066
rect 33416 34002 33468 34008
rect 33232 33992 33284 33998
rect 33232 33934 33284 33940
rect 33140 33652 33192 33658
rect 33140 33594 33192 33600
rect 32956 33108 33008 33114
rect 32956 33050 33008 33056
rect 32772 33040 32824 33046
rect 32772 32982 32824 32988
rect 32588 32020 32640 32026
rect 32588 31962 32640 31968
rect 32784 31822 32812 32982
rect 32772 31816 32824 31822
rect 32772 31758 32824 31764
rect 32404 30796 32456 30802
rect 32404 30738 32456 30744
rect 32784 29306 32812 31758
rect 33152 30258 33180 33594
rect 33244 32570 33272 33934
rect 33600 33924 33652 33930
rect 33600 33866 33652 33872
rect 33324 33040 33376 33046
rect 33324 32982 33376 32988
rect 33232 32564 33284 32570
rect 33232 32506 33284 32512
rect 33336 32026 33364 32982
rect 33612 32910 33640 33866
rect 33600 32904 33652 32910
rect 33600 32846 33652 32852
rect 33704 32366 33732 35550
rect 34164 34950 34192 36110
rect 34152 34944 34204 34950
rect 34152 34886 34204 34892
rect 34060 34604 34112 34610
rect 34060 34546 34112 34552
rect 33968 33516 34020 33522
rect 33968 33458 34020 33464
rect 33692 32360 33744 32366
rect 33692 32302 33744 32308
rect 33980 32230 34008 33458
rect 33968 32224 34020 32230
rect 33968 32166 34020 32172
rect 33324 32020 33376 32026
rect 33324 31962 33376 31968
rect 33508 31272 33560 31278
rect 33508 31214 33560 31220
rect 33416 31204 33468 31210
rect 33416 31146 33468 31152
rect 33428 30938 33456 31146
rect 33416 30932 33468 30938
rect 33416 30874 33468 30880
rect 33140 30252 33192 30258
rect 33140 30194 33192 30200
rect 32772 29300 32824 29306
rect 32772 29242 32824 29248
rect 30380 29164 30432 29170
rect 30380 29106 30432 29112
rect 28448 29028 28500 29034
rect 28448 28970 28500 28976
rect 29920 29028 29972 29034
rect 29920 28970 29972 28976
rect 20364 26206 20484 26234
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 20364 26042 20392 26206
rect 20352 26036 20404 26042
rect 20352 25978 20404 25984
rect 19432 25832 19484 25838
rect 19432 25774 19484 25780
rect 19444 22030 19472 25774
rect 28460 25770 28488 28970
rect 29000 26376 29052 26382
rect 29000 26318 29052 26324
rect 20260 25764 20312 25770
rect 20260 25706 20312 25712
rect 28448 25764 28500 25770
rect 28448 25706 28500 25712
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 20272 19514 20300 25706
rect 29012 23322 29040 26318
rect 29644 25288 29696 25294
rect 29644 25230 29696 25236
rect 29000 23316 29052 23322
rect 29000 23258 29052 23264
rect 28356 23112 28408 23118
rect 28356 23054 28408 23060
rect 24124 22024 24176 22030
rect 24124 21966 24176 21972
rect 20352 21956 20404 21962
rect 20352 21898 20404 21904
rect 20364 20602 20392 21898
rect 20352 20596 20404 20602
rect 20352 20538 20404 20544
rect 22008 20324 22060 20330
rect 22008 20266 22060 20272
rect 20260 19508 20312 19514
rect 20260 19450 20312 19456
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 16120 16244 16172 16250
rect 16120 16186 16172 16192
rect 17868 16244 17920 16250
rect 17868 16186 17920 16192
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 10336 10016 10456 10044
rect 4436 9920 4488 9926
rect 4436 9862 4488 9868
rect 4448 9586 4476 9862
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4448 7290 4476 7686
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 4448 7262 4660 7290
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3792 7200 3844 7206
rect 3792 7142 3844 7148
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3620 5914 3648 6190
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3712 5710 3740 7142
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3804 5302 3832 7142
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4632 6866 4660 7262
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4724 6730 4752 7414
rect 5460 7342 5488 8230
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 4804 7268 4856 7274
rect 4804 7210 4856 7216
rect 4816 7002 4844 7210
rect 4804 6996 4856 7002
rect 4804 6938 4856 6944
rect 5000 6934 5028 7278
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 4988 6928 5040 6934
rect 4988 6870 5040 6876
rect 4712 6724 4764 6730
rect 4712 6666 4764 6672
rect 5000 6458 5028 6870
rect 5184 6798 5212 7142
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 5460 6662 5488 7278
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 3792 5296 3844 5302
rect 3792 5238 3844 5244
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 5460 4554 5488 6598
rect 5448 4548 5500 4554
rect 5448 4490 5500 4496
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 8680 3534 8708 9658
rect 9312 5636 9364 5642
rect 9312 5578 9364 5584
rect 9324 4146 9352 5578
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9968 5166 9996 5510
rect 9956 5160 10008 5166
rect 9956 5102 10008 5108
rect 9968 5030 9996 5102
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 9784 4758 9812 4966
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 9968 4554 9996 4966
rect 9956 4548 10008 4554
rect 9956 4490 10008 4496
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 6644 3460 6696 3466
rect 6644 3402 6696 3408
rect 8300 3460 8352 3466
rect 8300 3402 8352 3408
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 6092 2508 6144 2514
rect 6092 2450 6144 2456
rect 2688 2440 2740 2446
rect 2688 2382 2740 2388
rect 3332 2440 3384 2446
rect 3332 2382 3384 2388
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 3344 1306 3372 2382
rect 3252 1278 3372 1306
rect 3252 800 3280 1278
rect 4724 800 4752 2382
rect 6104 1170 6132 2450
rect 6656 2446 6684 3402
rect 8312 3194 8340 3402
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 9968 3058 9996 4490
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 10152 3602 10180 4082
rect 10336 3670 10364 10016
rect 14292 8090 14320 12786
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 10416 7812 10468 7818
rect 10416 7754 10468 7760
rect 10428 7546 10456 7754
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 10888 5574 10916 5646
rect 10876 5568 10928 5574
rect 10876 5510 10928 5516
rect 10600 5024 10652 5030
rect 10600 4966 10652 4972
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10612 4622 10640 4966
rect 10600 4616 10652 4622
rect 10600 4558 10652 4564
rect 10600 4072 10652 4078
rect 10600 4014 10652 4020
rect 10324 3664 10376 3670
rect 10324 3606 10376 3612
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 6104 1142 6224 1170
rect 6196 800 6224 1142
rect 7668 800 7696 2926
rect 8772 2446 8800 2926
rect 9128 2508 9180 2514
rect 9128 2450 9180 2456
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 9140 800 9168 2450
rect 10612 800 10640 4014
rect 10704 3534 10732 4966
rect 10980 4826 11008 5646
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 11256 5166 11284 5510
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 11072 3466 11100 4422
rect 11900 4146 11928 5714
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 11060 3460 11112 3466
rect 11060 3402 11112 3408
rect 11992 3058 12020 5510
rect 12084 4690 12112 8026
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 13544 5840 13596 5846
rect 13544 5782 13596 5788
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 13084 5704 13136 5710
rect 13084 5646 13136 5652
rect 12072 4684 12124 4690
rect 12072 4626 12124 4632
rect 12084 4282 12112 4626
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 12084 3602 12112 4218
rect 12176 3738 12204 5646
rect 13096 5370 13124 5646
rect 13084 5364 13136 5370
rect 13084 5306 13136 5312
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 12256 5092 12308 5098
rect 12256 5034 12308 5040
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 12072 3596 12124 3602
rect 12072 3538 12124 3544
rect 12072 3460 12124 3466
rect 12072 3402 12124 3408
rect 12084 3194 12112 3402
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 12268 3058 12296 5034
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 12256 3052 12308 3058
rect 12256 2994 12308 3000
rect 11152 2984 11204 2990
rect 11152 2926 11204 2932
rect 11164 2446 11192 2926
rect 12452 2650 12480 4558
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12544 2514 12572 4422
rect 12636 2514 12664 4966
rect 13096 4826 13124 5102
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 13556 4690 13584 5782
rect 14016 5642 14044 6054
rect 14464 5840 14516 5846
rect 14464 5782 14516 5788
rect 14004 5636 14056 5642
rect 14004 5578 14056 5584
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 13728 5160 13780 5166
rect 13728 5102 13780 5108
rect 13544 4684 13596 4690
rect 13544 4626 13596 4632
rect 13176 4616 13228 4622
rect 13176 4558 13228 4564
rect 13188 4282 13216 4558
rect 13176 4276 13228 4282
rect 13176 4218 13228 4224
rect 13636 4072 13688 4078
rect 13740 4060 13768 5102
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13688 4032 13768 4060
rect 13636 4014 13688 4020
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 12084 800 12112 2450
rect 12912 2446 12940 2926
rect 13740 2922 13768 4032
rect 13832 3738 13860 4558
rect 14096 4480 14148 4486
rect 14096 4422 14148 4428
rect 13820 3732 13872 3738
rect 13820 3674 13872 3680
rect 14108 3058 14136 4422
rect 14384 4146 14412 5510
rect 14476 5370 14504 5782
rect 15752 5636 15804 5642
rect 15752 5578 15804 5584
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 14924 5364 14976 5370
rect 14924 5306 14976 5312
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14476 3942 14504 5102
rect 14936 4690 14964 5306
rect 14924 4684 14976 4690
rect 14924 4626 14976 4632
rect 14648 4140 14700 4146
rect 14648 4082 14700 4088
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14660 3738 14688 4082
rect 15016 4072 15068 4078
rect 15016 4014 15068 4020
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14556 3392 14608 3398
rect 14556 3334 14608 3340
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 13728 2916 13780 2922
rect 13728 2858 13780 2864
rect 14568 2514 14596 3334
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 13544 2372 13596 2378
rect 13544 2314 13596 2320
rect 13556 800 13584 2314
rect 15028 800 15056 4014
rect 15212 3534 15240 5510
rect 15764 5370 15792 5578
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 16132 5302 16160 16186
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17236 10674 17264 12582
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 17224 10668 17276 10674
rect 17224 10610 17276 10616
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 16856 10056 16908 10062
rect 16856 9998 16908 10004
rect 16488 5840 16540 5846
rect 16488 5782 16540 5788
rect 16120 5296 16172 5302
rect 16120 5238 16172 5244
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15304 3126 15332 4082
rect 15292 3120 15344 3126
rect 15292 3062 15344 3068
rect 15200 2984 15252 2990
rect 15200 2926 15252 2932
rect 15212 2446 15240 2926
rect 15488 2650 15516 5102
rect 16500 4622 16528 5782
rect 16672 4684 16724 4690
rect 16672 4626 16724 4632
rect 16488 4616 16540 4622
rect 16488 4558 16540 4564
rect 15660 4480 15712 4486
rect 15660 4422 15712 4428
rect 15844 4480 15896 4486
rect 15844 4422 15896 4428
rect 15672 3058 15700 4422
rect 15856 3194 15884 4422
rect 15844 3188 15896 3194
rect 15844 3130 15896 3136
rect 15660 3052 15712 3058
rect 15660 2994 15712 3000
rect 16500 2650 16528 4558
rect 16684 3738 16712 4626
rect 16672 3732 16724 3738
rect 16672 3674 16724 3680
rect 15476 2644 15528 2650
rect 15476 2586 15528 2592
rect 16488 2644 16540 2650
rect 16488 2586 16540 2592
rect 16868 2582 16896 9998
rect 17132 9920 17184 9926
rect 17132 9862 17184 9868
rect 17144 9722 17172 9862
rect 17132 9716 17184 9722
rect 17132 9658 17184 9664
rect 19352 7954 19380 10406
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19340 7948 19392 7954
rect 19340 7890 19392 7896
rect 20272 7818 20300 19450
rect 21640 19372 21692 19378
rect 21640 19314 21692 19320
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20916 16726 20944 16934
rect 20904 16720 20956 16726
rect 20904 16662 20956 16668
rect 21456 16720 21508 16726
rect 21456 16662 21508 16668
rect 20444 16448 20496 16454
rect 20444 16390 20496 16396
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 20456 16114 20484 16390
rect 20732 16250 20760 16390
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20916 10062 20944 16662
rect 21468 15570 21496 16662
rect 21456 15564 21508 15570
rect 21456 15506 21508 15512
rect 21468 15162 21496 15506
rect 21456 15156 21508 15162
rect 21456 15098 21508 15104
rect 20904 10056 20956 10062
rect 20904 9998 20956 10004
rect 20260 7812 20312 7818
rect 20260 7754 20312 7760
rect 20628 7812 20680 7818
rect 20628 7754 20680 7760
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 19260 6254 19288 7686
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 20640 7546 20668 7754
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 18512 6248 18564 6254
rect 18512 6190 18564 6196
rect 19248 6248 19300 6254
rect 19248 6190 19300 6196
rect 18524 5098 18552 6190
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 18512 5092 18564 5098
rect 18512 5034 18564 5040
rect 17684 5024 17736 5030
rect 17684 4966 17736 4972
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 17224 4480 17276 4486
rect 17224 4422 17276 4428
rect 17316 4480 17368 4486
rect 17316 4422 17368 4428
rect 16948 4072 17000 4078
rect 16948 4014 17000 4020
rect 16960 2854 16988 4014
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 16856 2576 16908 2582
rect 16856 2518 16908 2524
rect 17236 2514 17264 4422
rect 17328 3058 17356 4422
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 17420 3194 17448 3470
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 17696 3126 17724 4966
rect 19248 4752 19300 4758
rect 19248 4694 19300 4700
rect 18236 4616 18288 4622
rect 18236 4558 18288 4564
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 17960 3460 18012 3466
rect 17960 3402 18012 3408
rect 17972 3194 18000 3402
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 17684 3120 17736 3126
rect 17684 3062 17736 3068
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 17224 2508 17276 2514
rect 17224 2450 17276 2456
rect 18064 2446 18092 4014
rect 18248 3738 18276 4558
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 18236 3732 18288 3738
rect 18236 3674 18288 3680
rect 18800 3466 18828 4422
rect 19156 4072 19208 4078
rect 19156 4014 19208 4020
rect 18788 3460 18840 3466
rect 18788 3402 18840 3408
rect 19168 3194 19196 4014
rect 19260 3602 19288 4694
rect 19352 4486 19380 4966
rect 19340 4480 19392 4486
rect 19340 4422 19392 4428
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19156 3188 19208 3194
rect 19156 3130 19208 3136
rect 19260 2650 19288 3538
rect 19352 2990 19380 4422
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19984 3936 20036 3942
rect 19984 3878 20036 3884
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19444 3194 19472 3334
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19432 3188 19484 3194
rect 19432 3130 19484 3136
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 19996 2650 20024 3878
rect 20628 3120 20680 3126
rect 20626 3088 20628 3097
rect 20680 3088 20682 3097
rect 20626 3023 20682 3032
rect 20076 2984 20128 2990
rect 20076 2926 20128 2932
rect 19248 2644 19300 2650
rect 19248 2586 19300 2592
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 18144 2508 18196 2514
rect 18144 2450 18196 2456
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 16304 2372 16356 2378
rect 16304 2314 16356 2320
rect 16316 1170 16344 2314
rect 18156 1170 18184 2450
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 16316 1142 16528 1170
rect 16500 800 16528 1142
rect 17972 1142 18184 1170
rect 17972 800 18000 1142
rect 19996 898 20024 2450
rect 20088 2446 20116 2926
rect 20732 2446 20760 6054
rect 20904 2984 20956 2990
rect 20904 2926 20956 2932
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 19444 870 19564 898
rect 19444 800 19472 870
rect 1766 0 1822 800
rect 3238 0 3294 800
rect 4710 0 4766 800
rect 6182 0 6238 800
rect 7654 0 7710 800
rect 9126 0 9182 800
rect 10598 0 10654 800
rect 12070 0 12126 800
rect 13542 0 13598 800
rect 15014 0 15070 800
rect 16486 0 16542 800
rect 17958 0 18014 800
rect 19430 0 19486 800
rect 19536 762 19564 870
rect 19904 870 20024 898
rect 19904 762 19932 870
rect 20916 800 20944 2926
rect 21652 1358 21680 19314
rect 21824 18216 21876 18222
rect 21824 18158 21876 18164
rect 21836 16250 21864 18158
rect 21916 17536 21968 17542
rect 21916 17478 21968 17484
rect 21928 16726 21956 17478
rect 21916 16720 21968 16726
rect 21916 16662 21968 16668
rect 21824 16244 21876 16250
rect 21824 16186 21876 16192
rect 21916 16108 21968 16114
rect 21916 16050 21968 16056
rect 21928 15706 21956 16050
rect 21916 15700 21968 15706
rect 21916 15642 21968 15648
rect 22020 15502 22048 20266
rect 22468 19304 22520 19310
rect 22468 19246 22520 19252
rect 22480 18426 22508 19246
rect 24136 18426 24164 21966
rect 28172 21888 28224 21894
rect 28172 21830 28224 21836
rect 28184 21622 28212 21830
rect 28172 21616 28224 21622
rect 28172 21558 28224 21564
rect 27528 21480 27580 21486
rect 27528 21422 27580 21428
rect 24400 19848 24452 19854
rect 24400 19790 24452 19796
rect 22468 18420 22520 18426
rect 22468 18362 22520 18368
rect 24124 18420 24176 18426
rect 24124 18362 24176 18368
rect 23480 18148 23532 18154
rect 23480 18090 23532 18096
rect 23492 16794 23520 18090
rect 23480 16788 23532 16794
rect 23480 16730 23532 16736
rect 24412 16454 24440 19790
rect 24676 19780 24728 19786
rect 24676 19722 24728 19728
rect 24688 16590 24716 19722
rect 26976 19168 27028 19174
rect 26976 19110 27028 19116
rect 26988 18290 27016 19110
rect 26976 18284 27028 18290
rect 26976 18226 27028 18232
rect 27540 17882 27568 21422
rect 28368 20058 28396 23054
rect 29656 21690 29684 25230
rect 29932 21690 29960 28970
rect 30392 28762 30420 29106
rect 32128 29096 32180 29102
rect 32128 29038 32180 29044
rect 30380 28756 30432 28762
rect 30380 28698 30432 28704
rect 32140 25498 32168 29038
rect 33520 26586 33548 31214
rect 34072 30938 34100 34546
rect 34164 34406 34192 34886
rect 34152 34400 34204 34406
rect 34152 34342 34204 34348
rect 34152 33312 34204 33318
rect 34152 33254 34204 33260
rect 34164 32858 34192 33254
rect 34256 32978 34284 38270
rect 34334 38200 34390 38270
rect 36004 38270 36138 38298
rect 34518 38176 34574 38185
rect 34518 38111 34574 38120
rect 34532 35222 34560 38111
rect 35530 36544 35586 36553
rect 34934 36476 35242 36485
rect 35530 36479 35586 36488
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35348 36236 35400 36242
rect 35348 36178 35400 36184
rect 35360 35894 35388 36178
rect 35544 36106 35572 36479
rect 35900 36168 35952 36174
rect 35900 36110 35952 36116
rect 35532 36100 35584 36106
rect 35532 36042 35584 36048
rect 35360 35866 35480 35894
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34520 35216 34572 35222
rect 34520 35158 34572 35164
rect 34520 35080 34572 35086
rect 34520 35022 34572 35028
rect 34796 35080 34848 35086
rect 34796 35022 34848 35028
rect 34532 34678 34560 35022
rect 34704 35012 34756 35018
rect 34704 34954 34756 34960
rect 34610 34912 34666 34921
rect 34610 34847 34666 34856
rect 34624 34746 34652 34847
rect 34612 34740 34664 34746
rect 34612 34682 34664 34688
rect 34520 34672 34572 34678
rect 34520 34614 34572 34620
rect 34336 34536 34388 34542
rect 34336 34478 34388 34484
rect 34520 34536 34572 34542
rect 34520 34478 34572 34484
rect 34244 32972 34296 32978
rect 34244 32914 34296 32920
rect 34164 32842 34284 32858
rect 34164 32836 34296 32842
rect 34164 32830 34244 32836
rect 34244 32778 34296 32784
rect 34256 32502 34284 32778
rect 34244 32496 34296 32502
rect 34244 32438 34296 32444
rect 34256 31686 34284 32438
rect 34348 32434 34376 34478
rect 34428 33856 34480 33862
rect 34428 33798 34480 33804
rect 34440 32586 34468 33798
rect 34532 32774 34560 34478
rect 34612 33992 34664 33998
rect 34612 33934 34664 33940
rect 34520 32768 34572 32774
rect 34520 32710 34572 32716
rect 34440 32558 34560 32586
rect 34336 32428 34388 32434
rect 34336 32370 34388 32376
rect 34244 31680 34296 31686
rect 34244 31622 34296 31628
rect 34060 30932 34112 30938
rect 34060 30874 34112 30880
rect 34532 30326 34560 32558
rect 34624 31890 34652 33934
rect 34716 33862 34744 34954
rect 34704 33856 34756 33862
rect 34704 33798 34756 33804
rect 34704 33312 34756 33318
rect 34704 33254 34756 33260
rect 34612 31884 34664 31890
rect 34612 31826 34664 31832
rect 34612 31680 34664 31686
rect 34612 31622 34664 31628
rect 34624 30682 34652 31622
rect 34716 30802 34744 33254
rect 34808 32026 34836 35022
rect 35348 34672 35400 34678
rect 35348 34614 35400 34620
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35256 34196 35308 34202
rect 35256 34138 35308 34144
rect 35268 33833 35296 34138
rect 35254 33824 35310 33833
rect 35254 33759 35310 33768
rect 35360 33522 35388 34614
rect 35452 34202 35480 35866
rect 35912 35766 35940 36110
rect 35900 35760 35952 35766
rect 35900 35702 35952 35708
rect 35624 35012 35676 35018
rect 35624 34954 35676 34960
rect 35440 34196 35492 34202
rect 35440 34138 35492 34144
rect 35532 33856 35584 33862
rect 35532 33798 35584 33804
rect 35544 33658 35572 33798
rect 35532 33652 35584 33658
rect 35532 33594 35584 33600
rect 35348 33516 35400 33522
rect 35348 33458 35400 33464
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34796 32020 34848 32026
rect 34796 31962 34848 31968
rect 35360 31890 35388 33458
rect 35532 32836 35584 32842
rect 35532 32778 35584 32784
rect 35440 32768 35492 32774
rect 35440 32710 35492 32716
rect 35452 32026 35480 32710
rect 35440 32020 35492 32026
rect 35440 31962 35492 31968
rect 35348 31884 35400 31890
rect 35348 31826 35400 31832
rect 34796 31816 34848 31822
rect 34796 31758 34848 31764
rect 34808 30870 34836 31758
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34796 30864 34848 30870
rect 34796 30806 34848 30812
rect 34704 30796 34756 30802
rect 34704 30738 34756 30744
rect 35256 30728 35308 30734
rect 34624 30666 34836 30682
rect 35256 30670 35308 30676
rect 34624 30660 34848 30666
rect 34624 30654 34796 30660
rect 34796 30602 34848 30608
rect 34520 30320 34572 30326
rect 34520 30262 34572 30268
rect 34704 30048 34756 30054
rect 34704 29990 34756 29996
rect 34716 29850 34744 29990
rect 34808 29850 34836 30602
rect 35268 30258 35296 30670
rect 35360 30258 35388 31826
rect 35544 31822 35572 32778
rect 35532 31816 35584 31822
rect 35532 31758 35584 31764
rect 35532 31680 35584 31686
rect 35532 31622 35584 31628
rect 35544 31346 35572 31622
rect 35440 31340 35492 31346
rect 35440 31282 35492 31288
rect 35532 31340 35584 31346
rect 35532 31282 35584 31288
rect 35452 31226 35480 31282
rect 35636 31226 35664 34954
rect 35716 34128 35768 34134
rect 35716 34070 35768 34076
rect 35728 33930 35756 34070
rect 35808 34060 35860 34066
rect 35808 34002 35860 34008
rect 35820 33946 35848 34002
rect 36004 33946 36032 38270
rect 36082 38200 36138 38270
rect 37830 38200 37886 39000
rect 36176 36032 36228 36038
rect 36176 35974 36228 35980
rect 36084 35012 36136 35018
rect 36084 34954 36136 34960
rect 35716 33924 35768 33930
rect 35820 33918 36032 33946
rect 35716 33866 35768 33872
rect 35714 33824 35770 33833
rect 35714 33759 35770 33768
rect 35728 33658 35756 33759
rect 35716 33652 35768 33658
rect 35716 33594 35768 33600
rect 35900 33652 35952 33658
rect 35900 33594 35952 33600
rect 35714 33280 35770 33289
rect 35714 33215 35770 33224
rect 35728 32366 35756 33215
rect 35808 32428 35860 32434
rect 35808 32370 35860 32376
rect 35716 32360 35768 32366
rect 35716 32302 35768 32308
rect 35820 31482 35848 32370
rect 35808 31476 35860 31482
rect 35808 31418 35860 31424
rect 35452 31198 35664 31226
rect 35532 30592 35584 30598
rect 35532 30534 35584 30540
rect 35544 30326 35572 30534
rect 35532 30320 35584 30326
rect 35532 30262 35584 30268
rect 35256 30252 35308 30258
rect 35256 30194 35308 30200
rect 35348 30252 35400 30258
rect 35348 30194 35400 30200
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34704 29844 34756 29850
rect 34704 29786 34756 29792
rect 34796 29844 34848 29850
rect 34796 29786 34848 29792
rect 34716 29306 34744 29786
rect 34704 29300 34756 29306
rect 34704 29242 34756 29248
rect 34808 29186 34836 29786
rect 34624 29170 34836 29186
rect 34612 29164 34836 29170
rect 34664 29158 34836 29164
rect 34612 29106 34664 29112
rect 34796 29028 34848 29034
rect 34796 28970 34848 28976
rect 34808 28082 34836 28970
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35360 28762 35388 30194
rect 35912 30138 35940 33594
rect 36096 33114 36124 34954
rect 36188 34513 36216 35974
rect 36636 35556 36688 35562
rect 36636 35498 36688 35504
rect 36360 35488 36412 35494
rect 36360 35430 36412 35436
rect 36544 35488 36596 35494
rect 36544 35430 36596 35436
rect 36268 35080 36320 35086
rect 36268 35022 36320 35028
rect 36174 34504 36230 34513
rect 36174 34439 36230 34448
rect 36176 34128 36228 34134
rect 36176 34070 36228 34076
rect 36188 33658 36216 34070
rect 36280 33862 36308 35022
rect 36372 34134 36400 35430
rect 36556 35290 36584 35430
rect 36544 35284 36596 35290
rect 36544 35226 36596 35232
rect 36452 35216 36504 35222
rect 36452 35158 36504 35164
rect 36360 34128 36412 34134
rect 36360 34070 36412 34076
rect 36268 33856 36320 33862
rect 36268 33798 36320 33804
rect 36176 33652 36228 33658
rect 36176 33594 36228 33600
rect 36084 33108 36136 33114
rect 36084 33050 36136 33056
rect 36360 33108 36412 33114
rect 36360 33050 36412 33056
rect 36082 33008 36138 33017
rect 36082 32943 36138 32952
rect 36096 32502 36124 32943
rect 36176 32904 36228 32910
rect 36176 32846 36228 32852
rect 36268 32904 36320 32910
rect 36268 32846 36320 32852
rect 36084 32496 36136 32502
rect 36084 32438 36136 32444
rect 36188 32026 36216 32846
rect 36176 32020 36228 32026
rect 36176 31962 36228 31968
rect 36280 31414 36308 32846
rect 36372 32502 36400 33050
rect 36360 32496 36412 32502
rect 36360 32438 36412 32444
rect 36268 31408 36320 31414
rect 36268 31350 36320 31356
rect 36464 31142 36492 35158
rect 36544 33924 36596 33930
rect 36544 33866 36596 33872
rect 36556 32570 36584 33866
rect 36544 32564 36596 32570
rect 36544 32506 36596 32512
rect 36648 32298 36676 35498
rect 36912 34944 36964 34950
rect 36912 34886 36964 34892
rect 36728 34604 36780 34610
rect 36728 34546 36780 34552
rect 36636 32292 36688 32298
rect 36636 32234 36688 32240
rect 36740 31958 36768 34546
rect 36924 33590 36952 34886
rect 36912 33584 36964 33590
rect 36912 33526 36964 33532
rect 37188 32836 37240 32842
rect 37188 32778 37240 32784
rect 36820 32496 36872 32502
rect 36820 32438 36872 32444
rect 36728 31952 36780 31958
rect 36728 31894 36780 31900
rect 36832 31890 36860 32438
rect 37004 31952 37056 31958
rect 37004 31894 37056 31900
rect 36820 31884 36872 31890
rect 36820 31826 36872 31832
rect 36832 31482 36860 31826
rect 36820 31476 36872 31482
rect 36820 31418 36872 31424
rect 37016 31278 37044 31894
rect 37200 31657 37228 32778
rect 37186 31648 37242 31657
rect 37186 31583 37242 31592
rect 37004 31272 37056 31278
rect 37004 31214 37056 31220
rect 37844 31210 37872 38200
rect 37832 31204 37884 31210
rect 37832 31146 37884 31152
rect 36452 31136 36504 31142
rect 36452 31078 36504 31084
rect 35992 30728 36044 30734
rect 35992 30670 36044 30676
rect 36268 30728 36320 30734
rect 36268 30670 36320 30676
rect 36004 30394 36032 30670
rect 35992 30388 36044 30394
rect 35992 30330 36044 30336
rect 35820 30110 35940 30138
rect 35716 29844 35768 29850
rect 35716 29786 35768 29792
rect 35532 28960 35584 28966
rect 35532 28902 35584 28908
rect 35348 28756 35400 28762
rect 35348 28698 35400 28704
rect 35164 28552 35216 28558
rect 35164 28494 35216 28500
rect 34796 28076 34848 28082
rect 34796 28018 34848 28024
rect 35176 28014 35204 28494
rect 35164 28008 35216 28014
rect 35164 27950 35216 27956
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34520 27532 34572 27538
rect 34520 27474 34572 27480
rect 33508 26580 33560 26586
rect 33508 26522 33560 26528
rect 34532 26246 34560 27474
rect 35360 26994 35388 28698
rect 35544 28558 35572 28902
rect 35532 28552 35584 28558
rect 35532 28494 35584 28500
rect 35532 28416 35584 28422
rect 35532 28358 35584 28364
rect 35544 28218 35572 28358
rect 35532 28212 35584 28218
rect 35532 28154 35584 28160
rect 35440 28008 35492 28014
rect 35440 27950 35492 27956
rect 35452 27606 35480 27950
rect 35440 27600 35492 27606
rect 35440 27542 35492 27548
rect 35532 27396 35584 27402
rect 35532 27338 35584 27344
rect 35440 27328 35492 27334
rect 35440 27270 35492 27276
rect 35452 27130 35480 27270
rect 35544 27130 35572 27338
rect 35440 27124 35492 27130
rect 35440 27066 35492 27072
rect 35532 27124 35584 27130
rect 35532 27066 35584 27072
rect 35348 26988 35400 26994
rect 35348 26930 35400 26936
rect 34704 26784 34756 26790
rect 34704 26726 34756 26732
rect 34716 26450 34744 26726
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34704 26444 34756 26450
rect 34704 26386 34756 26392
rect 34520 26240 34572 26246
rect 34520 26182 34572 26188
rect 34532 25838 34560 26182
rect 34520 25832 34572 25838
rect 34520 25774 34572 25780
rect 32128 25492 32180 25498
rect 32128 25434 32180 25440
rect 34532 24138 34560 25774
rect 34716 25770 34744 26386
rect 35360 26234 35388 26930
rect 35360 26206 35480 26234
rect 34704 25764 34756 25770
rect 34704 25706 34756 25712
rect 34796 25764 34848 25770
rect 34796 25706 34848 25712
rect 34808 24818 34836 25706
rect 35348 25696 35400 25702
rect 35348 25638 35400 25644
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 35360 25498 35388 25638
rect 35348 25492 35400 25498
rect 35348 25434 35400 25440
rect 35452 25294 35480 26206
rect 35624 25832 35676 25838
rect 35624 25774 35676 25780
rect 35636 25498 35664 25774
rect 35624 25492 35676 25498
rect 35624 25434 35676 25440
rect 35164 25288 35216 25294
rect 35164 25230 35216 25236
rect 35440 25288 35492 25294
rect 35440 25230 35492 25236
rect 35176 24954 35204 25230
rect 35348 25152 35400 25158
rect 35348 25094 35400 25100
rect 35164 24948 35216 24954
rect 35164 24890 35216 24896
rect 35360 24818 35388 25094
rect 34796 24812 34848 24818
rect 34796 24754 34848 24760
rect 35348 24812 35400 24818
rect 35348 24754 35400 24760
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34520 24132 34572 24138
rect 34520 24074 34572 24080
rect 35256 24064 35308 24070
rect 35256 24006 35308 24012
rect 35348 24064 35400 24070
rect 35348 24006 35400 24012
rect 35268 23866 35296 24006
rect 35256 23860 35308 23866
rect 35256 23802 35308 23808
rect 35360 23798 35388 24006
rect 35348 23792 35400 23798
rect 35348 23734 35400 23740
rect 35452 23662 35480 25230
rect 35532 24948 35584 24954
rect 35532 24890 35584 24896
rect 35544 24342 35572 24890
rect 35532 24336 35584 24342
rect 35532 24278 35584 24284
rect 35440 23656 35492 23662
rect 35440 23598 35492 23604
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 29644 21684 29696 21690
rect 29644 21626 29696 21632
rect 29920 21684 29972 21690
rect 29920 21626 29972 21632
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 35452 21010 35480 23598
rect 35624 23520 35676 23526
rect 35624 23462 35676 23468
rect 35636 23118 35664 23462
rect 35624 23112 35676 23118
rect 35624 23054 35676 23060
rect 35636 22166 35664 23054
rect 35624 22160 35676 22166
rect 35624 22102 35676 22108
rect 35532 21888 35584 21894
rect 35532 21830 35584 21836
rect 35440 21004 35492 21010
rect 35440 20946 35492 20952
rect 35544 20942 35572 21830
rect 35532 20936 35584 20942
rect 35532 20878 35584 20884
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35728 20058 35756 29786
rect 35820 27538 35848 30110
rect 36280 29714 36308 30670
rect 37188 30660 37240 30666
rect 37188 30602 37240 30608
rect 37200 30025 37228 30602
rect 37186 30016 37242 30025
rect 37186 29951 37242 29960
rect 36268 29708 36320 29714
rect 36268 29650 36320 29656
rect 36084 29164 36136 29170
rect 36084 29106 36136 29112
rect 36096 28150 36124 29106
rect 36912 29096 36964 29102
rect 36912 29038 36964 29044
rect 36820 29028 36872 29034
rect 36820 28970 36872 28976
rect 36832 28762 36860 28970
rect 36820 28756 36872 28762
rect 36820 28698 36872 28704
rect 36924 28393 36952 29038
rect 36910 28384 36966 28393
rect 36910 28319 36966 28328
rect 36084 28144 36136 28150
rect 36084 28086 36136 28092
rect 35808 27532 35860 27538
rect 35808 27474 35860 27480
rect 35992 27464 36044 27470
rect 35992 27406 36044 27412
rect 36268 27464 36320 27470
rect 36268 27406 36320 27412
rect 36004 27130 36032 27406
rect 35992 27124 36044 27130
rect 35992 27066 36044 27072
rect 36280 26586 36308 27406
rect 37280 27396 37332 27402
rect 37280 27338 37332 27344
rect 37292 26761 37320 27338
rect 37278 26752 37334 26761
rect 37278 26687 37334 26696
rect 36268 26580 36320 26586
rect 36268 26522 36320 26528
rect 35900 25900 35952 25906
rect 35900 25842 35952 25848
rect 35912 24886 35940 25842
rect 37464 25832 37516 25838
rect 37464 25774 37516 25780
rect 37476 25129 37504 25774
rect 37462 25120 37518 25129
rect 37462 25055 37518 25064
rect 35900 24880 35952 24886
rect 35900 24822 35952 24828
rect 35992 24200 36044 24206
rect 35992 24142 36044 24148
rect 36268 24200 36320 24206
rect 36268 24142 36320 24148
rect 36004 23866 36032 24142
rect 36084 24132 36136 24138
rect 36084 24074 36136 24080
rect 35992 23860 36044 23866
rect 35992 23802 36044 23808
rect 36096 22778 36124 24074
rect 36280 23186 36308 24142
rect 37280 24132 37332 24138
rect 37280 24074 37332 24080
rect 37292 23497 37320 24074
rect 37278 23488 37334 23497
rect 37278 23423 37334 23432
rect 36268 23180 36320 23186
rect 36268 23122 36320 23128
rect 36084 22772 36136 22778
rect 36084 22714 36136 22720
rect 36096 22098 36124 22714
rect 36452 22568 36504 22574
rect 36452 22510 36504 22516
rect 36084 22092 36136 22098
rect 36084 22034 36136 22040
rect 36096 20482 36124 22034
rect 36464 20874 36492 22510
rect 37096 22432 37148 22438
rect 37096 22374 37148 22380
rect 36544 21956 36596 21962
rect 36544 21898 36596 21904
rect 36556 21690 36584 21898
rect 36544 21684 36596 21690
rect 36544 21626 36596 21632
rect 36452 20868 36504 20874
rect 36452 20810 36504 20816
rect 36004 20454 36124 20482
rect 36004 20330 36032 20454
rect 37108 20398 37136 22374
rect 37462 21856 37518 21865
rect 37462 21791 37518 21800
rect 37476 21622 37504 21791
rect 37464 21616 37516 21622
rect 37464 21558 37516 21564
rect 36084 20392 36136 20398
rect 36084 20334 36136 20340
rect 37096 20392 37148 20398
rect 37096 20334 37148 20340
rect 35992 20324 36044 20330
rect 35992 20266 36044 20272
rect 28356 20052 28408 20058
rect 28356 19994 28408 20000
rect 35716 20052 35768 20058
rect 35716 19994 35768 20000
rect 36004 19922 36032 20266
rect 36096 19922 36124 20334
rect 35992 19916 36044 19922
rect 35992 19858 36044 19864
rect 36084 19916 36136 19922
rect 36084 19858 36136 19864
rect 34612 19848 34664 19854
rect 34612 19790 34664 19796
rect 34624 18358 34652 19790
rect 34796 19304 34848 19310
rect 34796 19246 34848 19252
rect 34704 18624 34756 18630
rect 34704 18566 34756 18572
rect 34716 18426 34744 18566
rect 34808 18426 34836 19246
rect 35624 19168 35676 19174
rect 35624 19110 35676 19116
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35348 18760 35400 18766
rect 35348 18702 35400 18708
rect 34704 18420 34756 18426
rect 34704 18362 34756 18368
rect 34796 18420 34848 18426
rect 34796 18362 34848 18368
rect 34612 18352 34664 18358
rect 34612 18294 34664 18300
rect 27528 17876 27580 17882
rect 27528 17818 27580 17824
rect 27896 17808 27948 17814
rect 27896 17750 27948 17756
rect 24676 16584 24728 16590
rect 24676 16526 24728 16532
rect 22284 16448 22336 16454
rect 22284 16390 22336 16396
rect 24400 16448 24452 16454
rect 24400 16390 24452 16396
rect 22296 16250 22324 16390
rect 22284 16244 22336 16250
rect 22284 16186 22336 16192
rect 24412 15910 24440 16390
rect 25320 15972 25372 15978
rect 25320 15914 25372 15920
rect 23204 15904 23256 15910
rect 23204 15846 23256 15852
rect 24400 15904 24452 15910
rect 24400 15846 24452 15852
rect 22008 15496 22060 15502
rect 22008 15438 22060 15444
rect 22928 15496 22980 15502
rect 22928 15438 22980 15444
rect 22940 10266 22968 15438
rect 23216 13394 23244 15846
rect 23388 15360 23440 15366
rect 23388 15302 23440 15308
rect 23204 13388 23256 13394
rect 23204 13330 23256 13336
rect 22928 10260 22980 10266
rect 22928 10202 22980 10208
rect 23400 3058 23428 15302
rect 23756 13184 23808 13190
rect 23756 13126 23808 13132
rect 23768 10130 23796 13126
rect 23756 10124 23808 10130
rect 23756 10066 23808 10072
rect 24412 7206 24440 15846
rect 24860 15632 24912 15638
rect 24860 15574 24912 15580
rect 24872 13326 24900 15574
rect 25332 13938 25360 15914
rect 25320 13932 25372 13938
rect 25320 13874 25372 13880
rect 24860 13320 24912 13326
rect 24860 13262 24912 13268
rect 25964 13184 26016 13190
rect 25964 13126 26016 13132
rect 24400 7200 24452 7206
rect 24400 7142 24452 7148
rect 25976 5234 26004 13126
rect 27908 10674 27936 17750
rect 30196 17536 30248 17542
rect 30196 17478 30248 17484
rect 34520 17536 34572 17542
rect 34520 17478 34572 17484
rect 29460 13864 29512 13870
rect 29460 13806 29512 13812
rect 28908 13320 28960 13326
rect 28908 13262 28960 13268
rect 28920 10810 28948 13262
rect 28908 10804 28960 10810
rect 28908 10746 28960 10752
rect 29472 10674 29500 13806
rect 27896 10668 27948 10674
rect 27896 10610 27948 10616
rect 28540 10668 28592 10674
rect 28540 10610 28592 10616
rect 29460 10668 29512 10674
rect 29460 10610 29512 10616
rect 27344 10464 27396 10470
rect 27344 10406 27396 10412
rect 25964 5228 26016 5234
rect 25964 5170 26016 5176
rect 27160 5160 27212 5166
rect 27160 5102 27212 5108
rect 26240 5024 26292 5030
rect 26240 4966 26292 4972
rect 26148 4752 26200 4758
rect 26148 4694 26200 4700
rect 25320 4072 25372 4078
rect 25320 4014 25372 4020
rect 24860 3936 24912 3942
rect 24860 3878 24912 3884
rect 24872 3466 24900 3878
rect 24860 3460 24912 3466
rect 24860 3402 24912 3408
rect 22192 3052 22244 3058
rect 22192 2994 22244 3000
rect 23388 3052 23440 3058
rect 23388 2994 23440 3000
rect 22204 2514 22232 2994
rect 23940 2984 23992 2990
rect 23940 2926 23992 2932
rect 22192 2508 22244 2514
rect 22192 2450 22244 2456
rect 22836 2508 22888 2514
rect 22836 2450 22888 2456
rect 21640 1352 21692 1358
rect 21640 1294 21692 1300
rect 22388 870 22508 898
rect 22388 800 22416 870
rect 19536 734 19932 762
rect 20902 0 20958 800
rect 22374 0 22430 800
rect 22480 762 22508 870
rect 22848 762 22876 2450
rect 23952 2446 23980 2926
rect 23940 2440 23992 2446
rect 23940 2382 23992 2388
rect 24124 2372 24176 2378
rect 24044 2332 24124 2360
rect 24044 1170 24072 2332
rect 24124 2314 24176 2320
rect 23860 1142 24072 1170
rect 23860 800 23888 1142
rect 25332 800 25360 4014
rect 26160 2650 26188 4694
rect 26252 4486 26280 4966
rect 26332 4616 26384 4622
rect 26332 4558 26384 4564
rect 26240 4480 26292 4486
rect 26240 4422 26292 4428
rect 26252 4214 26280 4422
rect 26240 4208 26292 4214
rect 26240 4150 26292 4156
rect 26252 3194 26280 4150
rect 26344 3738 26372 4558
rect 26700 4480 26752 4486
rect 26700 4422 26752 4428
rect 27068 4480 27120 4486
rect 27068 4422 27120 4428
rect 26332 3732 26384 3738
rect 26332 3674 26384 3680
rect 26240 3188 26292 3194
rect 26240 3130 26292 3136
rect 26148 2644 26200 2650
rect 26148 2586 26200 2592
rect 26712 2446 26740 4422
rect 26976 4276 27028 4282
rect 26976 4218 27028 4224
rect 26988 4146 27016 4218
rect 26976 4140 27028 4146
rect 26976 4082 27028 4088
rect 26884 3936 26936 3942
rect 26884 3878 26936 3884
rect 26896 3534 26924 3878
rect 26988 3738 27016 4082
rect 26976 3732 27028 3738
rect 26976 3674 27028 3680
rect 27080 3534 27108 4422
rect 26884 3528 26936 3534
rect 26884 3470 26936 3476
rect 27068 3528 27120 3534
rect 27068 3470 27120 3476
rect 26792 3460 26844 3466
rect 26792 3402 26844 3408
rect 26804 3194 26832 3402
rect 27172 3194 27200 5102
rect 26792 3188 26844 3194
rect 26792 3130 26844 3136
rect 27160 3188 27212 3194
rect 27160 3130 27212 3136
rect 27356 3058 27384 10406
rect 28172 5160 28224 5166
rect 28172 5102 28224 5108
rect 27804 5024 27856 5030
rect 27804 4966 27856 4972
rect 27712 4684 27764 4690
rect 27712 4626 27764 4632
rect 27528 4072 27580 4078
rect 27528 4014 27580 4020
rect 27540 3602 27568 4014
rect 27528 3596 27580 3602
rect 27528 3538 27580 3544
rect 27724 3126 27752 4626
rect 27712 3120 27764 3126
rect 27712 3062 27764 3068
rect 27344 3052 27396 3058
rect 27344 2994 27396 3000
rect 26976 2984 27028 2990
rect 26976 2926 27028 2932
rect 26988 2446 27016 2926
rect 27816 2446 27844 4966
rect 28184 2854 28212 5102
rect 28448 4480 28500 4486
rect 28448 4422 28500 4428
rect 28460 3058 28488 4422
rect 28448 3052 28500 3058
rect 28448 2994 28500 3000
rect 28172 2848 28224 2854
rect 28172 2790 28224 2796
rect 28552 2650 28580 10610
rect 29552 7200 29604 7206
rect 29552 7142 29604 7148
rect 29564 5574 29592 7142
rect 30208 5914 30236 17478
rect 34532 17338 34560 17478
rect 34520 17332 34572 17338
rect 34520 17274 34572 17280
rect 34624 16794 34652 18294
rect 34808 18222 34836 18362
rect 34796 18216 34848 18222
rect 34796 18158 34848 18164
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35360 17678 35388 18702
rect 35636 18290 35664 19110
rect 36004 18426 36032 19858
rect 36084 19372 36136 19378
rect 36084 19314 36136 19320
rect 35992 18420 36044 18426
rect 35992 18362 36044 18368
rect 36096 18358 36124 19314
rect 36912 19304 36964 19310
rect 36912 19246 36964 19252
rect 36924 18601 36952 19246
rect 37108 18902 37136 20334
rect 37278 20224 37334 20233
rect 37278 20159 37334 20168
rect 37292 19922 37320 20159
rect 37280 19916 37332 19922
rect 37280 19858 37332 19864
rect 37096 18896 37148 18902
rect 37096 18838 37148 18844
rect 37004 18692 37056 18698
rect 37004 18634 37056 18640
rect 36910 18592 36966 18601
rect 36910 18527 36966 18536
rect 37016 18426 37044 18634
rect 37004 18420 37056 18426
rect 37004 18362 37056 18368
rect 36084 18352 36136 18358
rect 36084 18294 36136 18300
rect 35624 18284 35676 18290
rect 35624 18226 35676 18232
rect 35532 18080 35584 18086
rect 35532 18022 35584 18028
rect 35544 17678 35572 18022
rect 35256 17672 35308 17678
rect 35256 17614 35308 17620
rect 35348 17672 35400 17678
rect 35348 17614 35400 17620
rect 35532 17672 35584 17678
rect 35532 17614 35584 17620
rect 34704 17536 34756 17542
rect 34704 17478 34756 17484
rect 34612 16788 34664 16794
rect 34612 16730 34664 16736
rect 34624 16574 34652 16730
rect 34716 16726 34744 17478
rect 35268 17338 35296 17614
rect 35256 17332 35308 17338
rect 35256 17274 35308 17280
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34704 16720 34756 16726
rect 34704 16662 34756 16668
rect 34532 16546 34652 16574
rect 34532 15366 34560 16546
rect 35360 16114 35388 17614
rect 36820 17536 36872 17542
rect 36820 17478 36872 17484
rect 36832 17338 36860 17478
rect 36820 17332 36872 17338
rect 36820 17274 36872 17280
rect 36268 17128 36320 17134
rect 36268 17070 36320 17076
rect 36280 16590 36308 17070
rect 37186 16960 37242 16969
rect 37186 16895 37242 16904
rect 37200 16658 37228 16895
rect 37188 16652 37240 16658
rect 37188 16594 37240 16600
rect 35992 16584 36044 16590
rect 35992 16526 36044 16532
rect 36268 16584 36320 16590
rect 36268 16526 36320 16532
rect 35440 16448 35492 16454
rect 35440 16390 35492 16396
rect 35532 16448 35584 16454
rect 35532 16390 35584 16396
rect 35452 16250 35480 16390
rect 35440 16244 35492 16250
rect 35440 16186 35492 16192
rect 35544 16182 35572 16390
rect 36004 16250 36032 16526
rect 35992 16244 36044 16250
rect 35992 16186 36044 16192
rect 35532 16176 35584 16182
rect 35532 16118 35584 16124
rect 35348 16108 35400 16114
rect 35348 16050 35400 16056
rect 34704 15904 34756 15910
rect 34704 15846 34756 15852
rect 34716 15570 34744 15846
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34704 15564 34756 15570
rect 34704 15506 34756 15512
rect 34520 15360 34572 15366
rect 34520 15302 34572 15308
rect 34532 15178 34560 15302
rect 34440 15150 34560 15178
rect 34440 14958 34468 15150
rect 34428 14952 34480 14958
rect 34428 14894 34480 14900
rect 34440 13172 34468 14894
rect 34716 14890 34744 15506
rect 34704 14884 34756 14890
rect 34704 14826 34756 14832
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35360 14482 35388 16050
rect 36544 15428 36596 15434
rect 36544 15370 36596 15376
rect 36556 15026 36584 15370
rect 36910 15328 36966 15337
rect 36910 15263 36966 15272
rect 36924 15094 36952 15263
rect 36912 15088 36964 15094
rect 36912 15030 36964 15036
rect 36544 15020 36596 15026
rect 36544 14962 36596 14968
rect 35440 14952 35492 14958
rect 35440 14894 35492 14900
rect 35452 14618 35480 14894
rect 35532 14816 35584 14822
rect 35532 14758 35584 14764
rect 35716 14816 35768 14822
rect 35716 14758 35768 14764
rect 35440 14612 35492 14618
rect 35440 14554 35492 14560
rect 35348 14476 35400 14482
rect 35348 14418 35400 14424
rect 34796 14408 34848 14414
rect 34796 14350 34848 14356
rect 34808 14074 34836 14350
rect 34796 14068 34848 14074
rect 34796 14010 34848 14016
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34520 13184 34572 13190
rect 34440 13144 34520 13172
rect 34520 13126 34572 13132
rect 34532 12102 34560 13126
rect 35360 12850 35388 14418
rect 35452 13462 35480 14554
rect 35544 14414 35572 14758
rect 35532 14408 35584 14414
rect 35532 14350 35584 14356
rect 35728 13938 35756 14758
rect 35808 14272 35860 14278
rect 35808 14214 35860 14220
rect 35820 14074 35848 14214
rect 35808 14068 35860 14074
rect 35808 14010 35860 14016
rect 35716 13932 35768 13938
rect 35716 13874 35768 13880
rect 36268 13864 36320 13870
rect 36268 13806 36320 13812
rect 35440 13456 35492 13462
rect 35440 13398 35492 13404
rect 36280 13326 36308 13806
rect 37278 13696 37334 13705
rect 37278 13631 37334 13640
rect 37292 13394 37320 13631
rect 37280 13388 37332 13394
rect 37280 13330 37332 13336
rect 35992 13320 36044 13326
rect 35992 13262 36044 13268
rect 36268 13320 36320 13326
rect 36268 13262 36320 13268
rect 35532 13252 35584 13258
rect 35532 13194 35584 13200
rect 35440 13184 35492 13190
rect 35440 13126 35492 13132
rect 35452 12986 35480 13126
rect 35544 12986 35572 13194
rect 36004 12986 36032 13262
rect 35440 12980 35492 12986
rect 35440 12922 35492 12928
rect 35532 12980 35584 12986
rect 35532 12922 35584 12928
rect 35992 12980 36044 12986
rect 35992 12922 36044 12928
rect 35348 12844 35400 12850
rect 35348 12786 35400 12792
rect 34704 12640 34756 12646
rect 34704 12582 34756 12588
rect 34716 12306 34744 12582
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34704 12300 34756 12306
rect 34704 12242 34756 12248
rect 34520 12096 34572 12102
rect 34520 12038 34572 12044
rect 34532 11694 34560 12038
rect 34520 11688 34572 11694
rect 34520 11630 34572 11636
rect 34532 9994 34560 11630
rect 34716 11626 34744 12242
rect 34704 11620 34756 11626
rect 34704 11562 34756 11568
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35360 11218 35388 12786
rect 36544 12164 36596 12170
rect 36544 12106 36596 12112
rect 36556 11898 36584 12106
rect 37462 12064 37518 12073
rect 37462 11999 37518 12008
rect 36544 11892 36596 11898
rect 36544 11834 36596 11840
rect 37476 11830 37504 11999
rect 37464 11824 37516 11830
rect 37464 11766 37516 11772
rect 35440 11688 35492 11694
rect 35440 11630 35492 11636
rect 35452 11354 35480 11630
rect 35532 11552 35584 11558
rect 35532 11494 35584 11500
rect 35624 11552 35676 11558
rect 35624 11494 35676 11500
rect 35440 11348 35492 11354
rect 35440 11290 35492 11296
rect 35348 11212 35400 11218
rect 35348 11154 35400 11160
rect 34796 11144 34848 11150
rect 34796 11086 34848 11092
rect 34808 10810 34836 11086
rect 34796 10804 34848 10810
rect 34796 10746 34848 10752
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35360 10062 35388 11154
rect 35452 10198 35480 11290
rect 35544 11150 35572 11494
rect 35532 11144 35584 11150
rect 35532 11086 35584 11092
rect 35636 10674 35664 11494
rect 36820 11008 36872 11014
rect 36820 10950 36872 10956
rect 36832 10674 36860 10950
rect 35624 10668 35676 10674
rect 35624 10610 35676 10616
rect 36820 10668 36872 10674
rect 36820 10610 36872 10616
rect 36084 10600 36136 10606
rect 36084 10542 36136 10548
rect 35440 10192 35492 10198
rect 35440 10134 35492 10140
rect 36096 10130 36124 10542
rect 37278 10432 37334 10441
rect 37278 10367 37334 10376
rect 37292 10130 37320 10367
rect 35532 10124 35584 10130
rect 35532 10066 35584 10072
rect 36084 10124 36136 10130
rect 36084 10066 36136 10072
rect 37280 10124 37332 10130
rect 37280 10066 37332 10072
rect 35348 10056 35400 10062
rect 35348 9998 35400 10004
rect 34520 9988 34572 9994
rect 34520 9930 34572 9936
rect 31024 9920 31076 9926
rect 31024 9862 31076 9868
rect 31036 7478 31064 9862
rect 35360 9586 35388 9998
rect 35440 9920 35492 9926
rect 35440 9862 35492 9868
rect 35452 9722 35480 9862
rect 35440 9716 35492 9722
rect 35440 9658 35492 9664
rect 35544 9654 35572 10066
rect 35992 10056 36044 10062
rect 35992 9998 36044 10004
rect 35808 9988 35860 9994
rect 35808 9930 35860 9936
rect 35532 9648 35584 9654
rect 35532 9590 35584 9596
rect 35348 9580 35400 9586
rect 35348 9522 35400 9528
rect 34704 9376 34756 9382
rect 34704 9318 34756 9324
rect 34716 9178 34744 9318
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34704 9172 34756 9178
rect 34704 9114 34756 9120
rect 34520 8832 34572 8838
rect 34520 8774 34572 8780
rect 34532 8430 34560 8774
rect 34716 8634 34744 9114
rect 34704 8628 34756 8634
rect 34704 8570 34756 8576
rect 34520 8424 34572 8430
rect 34520 8366 34572 8372
rect 33692 7744 33744 7750
rect 33692 7686 33744 7692
rect 31024 7472 31076 7478
rect 31024 7414 31076 7420
rect 33508 7336 33560 7342
rect 33508 7278 33560 7284
rect 32404 6656 32456 6662
rect 32404 6598 32456 6604
rect 33048 6656 33100 6662
rect 33048 6598 33100 6604
rect 30196 5908 30248 5914
rect 30196 5850 30248 5856
rect 29092 5568 29144 5574
rect 29092 5510 29144 5516
rect 29552 5568 29604 5574
rect 29552 5510 29604 5516
rect 28632 4616 28684 4622
rect 28632 4558 28684 4564
rect 28724 4616 28776 4622
rect 28724 4558 28776 4564
rect 28644 4282 28672 4558
rect 28632 4276 28684 4282
rect 28632 4218 28684 4224
rect 28736 4146 28764 4558
rect 28724 4140 28776 4146
rect 28724 4082 28776 4088
rect 28632 4072 28684 4078
rect 28632 4014 28684 4020
rect 28540 2644 28592 2650
rect 28540 2586 28592 2592
rect 26700 2440 26752 2446
rect 26700 2382 26752 2388
rect 26976 2440 27028 2446
rect 26976 2382 27028 2388
rect 27160 2440 27212 2446
rect 27160 2382 27212 2388
rect 27804 2440 27856 2446
rect 27804 2382 27856 2388
rect 26804 870 26924 898
rect 26804 800 26832 870
rect 22480 734 22876 762
rect 23846 0 23902 800
rect 25318 0 25374 800
rect 26790 0 26846 800
rect 26896 762 26924 870
rect 27172 762 27200 2382
rect 28276 870 28396 898
rect 28276 800 28304 870
rect 26896 734 27200 762
rect 28262 0 28318 800
rect 28368 762 28396 870
rect 28644 762 28672 4014
rect 28736 2650 28764 4082
rect 29104 3534 29132 5510
rect 30208 5166 30236 5850
rect 32416 5778 32444 6598
rect 32404 5772 32456 5778
rect 32404 5714 32456 5720
rect 31392 5636 31444 5642
rect 31392 5578 31444 5584
rect 31404 5234 31432 5578
rect 32220 5568 32272 5574
rect 32220 5510 32272 5516
rect 31392 5228 31444 5234
rect 31392 5170 31444 5176
rect 29460 5160 29512 5166
rect 29460 5102 29512 5108
rect 29552 5160 29604 5166
rect 29552 5102 29604 5108
rect 30196 5160 30248 5166
rect 30196 5102 30248 5108
rect 30656 5160 30708 5166
rect 30656 5102 30708 5108
rect 29368 5092 29420 5098
rect 29368 5034 29420 5040
rect 29092 3528 29144 3534
rect 29092 3470 29144 3476
rect 29380 3058 29408 5034
rect 29472 4826 29500 5102
rect 29460 4820 29512 4826
rect 29460 4762 29512 4768
rect 29460 4684 29512 4690
rect 29460 4626 29512 4632
rect 29472 3670 29500 4626
rect 29564 3738 29592 5102
rect 30208 4690 30236 5102
rect 30288 5024 30340 5030
rect 30288 4966 30340 4972
rect 30196 4684 30248 4690
rect 30196 4626 30248 4632
rect 30104 4480 30156 4486
rect 30104 4422 30156 4428
rect 29736 4072 29788 4078
rect 29736 4014 29788 4020
rect 29552 3732 29604 3738
rect 29552 3674 29604 3680
rect 29460 3664 29512 3670
rect 29460 3606 29512 3612
rect 29552 3528 29604 3534
rect 29552 3470 29604 3476
rect 29564 3194 29592 3470
rect 29552 3188 29604 3194
rect 29552 3130 29604 3136
rect 29368 3052 29420 3058
rect 29368 2994 29420 3000
rect 29092 2984 29144 2990
rect 29092 2926 29144 2932
rect 28724 2644 28776 2650
rect 28724 2586 28776 2592
rect 29104 2446 29132 2926
rect 29092 2440 29144 2446
rect 29092 2382 29144 2388
rect 29748 800 29776 4014
rect 30116 3466 30144 4422
rect 30104 3460 30156 3466
rect 30104 3402 30156 3408
rect 30300 2514 30328 4966
rect 30472 4140 30524 4146
rect 30472 4082 30524 4088
rect 30484 3194 30512 4082
rect 30668 4010 30696 5102
rect 31404 4758 31432 5170
rect 31852 5092 31904 5098
rect 31852 5034 31904 5040
rect 31760 5024 31812 5030
rect 31760 4966 31812 4972
rect 31392 4752 31444 4758
rect 31392 4694 31444 4700
rect 31116 4684 31168 4690
rect 31116 4626 31168 4632
rect 31128 4282 31156 4626
rect 31116 4276 31168 4282
rect 31116 4218 31168 4224
rect 30656 4004 30708 4010
rect 30656 3946 30708 3952
rect 30668 3777 30696 3946
rect 30654 3768 30710 3777
rect 30654 3703 30710 3712
rect 31392 3460 31444 3466
rect 31392 3402 31444 3408
rect 31024 3392 31076 3398
rect 31024 3334 31076 3340
rect 31036 3194 31064 3334
rect 30472 3188 30524 3194
rect 30472 3130 30524 3136
rect 31024 3188 31076 3194
rect 31024 3130 31076 3136
rect 31404 3126 31432 3402
rect 31392 3120 31444 3126
rect 31392 3062 31444 3068
rect 31208 2848 31260 2854
rect 31208 2790 31260 2796
rect 30288 2508 30340 2514
rect 30288 2450 30340 2456
rect 31220 800 31248 2790
rect 31772 2446 31800 4966
rect 31864 3126 31892 5034
rect 32232 5030 32260 5510
rect 32416 5098 32444 5714
rect 32772 5160 32824 5166
rect 32772 5102 32824 5108
rect 32404 5092 32456 5098
rect 32404 5034 32456 5040
rect 31944 5024 31996 5030
rect 31944 4966 31996 4972
rect 32220 5024 32272 5030
rect 32220 4966 32272 4972
rect 32680 5024 32732 5030
rect 32680 4966 32732 4972
rect 31852 3120 31904 3126
rect 31852 3062 31904 3068
rect 31864 2650 31892 3062
rect 31956 3058 31984 4966
rect 32496 4140 32548 4146
rect 32496 4082 32548 4088
rect 32128 4072 32180 4078
rect 32128 4014 32180 4020
rect 32140 3738 32168 4014
rect 32128 3732 32180 3738
rect 32128 3674 32180 3680
rect 31944 3052 31996 3058
rect 31944 2994 31996 3000
rect 31852 2644 31904 2650
rect 31852 2586 31904 2592
rect 32508 2514 32536 4082
rect 32692 3466 32720 4966
rect 32784 4214 32812 5102
rect 32772 4208 32824 4214
rect 33060 4185 33088 6598
rect 33520 6458 33548 7278
rect 33704 6866 33732 7686
rect 34336 7336 34388 7342
rect 34336 7278 34388 7284
rect 33968 7200 34020 7206
rect 33968 7142 34020 7148
rect 34244 7200 34296 7206
rect 34244 7142 34296 7148
rect 33692 6860 33744 6866
rect 33692 6802 33744 6808
rect 33508 6452 33560 6458
rect 33508 6394 33560 6400
rect 33876 6112 33928 6118
rect 33876 6054 33928 6060
rect 33888 5914 33916 6054
rect 33876 5908 33928 5914
rect 33876 5850 33928 5856
rect 33980 5710 34008 7142
rect 34256 6866 34284 7142
rect 34244 6860 34296 6866
rect 34244 6802 34296 6808
rect 34152 6656 34204 6662
rect 34152 6598 34204 6604
rect 34060 6316 34112 6322
rect 34060 6258 34112 6264
rect 33876 5704 33928 5710
rect 33876 5646 33928 5652
rect 33968 5704 34020 5710
rect 33968 5646 34020 5652
rect 33888 4826 33916 5646
rect 33876 4820 33928 4826
rect 33876 4762 33928 4768
rect 33876 4684 33928 4690
rect 33876 4626 33928 4632
rect 33508 4616 33560 4622
rect 33508 4558 33560 4564
rect 32772 4150 32824 4156
rect 33046 4176 33102 4185
rect 32784 3738 32812 4150
rect 33046 4111 33102 4120
rect 32772 3732 32824 3738
rect 32772 3674 32824 3680
rect 32680 3460 32732 3466
rect 32680 3402 32732 3408
rect 33060 2922 33088 4111
rect 33140 3936 33192 3942
rect 33140 3878 33192 3884
rect 33152 3346 33180 3878
rect 33152 3318 33272 3346
rect 33048 2916 33100 2922
rect 33048 2858 33100 2864
rect 32496 2508 32548 2514
rect 32496 2450 32548 2456
rect 33140 2508 33192 2514
rect 33140 2450 33192 2456
rect 31760 2440 31812 2446
rect 31760 2382 31812 2388
rect 33152 1442 33180 2450
rect 33244 2446 33272 3318
rect 33520 3126 33548 4558
rect 33692 4548 33744 4554
rect 33692 4490 33744 4496
rect 33598 3768 33654 3777
rect 33598 3703 33654 3712
rect 33508 3120 33560 3126
rect 33508 3062 33560 3068
rect 33612 2650 33640 3703
rect 33704 3398 33732 4490
rect 33692 3392 33744 3398
rect 33692 3334 33744 3340
rect 33888 3058 33916 4626
rect 33876 3052 33928 3058
rect 33876 2994 33928 3000
rect 33980 2938 34008 5646
rect 34072 4808 34100 6258
rect 34164 6254 34192 6598
rect 34152 6248 34204 6254
rect 34152 6190 34204 6196
rect 34164 5846 34192 6190
rect 34152 5840 34204 5846
rect 34152 5782 34204 5788
rect 34244 5772 34296 5778
rect 34244 5714 34296 5720
rect 34256 5302 34284 5714
rect 34244 5296 34296 5302
rect 34244 5238 34296 5244
rect 34072 4780 34192 4808
rect 34060 4684 34112 4690
rect 34060 4626 34112 4632
rect 34072 3074 34100 4626
rect 34164 4214 34192 4780
rect 34152 4208 34204 4214
rect 34152 4150 34204 4156
rect 34164 3534 34192 4150
rect 34244 4140 34296 4146
rect 34244 4082 34296 4088
rect 34152 3528 34204 3534
rect 34152 3470 34204 3476
rect 34256 3194 34284 4082
rect 34348 3738 34376 7278
rect 34532 6662 34560 8366
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35360 7954 35388 9522
rect 35440 8424 35492 8430
rect 35440 8366 35492 8372
rect 35452 8090 35480 8366
rect 35532 8288 35584 8294
rect 35532 8230 35584 8236
rect 35624 8288 35676 8294
rect 35624 8230 35676 8236
rect 35440 8084 35492 8090
rect 35440 8026 35492 8032
rect 35348 7948 35400 7954
rect 35348 7890 35400 7896
rect 34704 7880 34756 7886
rect 34704 7822 34756 7828
rect 34796 7880 34848 7886
rect 34796 7822 34848 7828
rect 34520 6656 34572 6662
rect 34520 6598 34572 6604
rect 34532 6254 34560 6598
rect 34716 6338 34744 7822
rect 34808 7546 34836 7822
rect 34796 7540 34848 7546
rect 34796 7482 34848 7488
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35256 6656 35308 6662
rect 35256 6598 35308 6604
rect 35268 6458 35296 6598
rect 35256 6452 35308 6458
rect 35256 6394 35308 6400
rect 34716 6310 34836 6338
rect 35360 6322 35388 7890
rect 35452 6934 35480 8026
rect 35544 7886 35572 8230
rect 35532 7880 35584 7886
rect 35532 7822 35584 7828
rect 35636 7410 35664 8230
rect 35624 7404 35676 7410
rect 35624 7346 35676 7352
rect 35440 6928 35492 6934
rect 35440 6870 35492 6876
rect 34520 6248 34572 6254
rect 34520 6190 34572 6196
rect 34704 6248 34756 6254
rect 34704 6190 34756 6196
rect 34428 5636 34480 5642
rect 34428 5578 34480 5584
rect 34440 4026 34468 5578
rect 34532 5302 34560 6190
rect 34612 5704 34664 5710
rect 34612 5646 34664 5652
rect 34624 5302 34652 5646
rect 34520 5296 34572 5302
rect 34520 5238 34572 5244
rect 34612 5296 34664 5302
rect 34612 5238 34664 5244
rect 34532 4486 34560 5238
rect 34520 4480 34572 4486
rect 34520 4422 34572 4428
rect 34532 4146 34560 4422
rect 34520 4140 34572 4146
rect 34520 4082 34572 4088
rect 34610 4040 34666 4049
rect 34440 3998 34610 4026
rect 34610 3975 34666 3984
rect 34428 3936 34480 3942
rect 34428 3878 34480 3884
rect 34612 3936 34664 3942
rect 34612 3878 34664 3884
rect 34336 3732 34388 3738
rect 34336 3674 34388 3680
rect 34440 3602 34468 3878
rect 34624 3738 34652 3878
rect 34520 3732 34572 3738
rect 34520 3674 34572 3680
rect 34612 3732 34664 3738
rect 34612 3674 34664 3680
rect 34428 3596 34480 3602
rect 34428 3538 34480 3544
rect 34244 3188 34296 3194
rect 34244 3130 34296 3136
rect 34072 3046 34376 3074
rect 33980 2922 34284 2938
rect 33980 2916 34296 2922
rect 33980 2910 34244 2916
rect 34244 2858 34296 2864
rect 34348 2774 34376 3046
rect 34440 2990 34468 3538
rect 34532 3398 34560 3674
rect 34520 3392 34572 3398
rect 34520 3334 34572 3340
rect 34428 2984 34480 2990
rect 34428 2926 34480 2932
rect 34164 2746 34376 2774
rect 33600 2644 33652 2650
rect 33600 2586 33652 2592
rect 33232 2440 33284 2446
rect 33232 2382 33284 2388
rect 33060 1414 33180 1442
rect 32692 870 32812 898
rect 32692 800 32720 870
rect 28368 734 28672 762
rect 29734 0 29790 800
rect 31206 0 31262 800
rect 32678 0 32734 800
rect 32784 762 32812 870
rect 33060 762 33088 1414
rect 34164 800 34192 2746
rect 34440 2582 34468 2926
rect 34532 2582 34560 3334
rect 34428 2576 34480 2582
rect 34428 2518 34480 2524
rect 34520 2576 34572 2582
rect 34520 2518 34572 2524
rect 34716 2446 34744 6190
rect 34808 5166 34836 6310
rect 35256 6316 35308 6322
rect 35256 6258 35308 6264
rect 35348 6316 35400 6322
rect 35348 6258 35400 6264
rect 35268 6066 35296 6258
rect 35268 6038 35480 6066
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34888 5568 34940 5574
rect 34888 5510 34940 5516
rect 34796 5160 34848 5166
rect 34796 5102 34848 5108
rect 34900 5012 34928 5510
rect 34808 4984 34928 5012
rect 34808 4808 34836 4984
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34808 4780 34928 4808
rect 34796 4616 34848 4622
rect 34796 4558 34848 4564
rect 34808 4214 34836 4558
rect 34796 4208 34848 4214
rect 34796 4150 34848 4156
rect 34900 4060 34928 4780
rect 35452 4146 35480 6038
rect 35716 5704 35768 5710
rect 35716 5646 35768 5652
rect 35624 5636 35676 5642
rect 35624 5578 35676 5584
rect 35440 4140 35492 4146
rect 35440 4082 35492 4088
rect 34808 4032 34928 4060
rect 34808 3398 34836 4032
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34796 3392 34848 3398
rect 34796 3334 34848 3340
rect 35636 3058 35664 5578
rect 35728 3670 35756 5646
rect 35820 4690 35848 9930
rect 36004 9722 36032 9998
rect 35992 9716 36044 9722
rect 35992 9658 36044 9664
rect 36544 8900 36596 8906
rect 36544 8842 36596 8848
rect 36556 8634 36584 8842
rect 37462 8800 37518 8809
rect 37462 8735 37518 8744
rect 36544 8628 36596 8634
rect 36544 8570 36596 8576
rect 37476 8566 37504 8735
rect 37464 8560 37516 8566
rect 37464 8502 37516 8508
rect 37280 7812 37332 7818
rect 37280 7754 37332 7760
rect 36820 7744 36872 7750
rect 36820 7686 36872 7692
rect 36912 7744 36964 7750
rect 36912 7686 36964 7692
rect 36832 7546 36860 7686
rect 36820 7540 36872 7546
rect 36820 7482 36872 7488
rect 36176 7336 36228 7342
rect 36176 7278 36228 7284
rect 36188 6798 36216 7278
rect 35992 6792 36044 6798
rect 35992 6734 36044 6740
rect 36176 6792 36228 6798
rect 36176 6734 36228 6740
rect 36004 6458 36032 6734
rect 35992 6452 36044 6458
rect 35992 6394 36044 6400
rect 36176 6112 36228 6118
rect 36176 6054 36228 6060
rect 35900 5636 35952 5642
rect 35900 5578 35952 5584
rect 35912 5370 35940 5578
rect 35900 5364 35952 5370
rect 35900 5306 35952 5312
rect 36084 5160 36136 5166
rect 36084 5102 36136 5108
rect 36096 4826 36124 5102
rect 36084 4820 36136 4826
rect 36084 4762 36136 4768
rect 35808 4684 35860 4690
rect 35808 4626 35860 4632
rect 35900 4140 35952 4146
rect 35900 4082 35952 4088
rect 35716 3664 35768 3670
rect 35716 3606 35768 3612
rect 35348 3052 35400 3058
rect 35348 2994 35400 3000
rect 35624 3052 35676 3058
rect 35624 2994 35676 3000
rect 35360 2774 35388 2994
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 35360 2746 35572 2774
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34704 2440 34756 2446
rect 34704 2382 34756 2388
rect 35544 2258 35572 2746
rect 35912 2650 35940 4082
rect 36188 3534 36216 6054
rect 36544 5636 36596 5642
rect 36544 5578 36596 5584
rect 36556 4622 36584 5578
rect 36544 4616 36596 4622
rect 36544 4558 36596 4564
rect 36634 4176 36690 4185
rect 36634 4111 36636 4120
rect 36688 4111 36690 4120
rect 36636 4082 36688 4088
rect 36924 3942 36952 7686
rect 37186 7168 37242 7177
rect 37186 7103 37242 7112
rect 37200 6866 37228 7103
rect 37188 6860 37240 6866
rect 37188 6802 37240 6808
rect 37096 5024 37148 5030
rect 37096 4966 37148 4972
rect 37108 4622 37136 4966
rect 37096 4616 37148 4622
rect 37096 4558 37148 4564
rect 37004 4276 37056 4282
rect 37004 4218 37056 4224
rect 36912 3936 36964 3942
rect 36912 3878 36964 3884
rect 36176 3528 36228 3534
rect 36176 3470 36228 3476
rect 36924 3466 36952 3878
rect 36268 3460 36320 3466
rect 36268 3402 36320 3408
rect 36912 3460 36964 3466
rect 36912 3402 36964 3408
rect 36280 3097 36308 3402
rect 36266 3088 36322 3097
rect 36266 3023 36322 3032
rect 35900 2644 35952 2650
rect 35900 2586 35952 2592
rect 35544 2230 35664 2258
rect 34520 1352 34572 1358
rect 34520 1294 34572 1300
rect 32784 734 33088 762
rect 34150 0 34206 800
rect 34532 649 34560 1294
rect 35636 800 35664 2230
rect 37016 2122 37044 4218
rect 37108 3738 37136 4558
rect 37096 3732 37148 3738
rect 37096 3674 37148 3680
rect 37292 2650 37320 7754
rect 37646 5536 37702 5545
rect 37646 5471 37702 5480
rect 37660 4690 37688 5471
rect 37648 4684 37700 4690
rect 37648 4626 37700 4632
rect 37280 2644 37332 2650
rect 37280 2586 37332 2592
rect 37924 2372 37976 2378
rect 37924 2314 37976 2320
rect 37936 2281 37964 2314
rect 37922 2272 37978 2281
rect 37922 2207 37978 2216
rect 37016 2094 37136 2122
rect 37108 800 37136 2094
rect 34518 640 34574 649
rect 34518 575 34574 584
rect 35622 0 35678 800
rect 37094 0 37150 800
<< via2 >>
rect 3330 36488 3386 36544
rect 1582 33224 1638 33280
rect 1582 31592 1638 31648
rect 1582 30232 1638 30288
rect 1582 28328 1638 28384
rect 1582 26968 1638 27024
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4066 34856 4122 34912
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 938 25064 994 25120
rect 938 23432 994 23488
rect 1582 21936 1638 21992
rect 938 20168 994 20224
rect 1582 18536 1638 18592
rect 1582 16632 1638 16688
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 1582 15272 1638 15328
rect 938 13640 994 13696
rect 938 12008 994 12064
rect 938 10376 994 10432
rect 938 8744 994 8800
rect 1582 6976 1638 7032
rect 938 5480 994 5536
rect 938 3848 994 3904
rect 1582 2624 1638 2680
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 30010 34448 30066 34504
rect 32034 34448 32090 34504
rect 31666 32952 31722 33008
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 20626 3068 20628 3088
rect 20628 3068 20680 3088
rect 20680 3068 20682 3088
rect 20626 3032 20682 3068
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34518 38120 34574 38176
rect 35530 36488 35586 36544
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34610 34856 34666 34912
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 35254 33768 35310 33824
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 35714 33768 35770 33824
rect 35714 33224 35770 33280
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 36174 34448 36230 34504
rect 36082 32952 36138 33008
rect 37186 31592 37242 31648
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 37186 29960 37242 30016
rect 36910 28328 36966 28384
rect 37278 26696 37334 26752
rect 37462 25064 37518 25120
rect 37278 23432 37334 23488
rect 37462 21800 37518 21856
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 37278 20168 37334 20224
rect 36910 18536 36966 18592
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 37186 16904 37242 16960
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 36910 15272 36966 15328
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 37278 13640 37334 13696
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 37462 12008 37518 12064
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 37278 10376 37334 10432
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 30654 3712 30710 3768
rect 33046 4120 33102 4176
rect 33598 3712 33654 3768
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34610 3984 34666 4040
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 37462 8744 37518 8800
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 36634 4140 36690 4176
rect 36634 4120 36636 4140
rect 36636 4120 36688 4140
rect 36688 4120 36690 4140
rect 37186 7112 37242 7168
rect 36266 3032 36322 3088
rect 37646 5480 37702 5536
rect 37922 2216 37978 2272
rect 34518 584 34574 640
<< metal3 >>
rect 34513 38178 34579 38181
rect 38200 38178 39000 38208
rect 34513 38176 39000 38178
rect 34513 38120 34518 38176
rect 34574 38120 39000 38176
rect 34513 38118 39000 38120
rect 34513 38115 34579 38118
rect 38200 38088 39000 38118
rect 0 36546 800 36576
rect 3325 36546 3391 36549
rect 0 36544 3391 36546
rect 0 36488 3330 36544
rect 3386 36488 3391 36544
rect 0 36486 3391 36488
rect 0 36456 800 36486
rect 3325 36483 3391 36486
rect 35525 36546 35591 36549
rect 38200 36546 39000 36576
rect 35525 36544 39000 36546
rect 35525 36488 35530 36544
rect 35586 36488 39000 36544
rect 35525 36486 39000 36488
rect 35525 36483 35591 36486
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 38200 36456 39000 36486
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 0 34914 800 34944
rect 4061 34914 4127 34917
rect 0 34912 4127 34914
rect 0 34856 4066 34912
rect 4122 34856 4127 34912
rect 0 34854 4127 34856
rect 0 34824 800 34854
rect 4061 34851 4127 34854
rect 34605 34914 34671 34917
rect 38200 34914 39000 34944
rect 34605 34912 39000 34914
rect 34605 34856 34610 34912
rect 34666 34856 39000 34912
rect 34605 34854 39000 34856
rect 34605 34851 34671 34854
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 38200 34824 39000 34854
rect 19570 34783 19886 34784
rect 30005 34506 30071 34509
rect 32029 34506 32095 34509
rect 36169 34506 36235 34509
rect 30005 34504 36235 34506
rect 30005 34448 30010 34504
rect 30066 34448 32034 34504
rect 32090 34448 36174 34504
rect 36230 34448 36235 34504
rect 30005 34446 36235 34448
rect 30005 34443 30071 34446
rect 32029 34443 32095 34446
rect 36169 34443 36235 34446
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 35249 33826 35315 33829
rect 35709 33826 35775 33829
rect 35249 33824 35775 33826
rect 35249 33768 35254 33824
rect 35310 33768 35714 33824
rect 35770 33768 35775 33824
rect 35249 33766 35775 33768
rect 35249 33763 35315 33766
rect 35709 33763 35775 33766
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 0 33282 800 33312
rect 1577 33282 1643 33285
rect 0 33280 1643 33282
rect 0 33224 1582 33280
rect 1638 33224 1643 33280
rect 0 33222 1643 33224
rect 0 33192 800 33222
rect 1577 33219 1643 33222
rect 35709 33282 35775 33285
rect 38200 33282 39000 33312
rect 35709 33280 39000 33282
rect 35709 33224 35714 33280
rect 35770 33224 39000 33280
rect 35709 33222 39000 33224
rect 35709 33219 35775 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 38200 33192 39000 33222
rect 34930 33151 35246 33152
rect 31661 33010 31727 33013
rect 36077 33010 36143 33013
rect 31661 33008 36143 33010
rect 31661 32952 31666 33008
rect 31722 32952 36082 33008
rect 36138 32952 36143 33008
rect 31661 32950 36143 32952
rect 31661 32947 31727 32950
rect 36077 32947 36143 32950
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 0 31650 800 31680
rect 1577 31650 1643 31653
rect 0 31648 1643 31650
rect 0 31592 1582 31648
rect 1638 31592 1643 31648
rect 0 31590 1643 31592
rect 0 31560 800 31590
rect 1577 31587 1643 31590
rect 37181 31650 37247 31653
rect 38200 31650 39000 31680
rect 37181 31648 39000 31650
rect 37181 31592 37186 31648
rect 37242 31592 39000 31648
rect 37181 31590 39000 31592
rect 37181 31587 37247 31590
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 38200 31560 39000 31590
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 1577 30290 1643 30293
rect 798 30288 1643 30290
rect 798 30232 1582 30288
rect 1638 30232 1643 30288
rect 798 30230 1643 30232
rect 798 30048 858 30230
rect 1577 30227 1643 30230
rect 0 29958 858 30048
rect 37181 30018 37247 30021
rect 38200 30018 39000 30048
rect 37181 30016 39000 30018
rect 37181 29960 37186 30016
rect 37242 29960 39000 30016
rect 37181 29958 39000 29960
rect 0 29928 800 29958
rect 37181 29955 37247 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 38200 29928 39000 29958
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 0 28386 800 28416
rect 1577 28386 1643 28389
rect 0 28384 1643 28386
rect 0 28328 1582 28384
rect 1638 28328 1643 28384
rect 0 28326 1643 28328
rect 0 28296 800 28326
rect 1577 28323 1643 28326
rect 36905 28386 36971 28389
rect 38200 28386 39000 28416
rect 36905 28384 39000 28386
rect 36905 28328 36910 28384
rect 36966 28328 39000 28384
rect 36905 28326 39000 28328
rect 36905 28323 36971 28326
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 38200 28296 39000 28326
rect 19570 28255 19886 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 1577 27026 1643 27029
rect 982 27024 1643 27026
rect 982 26968 1582 27024
rect 1638 26968 1643 27024
rect 982 26966 1643 26968
rect 0 26754 800 26784
rect 982 26754 1042 26966
rect 1577 26963 1643 26966
rect 0 26694 1042 26754
rect 37273 26754 37339 26757
rect 38200 26754 39000 26784
rect 37273 26752 39000 26754
rect 37273 26696 37278 26752
rect 37334 26696 39000 26752
rect 37273 26694 39000 26696
rect 0 26664 800 26694
rect 37273 26691 37339 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 38200 26664 39000 26694
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 0 25122 800 25152
rect 933 25122 999 25125
rect 0 25120 999 25122
rect 0 25064 938 25120
rect 994 25064 999 25120
rect 0 25062 999 25064
rect 0 25032 800 25062
rect 933 25059 999 25062
rect 37457 25122 37523 25125
rect 38200 25122 39000 25152
rect 37457 25120 39000 25122
rect 37457 25064 37462 25120
rect 37518 25064 39000 25120
rect 37457 25062 39000 25064
rect 37457 25059 37523 25062
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 38200 25032 39000 25062
rect 19570 24991 19886 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 0 23490 800 23520
rect 933 23490 999 23493
rect 0 23488 999 23490
rect 0 23432 938 23488
rect 994 23432 999 23488
rect 0 23430 999 23432
rect 0 23400 800 23430
rect 933 23427 999 23430
rect 37273 23490 37339 23493
rect 38200 23490 39000 23520
rect 37273 23488 39000 23490
rect 37273 23432 37278 23488
rect 37334 23432 39000 23488
rect 37273 23430 39000 23432
rect 37273 23427 37339 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 38200 23400 39000 23430
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 1577 21994 1643 21997
rect 798 21992 1643 21994
rect 798 21936 1582 21992
rect 1638 21936 1643 21992
rect 798 21934 1643 21936
rect 798 21888 858 21934
rect 1577 21931 1643 21934
rect 0 21798 858 21888
rect 37457 21858 37523 21861
rect 38200 21858 39000 21888
rect 37457 21856 39000 21858
rect 37457 21800 37462 21856
rect 37518 21800 39000 21856
rect 37457 21798 39000 21800
rect 0 21768 800 21798
rect 37457 21795 37523 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 38200 21768 39000 21798
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 0 20226 800 20256
rect 933 20226 999 20229
rect 0 20224 999 20226
rect 0 20168 938 20224
rect 994 20168 999 20224
rect 0 20166 999 20168
rect 0 20136 800 20166
rect 933 20163 999 20166
rect 37273 20226 37339 20229
rect 38200 20226 39000 20256
rect 37273 20224 39000 20226
rect 37273 20168 37278 20224
rect 37334 20168 39000 20224
rect 37273 20166 39000 20168
rect 37273 20163 37339 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 38200 20136 39000 20166
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 0 18594 800 18624
rect 1577 18594 1643 18597
rect 0 18592 1643 18594
rect 0 18536 1582 18592
rect 1638 18536 1643 18592
rect 0 18534 1643 18536
rect 0 18504 800 18534
rect 1577 18531 1643 18534
rect 36905 18594 36971 18597
rect 38200 18594 39000 18624
rect 36905 18592 39000 18594
rect 36905 18536 36910 18592
rect 36966 18536 39000 18592
rect 36905 18534 39000 18536
rect 36905 18531 36971 18534
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 38200 18504 39000 18534
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 0 16962 800 16992
rect 37181 16962 37247 16965
rect 38200 16962 39000 16992
rect 0 16872 858 16962
rect 37181 16960 39000 16962
rect 37181 16904 37186 16960
rect 37242 16904 39000 16960
rect 37181 16902 39000 16904
rect 37181 16899 37247 16902
rect 798 16690 858 16872
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 38200 16872 39000 16902
rect 34930 16831 35246 16832
rect 1577 16690 1643 16693
rect 798 16688 1643 16690
rect 798 16632 1582 16688
rect 1638 16632 1643 16688
rect 798 16630 1643 16632
rect 1577 16627 1643 16630
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 0 15330 800 15360
rect 1577 15330 1643 15333
rect 0 15328 1643 15330
rect 0 15272 1582 15328
rect 1638 15272 1643 15328
rect 0 15270 1643 15272
rect 0 15240 800 15270
rect 1577 15267 1643 15270
rect 36905 15330 36971 15333
rect 38200 15330 39000 15360
rect 36905 15328 39000 15330
rect 36905 15272 36910 15328
rect 36966 15272 39000 15328
rect 36905 15270 39000 15272
rect 36905 15267 36971 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 38200 15240 39000 15270
rect 19570 15199 19886 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 0 13698 800 13728
rect 933 13698 999 13701
rect 0 13696 999 13698
rect 0 13640 938 13696
rect 994 13640 999 13696
rect 0 13638 999 13640
rect 0 13608 800 13638
rect 933 13635 999 13638
rect 37273 13698 37339 13701
rect 38200 13698 39000 13728
rect 37273 13696 39000 13698
rect 37273 13640 37278 13696
rect 37334 13640 39000 13696
rect 37273 13638 39000 13640
rect 37273 13635 37339 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 38200 13608 39000 13638
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 0 12066 800 12096
rect 933 12066 999 12069
rect 0 12064 999 12066
rect 0 12008 938 12064
rect 994 12008 999 12064
rect 0 12006 999 12008
rect 0 11976 800 12006
rect 933 12003 999 12006
rect 37457 12066 37523 12069
rect 38200 12066 39000 12096
rect 37457 12064 39000 12066
rect 37457 12008 37462 12064
rect 37518 12008 39000 12064
rect 37457 12006 39000 12008
rect 37457 12003 37523 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 38200 11976 39000 12006
rect 19570 11935 19886 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 0 10434 800 10464
rect 933 10434 999 10437
rect 0 10432 999 10434
rect 0 10376 938 10432
rect 994 10376 999 10432
rect 0 10374 999 10376
rect 0 10344 800 10374
rect 933 10371 999 10374
rect 37273 10434 37339 10437
rect 38200 10434 39000 10464
rect 37273 10432 39000 10434
rect 37273 10376 37278 10432
rect 37334 10376 39000 10432
rect 37273 10374 39000 10376
rect 37273 10371 37339 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 38200 10344 39000 10374
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 0 8802 800 8832
rect 933 8802 999 8805
rect 0 8800 999 8802
rect 0 8744 938 8800
rect 994 8744 999 8800
rect 0 8742 999 8744
rect 0 8712 800 8742
rect 933 8739 999 8742
rect 37457 8802 37523 8805
rect 38200 8802 39000 8832
rect 37457 8800 39000 8802
rect 37457 8744 37462 8800
rect 37518 8744 39000 8800
rect 37457 8742 39000 8744
rect 37457 8739 37523 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 38200 8712 39000 8742
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 0 7170 800 7200
rect 37181 7170 37247 7173
rect 38200 7170 39000 7200
rect 0 7110 1640 7170
rect 0 7080 800 7110
rect 1580 7037 1640 7110
rect 37181 7168 39000 7170
rect 37181 7112 37186 7168
rect 37242 7112 39000 7168
rect 37181 7110 39000 7112
rect 37181 7107 37247 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 38200 7080 39000 7110
rect 34930 7039 35246 7040
rect 1577 7032 1643 7037
rect 1577 6976 1582 7032
rect 1638 6976 1643 7032
rect 1577 6971 1643 6976
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 0 5538 800 5568
rect 933 5538 999 5541
rect 0 5536 999 5538
rect 0 5480 938 5536
rect 994 5480 999 5536
rect 0 5478 999 5480
rect 0 5448 800 5478
rect 933 5475 999 5478
rect 37641 5538 37707 5541
rect 38200 5538 39000 5568
rect 37641 5536 39000 5538
rect 37641 5480 37646 5536
rect 37702 5480 39000 5536
rect 37641 5478 39000 5480
rect 37641 5475 37707 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 38200 5448 39000 5478
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 33041 4178 33107 4181
rect 36629 4178 36695 4181
rect 33041 4176 36695 4178
rect 33041 4120 33046 4176
rect 33102 4120 36634 4176
rect 36690 4120 36695 4176
rect 33041 4118 36695 4120
rect 33041 4115 33107 4118
rect 36629 4115 36695 4118
rect 34605 4042 34671 4045
rect 34605 4040 35450 4042
rect 34605 3984 34610 4040
rect 34666 3984 35450 4040
rect 34605 3982 35450 3984
rect 34605 3979 34671 3982
rect 0 3906 800 3936
rect 933 3906 999 3909
rect 0 3904 999 3906
rect 0 3848 938 3904
rect 994 3848 999 3904
rect 0 3846 999 3848
rect 35390 3906 35450 3982
rect 38200 3906 39000 3936
rect 35390 3846 39000 3906
rect 0 3816 800 3846
rect 933 3843 999 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 38200 3816 39000 3846
rect 34930 3775 35246 3776
rect 30649 3770 30715 3773
rect 33593 3770 33659 3773
rect 30649 3768 33659 3770
rect 30649 3712 30654 3768
rect 30710 3712 33598 3768
rect 33654 3712 33659 3768
rect 30649 3710 33659 3712
rect 30649 3707 30715 3710
rect 33593 3707 33659 3710
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 20621 3090 20687 3093
rect 36261 3090 36327 3093
rect 20621 3088 36327 3090
rect 20621 3032 20626 3088
rect 20682 3032 36266 3088
rect 36322 3032 36327 3088
rect 20621 3030 36327 3032
rect 20621 3027 20687 3030
rect 36261 3027 36327 3030
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 1577 2680 1643 2685
rect 1577 2624 1582 2680
rect 1638 2624 1643 2680
rect 1577 2619 1643 2624
rect 0 2274 800 2304
rect 1580 2274 1640 2619
rect 0 2214 1640 2274
rect 37917 2274 37983 2277
rect 38200 2274 39000 2304
rect 37917 2272 39000 2274
rect 37917 2216 37922 2272
rect 37978 2216 39000 2272
rect 37917 2214 39000 2216
rect 0 2184 800 2214
rect 37917 2211 37983 2214
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 38200 2184 39000 2214
rect 19570 2143 19886 2144
rect 34513 642 34579 645
rect 38200 642 39000 672
rect 34513 640 39000 642
rect 34513 584 34518 640
rect 34574 584 39000 640
rect 34513 582 39000 584
rect 34513 579 34579 582
rect 38200 552 39000 582
<< via3 >>
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 36480 4528 36496
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 35936 19888 36496
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 36480 35248 36496
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__and2b_1  _088_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15180 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _089_
timestamp 1688980957
transform -1 0 16836 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _090_
timestamp 1688980957
transform 1 0 18492 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _091_
timestamp 1688980957
transform -1 0 20516 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _092_
timestamp 1688980957
transform -1 0 22448 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _093_
timestamp 1688980957
transform -1 0 25392 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _094_
timestamp 1688980957
transform -1 0 26772 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _095_
timestamp 1688980957
transform -1 0 27968 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _096_
timestamp 1688980957
transform -1 0 29072 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _097_
timestamp 1688980957
transform 1 0 29624 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _098_
timestamp 1688980957
transform -1 0 37076 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _099_
timestamp 1688980957
transform -1 0 35972 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _100_
timestamp 1688980957
transform 1 0 32568 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _101_
timestamp 1688980957
transform 1 0 27048 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _102_
timestamp 1688980957
transform 1 0 25760 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _103_
timestamp 1688980957
transform -1 0 25392 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _104_
timestamp 1688980957
transform 1 0 26312 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _105_
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _106_
timestamp 1688980957
transform 1 0 29624 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _107_
timestamp 1688980957
transform -1 0 31924 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _108_
timestamp 1688980957
transform -1 0 34500 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _109_
timestamp 1688980957
transform -1 0 35604 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _110_
timestamp 1688980957
transform 1 0 32200 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _111_
timestamp 1688980957
transform -1 0 35972 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _112_
timestamp 1688980957
transform 1 0 34776 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _113_
timestamp 1688980957
transform 1 0 34408 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _114_
timestamp 1688980957
transform 1 0 34776 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _115_
timestamp 1688980957
transform 1 0 34408 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _116_
timestamp 1688980957
transform 1 0 34776 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _117_
timestamp 1688980957
transform 1 0 34408 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _118_
timestamp 1688980957
transform 1 0 34776 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _119_
timestamp 1688980957
transform 1 0 34408 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _120_
timestamp 1688980957
transform -1 0 37444 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _121_
timestamp 1688980957
transform -1 0 36064 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _122_
timestamp 1688980957
transform 1 0 34776 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _123_
timestamp 1688980957
transform 1 0 34408 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _124_
timestamp 1688980957
transform 1 0 34776 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _125_
timestamp 1688980957
transform 1 0 34408 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _126_
timestamp 1688980957
transform 1 0 34776 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _127_
timestamp 1688980957
transform 1 0 34776 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _128_
timestamp 1688980957
transform -1 0 32752 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _129_
timestamp 1688980957
transform -1 0 37444 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _130_
timestamp 1688980957
transform -1 0 37444 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _131_
timestamp 1688980957
transform 1 0 21068 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _132_
timestamp 1688980957
transform 1 0 11592 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _133_
timestamp 1688980957
transform 1 0 9384 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _134_
timestamp 1688980957
transform 1 0 10120 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _135_
timestamp 1688980957
transform -1 0 13984 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _136_
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _137_
timestamp 1688980957
transform -1 0 15732 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _138_
timestamp 1688980957
transform -1 0 19412 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _139_
timestamp 1688980957
transform 1 0 18400 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _140_
timestamp 1688980957
transform 1 0 17112 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _141_
timestamp 1688980957
transform -1 0 12328 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _142_
timestamp 1688980957
transform -1 0 3956 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _143_
timestamp 1688980957
transform -1 0 5060 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _144_
timestamp 1688980957
transform -1 0 4140 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _145_
timestamp 1688980957
transform -1 0 4876 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _146_
timestamp 1688980957
transform -1 0 5428 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _147_
timestamp 1688980957
transform -1 0 5060 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _148_
timestamp 1688980957
transform -1 0 5428 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _149_
timestamp 1688980957
transform -1 0 5060 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _150_
timestamp 1688980957
transform -1 0 4876 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _151_
timestamp 1688980957
transform -1 0 4232 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _152_
timestamp 1688980957
transform -1 0 5060 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _153_
timestamp 1688980957
transform -1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _154_
timestamp 1688980957
transform -1 0 3404 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _155_
timestamp 1688980957
transform -1 0 4140 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _156_
timestamp 1688980957
transform -1 0 4140 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _157_
timestamp 1688980957
transform -1 0 4140 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _158_
timestamp 1688980957
transform -1 0 4140 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _159_
timestamp 1688980957
transform -1 0 4140 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _160_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4968 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _161_
timestamp 1688980957
transform -1 0 17296 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _162_
timestamp 1688980957
transform -1 0 20792 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _163_
timestamp 1688980957
transform 1 0 21436 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _164_
timestamp 1688980957
transform -1 0 20884 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _165_
timestamp 1688980957
transform 1 0 12788 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _166_
timestamp 1688980957
transform 1 0 3772 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _167_
timestamp 1688980957
transform 1 0 2852 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _168_
timestamp 1688980957
transform -1 0 4876 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _169_
timestamp 1688980957
transform 1 0 1472 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _170_
timestamp 1688980957
transform -1 0 4324 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _171_
timestamp 1688980957
transform -1 0 6900 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _172_
timestamp 1688980957
transform 1 0 7176 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _173_
timestamp 1688980957
transform -1 0 9476 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _174_
timestamp 1688980957
transform -1 0 12052 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _175_
timestamp 1688980957
transform 1 0 12696 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _176_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14720 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _177_
timestamp 1688980957
transform -1 0 16284 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _178_
timestamp 1688980957
transform -1 0 18308 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _179_
timestamp 1688980957
transform -1 0 20700 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _180_
timestamp 1688980957
transform -1 0 22632 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _181_
timestamp 1688980957
transform 1 0 22816 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _182_
timestamp 1688980957
transform -1 0 26312 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _183_
timestamp 1688980957
transform 1 0 26496 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _184_
timestamp 1688980957
transform 1 0 27968 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _185_
timestamp 1688980957
transform 1 0 29808 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _186_
timestamp 1688980957
transform 1 0 31648 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _187_
timestamp 1688980957
transform -1 0 34592 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _188_
timestamp 1688980957
transform -1 0 33580 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _189_
timestamp 1688980957
transform 1 0 28244 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _190_
timestamp 1688980957
transform -1 0 28428 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _191_
timestamp 1688980957
transform 1 0 24656 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _192_
timestamp 1688980957
transform 1 0 27600 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _193_
timestamp 1688980957
transform 1 0 27508 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _194_
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _195_
timestamp 1688980957
transform 1 0 31004 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _196_
timestamp 1688980957
transform 1 0 32476 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _197_
timestamp 1688980957
transform 1 0 33120 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _198_
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _199_
timestamp 1688980957
transform 1 0 32752 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _200_
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _201_
timestamp 1688980957
transform 1 0 35420 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _202_
timestamp 1688980957
transform 1 0 35420 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _203_
timestamp 1688980957
transform 1 0 35420 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _204_
timestamp 1688980957
transform 1 0 35420 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _205_
timestamp 1688980957
transform 1 0 35420 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _206_
timestamp 1688980957
transform 1 0 35420 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _207_
timestamp 1688980957
transform 1 0 35420 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _208_
timestamp 1688980957
transform -1 0 36892 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _209_
timestamp 1688980957
transform 1 0 35420 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _210_
timestamp 1688980957
transform 1 0 35420 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _211_
timestamp 1688980957
transform 1 0 35420 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _212_
timestamp 1688980957
transform 1 0 35420 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _213_
timestamp 1688980957
transform 1 0 35420 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _214_
timestamp 1688980957
transform 1 0 35420 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _215_
timestamp 1688980957
transform 1 0 35420 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _216_
timestamp 1688980957
transform 1 0 35420 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _217_
timestamp 1688980957
transform -1 0 35420 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _218_
timestamp 1688980957
transform -1 0 36892 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _219_
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _220_
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _221_
timestamp 1688980957
transform 1 0 10764 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _222_
timestamp 1688980957
transform -1 0 12144 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _223_
timestamp 1688980957
transform 1 0 11776 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _224_
timestamp 1688980957
transform -1 0 14720 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _225_
timestamp 1688980957
transform -1 0 16008 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _226_
timestamp 1688980957
transform -1 0 17480 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _227_
timestamp 1688980957
transform -1 0 18952 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _228_
timestamp 1688980957
transform 1 0 17388 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _229_
timestamp 1688980957
transform 1 0 14168 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _230_
timestamp 1688980957
transform 1 0 2208 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _231_
timestamp 1688980957
transform 1 0 1932 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _232_
timestamp 1688980957
transform -1 0 3404 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _233_
timestamp 1688980957
transform 1 0 1932 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _234_
timestamp 1688980957
transform 1 0 1932 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _235_
timestamp 1688980957
transform 1 0 1932 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _236_
timestamp 1688980957
transform 1 0 1932 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _237_
timestamp 1688980957
transform -1 0 3404 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _238_
timestamp 1688980957
transform -1 0 3404 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _239_
timestamp 1688980957
transform 1 0 1932 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _240_
timestamp 1688980957
transform -1 0 3404 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _241_
timestamp 1688980957
transform -1 0 3404 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _242_
timestamp 1688980957
transform 1 0 1932 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _243_
timestamp 1688980957
transform 1 0 1932 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _244_
timestamp 1688980957
transform 1 0 1932 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _245_
timestamp 1688980957
transform 1 0 1932 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _246_
timestamp 1688980957
transform -1 0 3404 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _247_
timestamp 1688980957
transform -1 0 3404 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _248_
timestamp 1688980957
transform 1 0 1932 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _249_
timestamp 1688980957
transform -1 0 14904 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _250_
timestamp 1688980957
transform -1 0 20792 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _251_
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _252_
timestamp 1688980957
transform 1 0 20148 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _253_
timestamp 1688980957
transform 1 0 15456 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _254_
timestamp 1688980957
transform 1 0 4692 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _255_
timestamp 1688980957
transform -1 0 4324 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _256_
timestamp 1688980957
transform -1 0 3404 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _257_
timestamp 1688980957
transform 1 0 1932 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _258_
timestamp 1688980957
transform -1 0 4232 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _259_
timestamp 1688980957
transform -1 0 5888 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _260_
timestamp 1688980957
transform -1 0 7360 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _261_
timestamp 1688980957
transform -1 0 8832 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _262_
timestamp 1688980957
transform -1 0 11408 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _263_
timestamp 1688980957
transform -1 0 13616 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A_N dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15364 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A_N
timestamp 1688980957
transform 1 0 16836 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A_N
timestamp 1688980957
transform 1 0 18308 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A_N
timestamp 1688980957
transform 1 0 20700 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A_N
timestamp 1688980957
transform 1 0 22632 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A_N
timestamp 1688980957
transform 1 0 25392 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A_N
timestamp 1688980957
transform 1 0 26956 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A_N
timestamp 1688980957
transform 1 0 27968 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A_N
timestamp 1688980957
transform 1 0 28704 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A_N
timestamp 1688980957
transform 1 0 32660 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A_N
timestamp 1688980957
transform 1 0 36340 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A_N
timestamp 1688980957
transform -1 0 37260 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A_N
timestamp 1688980957
transform 1 0 32292 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A_N
timestamp 1688980957
transform -1 0 27968 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A_N
timestamp 1688980957
transform 1 0 26312 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A_N
timestamp 1688980957
transform 1 0 25392 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A_N
timestamp 1688980957
transform 1 0 25208 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A_N
timestamp 1688980957
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A_N
timestamp 1688980957
transform 1 0 30176 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A_N
timestamp 1688980957
transform -1 0 33304 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A_N
timestamp 1688980957
transform 1 0 34776 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A_N
timestamp 1688980957
transform 1 0 36708 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A_N
timestamp 1688980957
transform 1 0 35236 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A_N
timestamp 1688980957
transform -1 0 37260 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A_N
timestamp 1688980957
transform 1 0 34408 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A_N
timestamp 1688980957
transform 1 0 34960 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A_N
timestamp 1688980957
transform 1 0 34408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A_N
timestamp 1688980957
transform 1 0 34960 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A_N
timestamp 1688980957
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A_N
timestamp 1688980957
transform 1 0 34960 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A_N
timestamp 1688980957
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A_N
timestamp 1688980957
transform 1 0 34224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A_N
timestamp 1688980957
transform -1 0 36892 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A_N
timestamp 1688980957
transform 1 0 36064 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A_N
timestamp 1688980957
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A_N
timestamp 1688980957
transform 1 0 34960 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A_N
timestamp 1688980957
transform 1 0 34408 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A_N
timestamp 1688980957
transform 1 0 34960 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A_N
timestamp 1688980957
transform 1 0 36708 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__A_N
timestamp 1688980957
transform 1 0 36708 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__128__A_N
timestamp 1688980957
transform 1 0 33488 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A_N
timestamp 1688980957
transform -1 0 36156 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__A_N
timestamp 1688980957
transform -1 0 37536 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__A_N
timestamp 1688980957
transform 1 0 21804 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__B
timestamp 1688980957
transform -1 0 21068 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__A_N
timestamp 1688980957
transform -1 0 12512 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A_N
timestamp 1688980957
transform 1 0 9936 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A_N
timestamp 1688980957
transform 1 0 10672 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A_N
timestamp 1688980957
transform 1 0 13984 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__A_N
timestamp 1688980957
transform 1 0 14812 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__A_N
timestamp 1688980957
transform 1 0 15916 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__A_N
timestamp 1688980957
transform -1 0 20700 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A_N
timestamp 1688980957
transform 1 0 19412 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A_N
timestamp 1688980957
transform 1 0 17848 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__A_N
timestamp 1688980957
transform 1 0 12512 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A_N
timestamp 1688980957
transform 1 0 4416 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A_N
timestamp 1688980957
transform 1 0 5244 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__153__A_N
timestamp 1688980957
transform 1 0 5888 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A_N
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A_N
timestamp 1688980957
transform 1 0 4324 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A_N
timestamp 1688980957
transform 1 0 4324 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A_N
timestamp 1688980957
transform 1 0 4324 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A_N
timestamp 1688980957
transform 1 0 4324 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__161__A_N
timestamp 1688980957
transform 1 0 17296 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__A_N
timestamp 1688980957
transform 1 0 20976 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__A_N
timestamp 1688980957
transform 1 0 21988 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__164__A_N
timestamp 1688980957
transform -1 0 20332 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__165__A_N
timestamp 1688980957
transform 1 0 13524 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__166__A_N
timestamp 1688980957
transform 1 0 4508 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__A_N
timestamp 1688980957
transform 1 0 3956 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__A_N
timestamp 1688980957
transform 1 0 9660 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A_N
timestamp 1688980957
transform 1 0 12052 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__175__A_N
timestamp 1688980957
transform 1 0 13248 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__179__CLK
timestamp 1688980957
transform 1 0 20884 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__CLK
timestamp 1688980957
transform 1 0 23000 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__CLK
timestamp 1688980957
transform 1 0 24564 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__CLK
timestamp 1688980957
transform -1 0 27324 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__183__CLK
timestamp 1688980957
transform -1 0 28612 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__CLK
timestamp 1688980957
transform -1 0 31648 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__185__CLK
timestamp 1688980957
transform -1 0 31556 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__CLK
timestamp 1688980957
transform -1 0 30084 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__CLK
timestamp 1688980957
transform -1 0 31096 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__191__CLK
timestamp 1688980957
transform 1 0 26312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__CLK
timestamp 1688980957
transform 1 0 29072 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__CLK
timestamp 1688980957
transform -1 0 29624 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__CLK
timestamp 1688980957
transform 1 0 29716 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__CLK
timestamp 1688980957
transform -1 0 33304 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__CLK
timestamp 1688980957
transform -1 0 26220 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__250__CLK
timestamp 1688980957
transform 1 0 20976 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__CLK
timestamp 1688980957
transform 1 0 23460 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__CLK
timestamp 1688980957
transform 1 0 22172 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0__f_wb_clk_i_A
timestamp 1688980957
transform -1 0 10028 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1__f_wb_clk_i_A
timestamp 1688980957
transform 1 0 12420 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2__f_wb_clk_i_A
timestamp 1688980957
transform 1 0 7268 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3__f_wb_clk_i_A
timestamp 1688980957
transform 1 0 9844 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4__f_wb_clk_i_A
timestamp 1688980957
transform -1 0 28612 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5__f_wb_clk_i_A
timestamp 1688980957
transform 1 0 31004 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6__f_wb_clk_i_A
timestamp 1688980957
transform 1 0 28428 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7__f_wb_clk_i_A
timestamp 1688980957
transform 1 0 31004 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout90_A
timestamp 1688980957
transform 1 0 16836 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout91_A
timestamp 1688980957
transform -1 0 1932 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout92_A
timestamp 1688980957
transform 1 0 17848 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout93_A
timestamp 1688980957
transform 1 0 36708 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout94_A
timestamp 1688980957
transform 1 0 35328 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout95_A
timestamp 1688980957
transform 1 0 36984 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold330_A
timestamp 1688980957
transform 1 0 16928 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 21712 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_wb_clk_i
timestamp 1688980957
transform -1 0 9660 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_wb_clk_i
timestamp 1688980957
transform 1 0 10396 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_wb_clk_i
timestamp 1688980957
transform -1 0 7084 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_wb_clk_i
timestamp 1688980957
transform -1 0 9660 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_wb_clk_i
timestamp 1688980957
transform 1 0 28612 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_wb_clk_i
timestamp 1688980957
transform 1 0 31188 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_wb_clk_i
timestamp 1688980957
transform -1 0 30452 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_wb_clk_i
timestamp 1688980957
transform 1 0 31188 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout90 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout91
timestamp 1688980957
transform -1 0 1932 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout92 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17664 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout93 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 35420 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout94
timestamp 1688980957
transform 1 0 35512 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout95
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout96
timestamp 1688980957
transform -1 0 37444 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_9 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_19 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_23
timestamp 1688980957
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_29 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_65 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_91
timestamp 1688980957
transform 1 0 9476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_95
timestamp 1688980957
transform 1 0 9844 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_177
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1688980957
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_234 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22632 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_246
timestamp 1688980957
transform 1 0 23736 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_269
timestamp 1688980957
transform 1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1688980957
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_346 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32936 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_350
timestamp 1688980957
transform 1 0 33304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 1688980957
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 1688980957
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_22
timestamp 1688980957
transform 1 0 3128 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_34
timestamp 1688980957
transform 1 0 4232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_46
timestamp 1688980957
transform 1 0 5336 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 1688980957
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_63
timestamp 1688980957
transform 1 0 6900 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_80
timestamp 1688980957
transform 1 0 8464 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_86
timestamp 1688980957
transform 1 0 9016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_96
timestamp 1688980957
transform 1 0 9936 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_102
timestamp 1688980957
transform 1 0 10488 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_120
timestamp 1688980957
transform 1 0 12144 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_124
timestamp 1688980957
transform 1 0 12512 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_136
timestamp 1688980957
transform 1 0 13616 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_142
timestamp 1688980957
transform 1 0 14168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_199
timestamp 1688980957
transform 1 0 19412 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_209
timestamp 1688980957
transform 1 0 20332 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_213
timestamp 1688980957
transform 1 0 20700 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_221
timestamp 1688980957
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_250
timestamp 1688980957
transform 1 0 24104 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_306
timestamp 1688980957
transform 1 0 29256 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_310
timestamp 1688980957
transform 1 0 29624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_322
timestamp 1688980957
transform 1 0 30728 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_326
timestamp 1688980957
transform 1 0 31096 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_346
timestamp 1688980957
transform 1 0 32936 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_350
timestamp 1688980957
transform 1 0 33304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_375
timestamp 1688980957
transform 1 0 35604 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_385
timestamp 1688980957
transform 1 0 36524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_389
timestamp 1688980957
transform 1 0 36892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_19
timestamp 1688980957
transform 1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_68
timestamp 1688980957
transform 1 0 7360 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_74
timestamp 1688980957
transform 1 0 7912 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_93
timestamp 1688980957
transform 1 0 9660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_137
timestamp 1688980957
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_145
timestamp 1688980957
transform 1 0 14444 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_194
timestamp 1688980957
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_205
timestamp 1688980957
transform 1 0 19964 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_217
timestamp 1688980957
transform 1 0 21068 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_229
timestamp 1688980957
transform 1 0 22172 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_241
timestamp 1688980957
transform 1 0 23276 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_249
timestamp 1688980957
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_272
timestamp 1688980957
transform 1 0 26128 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_276
timestamp 1688980957
transform 1 0 26496 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_304
timestamp 1688980957
transform 1 0 29072 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_395
timestamp 1688980957
transform 1 0 37444 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_9
timestamp 1688980957
transform 1 0 1932 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_19
timestamp 1688980957
transform 1 0 2852 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_31
timestamp 1688980957
transform 1 0 3956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_43
timestamp 1688980957
transform 1 0 5060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_87
timestamp 1688980957
transform 1 0 9108 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_148
timestamp 1688980957
transform 1 0 14720 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_189
timestamp 1688980957
transform 1 0 18492 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_195
timestamp 1688980957
transform 1 0 19044 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_204
timestamp 1688980957
transform 1 0 19872 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_216
timestamp 1688980957
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_257
timestamp 1688980957
transform 1 0 24748 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_303
timestamp 1688980957
transform 1 0 28980 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_345
timestamp 1688980957
transform 1 0 32844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_364
timestamp 1688980957
transform 1 0 34592 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_368
timestamp 1688980957
transform 1 0 34960 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_388
timestamp 1688980957
transform 1 0 36800 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_19
timestamp 1688980957
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_89
timestamp 1688980957
transform 1 0 9292 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_120
timestamp 1688980957
transform 1 0 12144 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_149
timestamp 1688980957
transform 1 0 14812 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_159
timestamp 1688980957
transform 1 0 15732 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_176
timestamp 1688980957
transform 1 0 17296 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_194
timestamp 1688980957
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_201
timestamp 1688980957
transform 1 0 19596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_213
timestamp 1688980957
transform 1 0 20700 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_225
timestamp 1688980957
transform 1 0 21804 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_237
timestamp 1688980957
transform 1 0 22908 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_249
timestamp 1688980957
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_261
timestamp 1688980957
transform 1 0 25116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_266
timestamp 1688980957
transform 1 0 25576 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_306
timestamp 1688980957
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_379
timestamp 1688980957
transform 1 0 35972 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_9
timestamp 1688980957
transform 1 0 1932 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_147
timestamp 1688980957
transform 1 0 14628 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_158
timestamp 1688980957
transform 1 0 15640 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_165
timestamp 1688980957
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_173
timestamp 1688980957
transform 1 0 17020 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_180
timestamp 1688980957
transform 1 0 17664 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_184
timestamp 1688980957
transform 1 0 18032 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_196
timestamp 1688980957
transform 1 0 19136 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_208
timestamp 1688980957
transform 1 0 20240 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_220
timestamp 1688980957
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_276
timestamp 1688980957
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_291
timestamp 1688980957
transform 1 0 27876 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_326
timestamp 1688980957
transform 1 0 31096 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_369
timestamp 1688980957
transform 1 0 35052 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_389
timestamp 1688980957
transform 1 0 36892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_9
timestamp 1688980957
transform 1 0 1932 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_103
timestamp 1688980957
transform 1 0 10580 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_106
timestamp 1688980957
transform 1 0 10856 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_115
timestamp 1688980957
transform 1 0 11684 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_132
timestamp 1688980957
transform 1 0 13248 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_147
timestamp 1688980957
transform 1 0 14628 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_151
timestamp 1688980957
transform 1 0 14996 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_159
timestamp 1688980957
transform 1 0 15732 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_163
timestamp 1688980957
transform 1 0 16100 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_175
timestamp 1688980957
transform 1 0 17204 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_187
timestamp 1688980957
transform 1 0 18308 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_306
timestamp 1688980957
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_313
timestamp 1688980957
transform 1 0 29900 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_318
timestamp 1688980957
transform 1 0 30360 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_379
timestamp 1688980957
transform 1 0 35972 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_393
timestamp 1688980957
transform 1 0 37260 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_35
timestamp 1688980957
transform 1 0 4324 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_47
timestamp 1688980957
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_142
timestamp 1688980957
transform 1 0 14168 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_154
timestamp 1688980957
transform 1 0 15272 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_166
timestamp 1688980957
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_197
timestamp 1688980957
transform 1 0 19228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_209
timestamp 1688980957
transform 1 0 20332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_221
timestamp 1688980957
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_357
timestamp 1688980957
transform 1 0 33948 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_389
timestamp 1688980957
transform 1 0 36892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_25
timestamp 1688980957
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_43
timestamp 1688980957
transform 1 0 5060 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_47
timestamp 1688980957
transform 1 0 5428 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_59
timestamp 1688980957
transform 1 0 6532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_71
timestamp 1688980957
transform 1 0 7636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_339
timestamp 1688980957
transform 1 0 32292 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_25
timestamp 1688980957
transform 1 0 3404 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_50
timestamp 1688980957
transform 1 0 5704 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_54
timestamp 1688980957
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_97
timestamp 1688980957
transform 1 0 10028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_109
timestamp 1688980957
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1688980957
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_319
timestamp 1688980957
transform 1 0 30452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_331
timestamp 1688980957
transform 1 0 31556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1688980957
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1688980957
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_25
timestamp 1688980957
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_37
timestamp 1688980957
transform 1 0 4508 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_49
timestamp 1688980957
transform 1 0 5612 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_61
timestamp 1688980957
transform 1 0 6716 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_73
timestamp 1688980957
transform 1 0 7820 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_81
timestamp 1688980957
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_125
timestamp 1688980957
transform 1 0 12604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_137
timestamp 1688980957
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_205
timestamp 1688980957
transform 1 0 19964 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_217
timestamp 1688980957
transform 1 0 21068 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_229
timestamp 1688980957
transform 1 0 22172 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_241
timestamp 1688980957
transform 1 0 23276 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_249
timestamp 1688980957
transform 1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1688980957
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1688980957
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_345
timestamp 1688980957
transform 1 0 32844 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_353
timestamp 1688980957
transform 1 0 33580 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_395
timestamp 1688980957
transform 1 0 37444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_25
timestamp 1688980957
transform 1 0 3404 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_29
timestamp 1688980957
transform 1 0 3772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_41
timestamp 1688980957
transform 1 0 4876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_53
timestamp 1688980957
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1688980957
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1688980957
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1688980957
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1688980957
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1688980957
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1688980957
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1688980957
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1688980957
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1688980957
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_361
timestamp 1688980957
transform 1 0 34316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_9
timestamp 1688980957
transform 1 0 1932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1688980957
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1688980957
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1688980957
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1688980957
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1688980957
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1688980957
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 1688980957
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1688980957
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1688980957
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1688980957
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1688980957
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1688980957
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1688980957
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1688980957
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 1688980957
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 1688980957
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1688980957
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_370
timestamp 1688980957
transform 1 0 35144 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_389
timestamp 1688980957
transform 1 0 36892 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_395
timestamp 1688980957
transform 1 0 37444 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_33
timestamp 1688980957
transform 1 0 4140 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_45
timestamp 1688980957
transform 1 0 5244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 1688980957
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1688980957
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1688980957
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1688980957
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1688980957
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1688980957
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1688980957
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1688980957
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1688980957
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 1688980957
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 1688980957
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 1688980957
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1688980957
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1688980957
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1688980957
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1688980957
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1688980957
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1688980957
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1688980957
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 1688980957
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 1688980957
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_329
timestamp 1688980957
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 1688980957
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_349
timestamp 1688980957
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_361
timestamp 1688980957
transform 1 0 34316 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_389
timestamp 1688980957
transform 1 0 36892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_393
timestamp 1688980957
transform 1 0 37260 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_37
timestamp 1688980957
transform 1 0 4508 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_49
timestamp 1688980957
transform 1 0 5612 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_61
timestamp 1688980957
transform 1 0 6716 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_71
timestamp 1688980957
transform 1 0 7636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1688980957
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1688980957
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1688980957
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1688980957
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1688980957
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1688980957
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_165
timestamp 1688980957
transform 1 0 16284 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_171
timestamp 1688980957
transform 1 0 16836 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 1688980957
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 1688980957
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1688980957
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 1688980957
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 1688980957
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_233
timestamp 1688980957
transform 1 0 22540 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_245
timestamp 1688980957
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1688980957
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1688980957
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 1688980957
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_289
timestamp 1688980957
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_301
timestamp 1688980957
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1688980957
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_321
timestamp 1688980957
transform 1 0 30636 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_347
timestamp 1688980957
transform 1 0 33028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_359
timestamp 1688980957
transform 1 0 34132 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_365
timestamp 1688980957
transform 1 0 34684 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_9
timestamp 1688980957
transform 1 0 1932 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_33
timestamp 1688980957
transform 1 0 4140 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_37
timestamp 1688980957
transform 1 0 4508 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_49
timestamp 1688980957
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1688980957
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1688980957
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1688980957
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1688980957
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1688980957
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1688980957
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1688980957
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 1688980957
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1688980957
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_183
timestamp 1688980957
transform 1 0 17940 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_195
timestamp 1688980957
transform 1 0 19044 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_207
timestamp 1688980957
transform 1 0 20148 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_219
timestamp 1688980957
transform 1 0 21252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1688980957
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 1688980957
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_249
timestamp 1688980957
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_261
timestamp 1688980957
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_273
timestamp 1688980957
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1688980957
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_281
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_293
timestamp 1688980957
transform 1 0 28060 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_301
timestamp 1688980957
transform 1 0 28796 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_310
timestamp 1688980957
transform 1 0 29624 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_322
timestamp 1688980957
transform 1 0 30728 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_334
timestamp 1688980957
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_337
timestamp 1688980957
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_349
timestamp 1688980957
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_361
timestamp 1688980957
transform 1 0 34316 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_367
timestamp 1688980957
transform 1 0 34868 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_385
timestamp 1688980957
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_391
timestamp 1688980957
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_393
timestamp 1688980957
transform 1 0 37260 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_25
timestamp 1688980957
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_37
timestamp 1688980957
transform 1 0 4508 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_49
timestamp 1688980957
transform 1 0 5612 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_61
timestamp 1688980957
transform 1 0 6716 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_73
timestamp 1688980957
transform 1 0 7820 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_81
timestamp 1688980957
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1688980957
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1688980957
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1688980957
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1688980957
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 1688980957
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 1688980957
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 1688980957
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 1688980957
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1688980957
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 1688980957
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_221
timestamp 1688980957
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_233
timestamp 1688980957
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_245
timestamp 1688980957
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1688980957
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 1688980957
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 1688980957
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 1688980957
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 1688980957
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1688980957
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_321
timestamp 1688980957
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_333
timestamp 1688980957
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_345
timestamp 1688980957
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_357
timestamp 1688980957
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_363
timestamp 1688980957
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_389
timestamp 1688980957
transform 1 0 36892 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_395
timestamp 1688980957
transform 1 0 37444 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_33
timestamp 1688980957
transform 1 0 4140 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_37
timestamp 1688980957
transform 1 0 4508 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_49
timestamp 1688980957
transform 1 0 5612 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1688980957
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1688980957
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1688980957
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1688980957
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 1688980957
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 1688980957
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1688980957
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 1688980957
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_193
timestamp 1688980957
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_205
timestamp 1688980957
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 1688980957
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1688980957
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 1688980957
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 1688980957
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 1688980957
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 1688980957
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1688980957
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1688980957
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 1688980957
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 1688980957
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_329
timestamp 1688980957
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_335
timestamp 1688980957
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_337
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_349
timestamp 1688980957
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_361
timestamp 1688980957
transform 1 0 34316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_393
timestamp 1688980957
transform 1 0 37260 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_9
timestamp 1688980957
transform 1 0 1932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1688980957
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1688980957
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1688980957
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1688980957
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1688980957
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1688980957
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1688980957
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1688980957
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 1688980957
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_165
timestamp 1688980957
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 1688980957
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_189
timestamp 1688980957
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1688980957
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_209
timestamp 1688980957
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_221
timestamp 1688980957
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_233
timestamp 1688980957
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_245
timestamp 1688980957
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1688980957
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1688980957
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 1688980957
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 1688980957
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_301
timestamp 1688980957
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1688980957
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_321
timestamp 1688980957
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_333
timestamp 1688980957
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_345
timestamp 1688980957
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_357
timestamp 1688980957
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_363
timestamp 1688980957
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_365
timestamp 1688980957
transform 1 0 34684 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_370
timestamp 1688980957
transform 1 0 35144 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_389
timestamp 1688980957
transform 1 0 36892 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_395
timestamp 1688980957
transform 1 0 37444 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_33
timestamp 1688980957
transform 1 0 4140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_45
timestamp 1688980957
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_53
timestamp 1688980957
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1688980957
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1688980957
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1688980957
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1688980957
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1688980957
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1688980957
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_137
timestamp 1688980957
transform 1 0 13708 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_141
timestamp 1688980957
transform 1 0 14076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_158
timestamp 1688980957
transform 1 0 15640 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1688980957
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 1688980957
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_193
timestamp 1688980957
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_205
timestamp 1688980957
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_217
timestamp 1688980957
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1688980957
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_237
timestamp 1688980957
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_249
timestamp 1688980957
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_261
timestamp 1688980957
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_273
timestamp 1688980957
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1688980957
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1688980957
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1688980957
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_317
timestamp 1688980957
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_329
timestamp 1688980957
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_335
timestamp 1688980957
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_337
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_349
timestamp 1688980957
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_361
timestamp 1688980957
transform 1 0 34316 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_389
timestamp 1688980957
transform 1 0 36892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_393
timestamp 1688980957
transform 1 0 37260 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_37
timestamp 1688980957
transform 1 0 4508 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_49
timestamp 1688980957
transform 1 0 5612 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_57
timestamp 1688980957
transform 1 0 6348 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_67
timestamp 1688980957
transform 1 0 7268 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_79
timestamp 1688980957
transform 1 0 8372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1688980957
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_97
timestamp 1688980957
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 1688980957
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 1688980957
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 1688980957
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1688980957
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 1688980957
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 1688980957
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 1688980957
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 1688980957
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 1688980957
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_221
timestamp 1688980957
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_233
timestamp 1688980957
transform 1 0 22540 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_247
timestamp 1688980957
transform 1 0 23828 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1688980957
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_265
timestamp 1688980957
transform 1 0 25484 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_271
timestamp 1688980957
transform 1 0 26036 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_283
timestamp 1688980957
transform 1 0 27140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_295
timestamp 1688980957
transform 1 0 28244 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1688980957
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_321
timestamp 1688980957
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_333
timestamp 1688980957
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_345
timestamp 1688980957
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_357
timestamp 1688980957
transform 1 0 33948 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_361
timestamp 1688980957
transform 1 0 34316 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_365
timestamp 1688980957
transform 1 0 34684 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_9
timestamp 1688980957
transform 1 0 1932 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_33
timestamp 1688980957
transform 1 0 4140 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_37
timestamp 1688980957
transform 1 0 4508 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_49
timestamp 1688980957
transform 1 0 5612 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1688980957
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1688980957
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1688980957
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1688980957
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 1688980957
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 1688980957
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 1688980957
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1688980957
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 1688980957
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_193
timestamp 1688980957
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_205
timestamp 1688980957
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_217
timestamp 1688980957
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1688980957
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1688980957
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 1688980957
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_261
timestamp 1688980957
transform 1 0 25116 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_271
timestamp 1688980957
transform 1 0 26036 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1688980957
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 1688980957
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 1688980957
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_317
timestamp 1688980957
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_329
timestamp 1688980957
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_335
timestamp 1688980957
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_337
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_349
timestamp 1688980957
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_361
timestamp 1688980957
transform 1 0 34316 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_367
timestamp 1688980957
transform 1 0 34868 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_385
timestamp 1688980957
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_391
timestamp 1688980957
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_393
timestamp 1688980957
transform 1 0 37260 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_25
timestamp 1688980957
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_37
timestamp 1688980957
transform 1 0 4508 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_49
timestamp 1688980957
transform 1 0 5612 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_61
timestamp 1688980957
transform 1 0 6716 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_73
timestamp 1688980957
transform 1 0 7820 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_81
timestamp 1688980957
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1688980957
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1688980957
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 1688980957
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1688980957
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1688980957
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 1688980957
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 1688980957
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 1688980957
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 1688980957
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1688980957
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 1688980957
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_221
timestamp 1688980957
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_233
timestamp 1688980957
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_245
timestamp 1688980957
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1688980957
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1688980957
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 1688980957
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 1688980957
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 1688980957
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1688980957
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_321
timestamp 1688980957
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_333
timestamp 1688980957
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_345
timestamp 1688980957
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_357
timestamp 1688980957
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_363
timestamp 1688980957
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_389
timestamp 1688980957
transform 1 0 36892 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_395
timestamp 1688980957
transform 1 0 37444 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_33
timestamp 1688980957
transform 1 0 4140 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_37
timestamp 1688980957
transform 1 0 4508 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_49
timestamp 1688980957
transform 1 0 5612 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1688980957
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1688980957
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1688980957
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1688980957
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1688980957
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 1688980957
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 1688980957
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1688980957
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1688980957
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 1688980957
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_193
timestamp 1688980957
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_205
timestamp 1688980957
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 1688980957
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1688980957
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_229
timestamp 1688980957
transform 1 0 22172 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_241
timestamp 1688980957
transform 1 0 23276 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_253
timestamp 1688980957
transform 1 0 24380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_265
timestamp 1688980957
transform 1 0 25484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_277
timestamp 1688980957
transform 1 0 26588 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 1688980957
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 1688980957
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_317
timestamp 1688980957
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_329
timestamp 1688980957
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_335
timestamp 1688980957
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_337
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_349
timestamp 1688980957
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_361
timestamp 1688980957
transform 1 0 34316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_393
timestamp 1688980957
transform 1 0 37260 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_9
timestamp 1688980957
transform 1 0 1932 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_25
timestamp 1688980957
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_33
timestamp 1688980957
transform 1 0 4140 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_37
timestamp 1688980957
transform 1 0 4508 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_49
timestamp 1688980957
transform 1 0 5612 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_61
timestamp 1688980957
transform 1 0 6716 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_73
timestamp 1688980957
transform 1 0 7820 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_81
timestamp 1688980957
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1688980957
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_109
timestamp 1688980957
transform 1 0 11132 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_115
timestamp 1688980957
transform 1 0 11684 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_122
timestamp 1688980957
transform 1 0 12328 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_126
timestamp 1688980957
transform 1 0 12696 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_138
timestamp 1688980957
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 1688980957
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 1688980957
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 1688980957
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 1688980957
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1688980957
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_209
timestamp 1688980957
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_235
timestamp 1688980957
transform 1 0 22724 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_247
timestamp 1688980957
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1688980957
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 1688980957
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_277
timestamp 1688980957
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_289
timestamp 1688980957
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 1688980957
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1688980957
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_321
timestamp 1688980957
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_333
timestamp 1688980957
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_345
timestamp 1688980957
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_357
timestamp 1688980957
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_363
timestamp 1688980957
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_365
timestamp 1688980957
transform 1 0 34684 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_370
timestamp 1688980957
transform 1 0 35144 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_389
timestamp 1688980957
transform 1 0 36892 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_395
timestamp 1688980957
transform 1 0 37444 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_9
timestamp 1688980957
transform 1 0 1932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_27
timestamp 1688980957
transform 1 0 3588 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_35
timestamp 1688980957
transform 1 0 4324 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1688980957
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1688980957
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1688980957
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1688980957
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1688980957
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1688980957
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1688980957
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_125
timestamp 1688980957
transform 1 0 12604 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_133
timestamp 1688980957
transform 1 0 13340 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 1688980957
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1688980957
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1688980957
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1688980957
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1688980957
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 1688980957
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_205
timestamp 1688980957
transform 1 0 19964 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1688980957
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_241
timestamp 1688980957
transform 1 0 23276 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_245
timestamp 1688980957
transform 1 0 23644 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_257
timestamp 1688980957
transform 1 0 24748 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_269
timestamp 1688980957
transform 1 0 25852 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_277
timestamp 1688980957
transform 1 0 26588 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1688980957
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 1688980957
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_317
timestamp 1688980957
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_329
timestamp 1688980957
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_335
timestamp 1688980957
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_337
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_349
timestamp 1688980957
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_361
timestamp 1688980957
transform 1 0 34316 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_389
timestamp 1688980957
transform 1 0 36892 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_393
timestamp 1688980957
transform 1 0 37260 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_37
timestamp 1688980957
transform 1 0 4508 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_55
timestamp 1688980957
transform 1 0 6164 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_67
timestamp 1688980957
transform 1 0 7268 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_79
timestamp 1688980957
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1688980957
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1688980957
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1688980957
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1688980957
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1688980957
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_153
timestamp 1688980957
transform 1 0 15180 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_172
timestamp 1688980957
transform 1 0 16928 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_184
timestamp 1688980957
transform 1 0 18032 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_205
timestamp 1688980957
transform 1 0 19964 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_215
timestamp 1688980957
transform 1 0 20884 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_223
timestamp 1688980957
transform 1 0 21620 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_227
timestamp 1688980957
transform 1 0 21988 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_231
timestamp 1688980957
transform 1 0 22356 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_243
timestamp 1688980957
transform 1 0 23460 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1688980957
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 1688980957
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 1688980957
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 1688980957
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 1688980957
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 1688980957
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1688980957
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_321
timestamp 1688980957
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_333
timestamp 1688980957
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_345
timestamp 1688980957
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_357
timestamp 1688980957
transform 1 0 33948 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_361
timestamp 1688980957
transform 1 0 34316 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_365
timestamp 1688980957
transform 1 0 34684 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_9
timestamp 1688980957
transform 1 0 1932 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_43
timestamp 1688980957
transform 1 0 5060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1688980957
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 1688980957
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 1688980957
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 1688980957
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1688980957
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1688980957
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 1688980957
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 1688980957
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 1688980957
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1688980957
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 1688980957
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_193
timestamp 1688980957
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_205
timestamp 1688980957
transform 1 0 19964 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_213
timestamp 1688980957
transform 1 0 20700 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 1688980957
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1688980957
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 1688980957
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 1688980957
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_261
timestamp 1688980957
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 1688980957
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1688980957
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 1688980957
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 1688980957
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_317
timestamp 1688980957
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_329
timestamp 1688980957
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_335
timestamp 1688980957
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_337
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_349
timestamp 1688980957
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_361
timestamp 1688980957
transform 1 0 34316 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_367
timestamp 1688980957
transform 1 0 34868 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_385
timestamp 1688980957
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_391
timestamp 1688980957
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_393
timestamp 1688980957
transform 1 0 37260 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_37
timestamp 1688980957
transform 1 0 4508 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_49
timestamp 1688980957
transform 1 0 5612 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_61
timestamp 1688980957
transform 1 0 6716 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_69
timestamp 1688980957
transform 1 0 7452 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_78
timestamp 1688980957
transform 1 0 8280 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1688980957
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1688980957
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1688980957
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1688980957
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1688980957
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1688980957
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 1688980957
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 1688980957
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 1688980957
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1688980957
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 1688980957
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 1688980957
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_233
timestamp 1688980957
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 1688980957
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1688980957
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 1688980957
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_277
timestamp 1688980957
transform 1 0 26588 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_281
timestamp 1688980957
transform 1 0 26956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_288
timestamp 1688980957
transform 1 0 27600 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_292
timestamp 1688980957
transform 1 0 27968 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_304
timestamp 1688980957
transform 1 0 29072 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_321
timestamp 1688980957
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_333
timestamp 1688980957
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_345
timestamp 1688980957
transform 1 0 32844 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_353
timestamp 1688980957
transform 1 0 33580 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_389
timestamp 1688980957
transform 1 0 36892 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_395
timestamp 1688980957
transform 1 0 37444 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_34
timestamp 1688980957
transform 1 0 4232 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_38
timestamp 1688980957
transform 1 0 4600 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_50
timestamp 1688980957
transform 1 0 5704 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1688980957
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1688980957
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 1688980957
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 1688980957
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1688980957
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1688980957
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1688980957
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 1688980957
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 1688980957
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1688980957
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1688980957
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_193
timestamp 1688980957
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 1688980957
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 1688980957
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1688980957
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_233
timestamp 1688980957
transform 1 0 22540 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_245
timestamp 1688980957
transform 1 0 23644 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_251
timestamp 1688980957
transform 1 0 24196 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_263
timestamp 1688980957
transform 1 0 25300 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_275
timestamp 1688980957
transform 1 0 26404 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1688980957
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1688980957
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 1688980957
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_317
timestamp 1688980957
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_329
timestamp 1688980957
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 1688980957
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_337
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_349
timestamp 1688980957
transform 1 0 33212 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_357
timestamp 1688980957
transform 1 0 33948 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_385
timestamp 1688980957
transform 1 0 36524 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_389
timestamp 1688980957
transform 1 0 36892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_393
timestamp 1688980957
transform 1 0 37260 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_25
timestamp 1688980957
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_37
timestamp 1688980957
transform 1 0 4508 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_49
timestamp 1688980957
transform 1 0 5612 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_61
timestamp 1688980957
transform 1 0 6716 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_73
timestamp 1688980957
transform 1 0 7820 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_81
timestamp 1688980957
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1688980957
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1688980957
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 1688980957
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 1688980957
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1688980957
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1688980957
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 1688980957
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 1688980957
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 1688980957
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1688980957
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 1688980957
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 1688980957
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 1688980957
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 1688980957
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1688980957
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1688980957
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 1688980957
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 1688980957
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_301
timestamp 1688980957
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1688980957
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_321
timestamp 1688980957
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_333
timestamp 1688980957
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_345
timestamp 1688980957
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_357
timestamp 1688980957
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_363
timestamp 1688980957
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_395
timestamp 1688980957
transform 1 0 37444 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_31
timestamp 1688980957
transform 1 0 3956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_43
timestamp 1688980957
transform 1 0 5060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1688980957
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1688980957
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1688980957
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 1688980957
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1688980957
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1688980957
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1688980957
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1688980957
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 1688980957
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 1688980957
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1688980957
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 1688980957
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_193
timestamp 1688980957
transform 1 0 18860 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_201
timestamp 1688980957
transform 1 0 19596 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1688980957
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 1688980957
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 1688980957
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 1688980957
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1688980957
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_289
timestamp 1688980957
transform 1 0 27692 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_301
timestamp 1688980957
transform 1 0 28796 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_313
timestamp 1688980957
transform 1 0 29900 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_325
timestamp 1688980957
transform 1 0 31004 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_333
timestamp 1688980957
transform 1 0 31740 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_337
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_349
timestamp 1688980957
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_361
timestamp 1688980957
transform 1 0 34316 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_367
timestamp 1688980957
transform 1 0 34868 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_393
timestamp 1688980957
transform 1 0 37260 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1688980957
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1688980957
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1688980957
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1688980957
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1688980957
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1688980957
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1688980957
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1688980957
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1688980957
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1688980957
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1688980957
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 1688980957
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 1688980957
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 1688980957
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1688980957
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1688980957
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1688980957
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 1688980957
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 1688980957
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1688980957
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_269
timestamp 1688980957
transform 1 0 25852 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_273
timestamp 1688980957
transform 1 0 26220 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_285
timestamp 1688980957
transform 1 0 27324 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_297
timestamp 1688980957
transform 1 0 28428 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_305
timestamp 1688980957
transform 1 0 29164 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 1688980957
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_321
timestamp 1688980957
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_333
timestamp 1688980957
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_345
timestamp 1688980957
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_357
timestamp 1688980957
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_363
timestamp 1688980957
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_365
timestamp 1688980957
transform 1 0 34684 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_371
timestamp 1688980957
transform 1 0 35236 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_33
timestamp 1688980957
transform 1 0 4140 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_45
timestamp 1688980957
transform 1 0 5244 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_53
timestamp 1688980957
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1688980957
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 1688980957
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 1688980957
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_105
timestamp 1688980957
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1688980957
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_137
timestamp 1688980957
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_149
timestamp 1688980957
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_161
timestamp 1688980957
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1688980957
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 1688980957
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_193
timestamp 1688980957
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_205
timestamp 1688980957
transform 1 0 19964 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_214
timestamp 1688980957
transform 1 0 20792 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_218
timestamp 1688980957
transform 1 0 21160 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 1688980957
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_249
timestamp 1688980957
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_261
timestamp 1688980957
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_273
timestamp 1688980957
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 1688980957
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 1688980957
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_305
timestamp 1688980957
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_317
timestamp 1688980957
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_329
timestamp 1688980957
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_335
timestamp 1688980957
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_337
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_349
timestamp 1688980957
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_361
timestamp 1688980957
transform 1 0 34316 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_367
timestamp 1688980957
transform 1 0 34868 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_385
timestamp 1688980957
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_391
timestamp 1688980957
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_393
timestamp 1688980957
transform 1 0 37260 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_9
timestamp 1688980957
transform 1 0 1932 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_43
timestamp 1688980957
transform 1 0 5060 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_55
timestamp 1688980957
transform 1 0 6164 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_67
timestamp 1688980957
transform 1 0 7268 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_79
timestamp 1688980957
transform 1 0 8372 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1688980957
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_97
timestamp 1688980957
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_109
timestamp 1688980957
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_121
timestamp 1688980957
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_133
timestamp 1688980957
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1688980957
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_153
timestamp 1688980957
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_165
timestamp 1688980957
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_177
timestamp 1688980957
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_189
timestamp 1688980957
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1688980957
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_209
timestamp 1688980957
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_221
timestamp 1688980957
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_233
timestamp 1688980957
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_245
timestamp 1688980957
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 1688980957
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_265
timestamp 1688980957
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_277
timestamp 1688980957
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_289
timestamp 1688980957
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_301
timestamp 1688980957
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_307
timestamp 1688980957
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_309
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_321
timestamp 1688980957
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_333
timestamp 1688980957
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_345
timestamp 1688980957
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_357
timestamp 1688980957
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_363
timestamp 1688980957
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_389
timestamp 1688980957
transform 1 0 36892 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_395
timestamp 1688980957
transform 1 0 37444 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_9
timestamp 1688980957
transform 1 0 1932 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_33
timestamp 1688980957
transform 1 0 4140 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_45
timestamp 1688980957
transform 1 0 5244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_53
timestamp 1688980957
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1688980957
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_81
timestamp 1688980957
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_93
timestamp 1688980957
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_105
timestamp 1688980957
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1688980957
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 1688980957
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_137
timestamp 1688980957
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_149
timestamp 1688980957
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_161
timestamp 1688980957
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1688980957
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_181
timestamp 1688980957
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_193
timestamp 1688980957
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_205
timestamp 1688980957
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_217
timestamp 1688980957
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1688980957
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_237
timestamp 1688980957
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_249
timestamp 1688980957
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_261
timestamp 1688980957
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_273
timestamp 1688980957
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 1688980957
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_293
timestamp 1688980957
transform 1 0 28060 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_311
timestamp 1688980957
transform 1 0 29716 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_315
timestamp 1688980957
transform 1 0 30084 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_327
timestamp 1688980957
transform 1 0 31188 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_335
timestamp 1688980957
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_337
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_349
timestamp 1688980957
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_361
timestamp 1688980957
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_373
timestamp 1688980957
transform 1 0 35420 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_393
timestamp 1688980957
transform 1 0 37260 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_25
timestamp 1688980957
transform 1 0 3404 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_37
timestamp 1688980957
transform 1 0 4508 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_49
timestamp 1688980957
transform 1 0 5612 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_61
timestamp 1688980957
transform 1 0 6716 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_73
timestamp 1688980957
transform 1 0 7820 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_81
timestamp 1688980957
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 1688980957
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 1688980957
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 1688980957
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 1688980957
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1688980957
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_153
timestamp 1688980957
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_165
timestamp 1688980957
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_177
timestamp 1688980957
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_189
timestamp 1688980957
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1688980957
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_214
timestamp 1688980957
transform 1 0 20792 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_218
timestamp 1688980957
transform 1 0 21160 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_230
timestamp 1688980957
transform 1 0 22264 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_242
timestamp 1688980957
transform 1 0 23368 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_250
timestamp 1688980957
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_265
timestamp 1688980957
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_277
timestamp 1688980957
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_289
timestamp 1688980957
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_301
timestamp 1688980957
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 1688980957
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 1688980957
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_321
timestamp 1688980957
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_333
timestamp 1688980957
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_345
timestamp 1688980957
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_357
timestamp 1688980957
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_363
timestamp 1688980957
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_365
timestamp 1688980957
transform 1 0 34684 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_373
timestamp 1688980957
transform 1 0 35420 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_389
timestamp 1688980957
transform 1 0 36892 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_395
timestamp 1688980957
transform 1 0 37444 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_33
timestamp 1688980957
transform 1 0 4140 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_45
timestamp 1688980957
transform 1 0 5244 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_53
timestamp 1688980957
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 1688980957
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_81
timestamp 1688980957
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_93
timestamp 1688980957
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_105
timestamp 1688980957
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1688980957
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_125
timestamp 1688980957
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_137
timestamp 1688980957
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_149
timestamp 1688980957
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_161
timestamp 1688980957
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1688980957
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_181
timestamp 1688980957
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_193
timestamp 1688980957
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_205
timestamp 1688980957
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_217
timestamp 1688980957
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1688980957
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_237
timestamp 1688980957
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_249
timestamp 1688980957
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_261
timestamp 1688980957
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_273
timestamp 1688980957
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1688980957
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_293
timestamp 1688980957
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_305
timestamp 1688980957
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_317
timestamp 1688980957
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_329
timestamp 1688980957
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_335
timestamp 1688980957
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_337
timestamp 1688980957
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_349
timestamp 1688980957
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_361
timestamp 1688980957
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_373
timestamp 1688980957
transform 1 0 35420 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_379
timestamp 1688980957
transform 1 0 35972 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_382
timestamp 1688980957
transform 1 0 36248 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_393
timestamp 1688980957
transform 1 0 37260 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_9
timestamp 1688980957
transform 1 0 1932 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1688980957
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 1688980957
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 1688980957
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1688980957
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_97
timestamp 1688980957
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_109
timestamp 1688980957
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_121
timestamp 1688980957
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_133
timestamp 1688980957
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1688980957
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_153
timestamp 1688980957
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_165
timestamp 1688980957
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_177
timestamp 1688980957
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_189
timestamp 1688980957
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 1688980957
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_209
timestamp 1688980957
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_221
timestamp 1688980957
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_233
timestamp 1688980957
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_245
timestamp 1688980957
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 1688980957
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_265
timestamp 1688980957
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_277
timestamp 1688980957
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_289
timestamp 1688980957
transform 1 0 27692 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_295
timestamp 1688980957
transform 1 0 28244 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_304
timestamp 1688980957
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_321
timestamp 1688980957
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_333
timestamp 1688980957
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_345
timestamp 1688980957
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_357
timestamp 1688980957
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_363
timestamp 1688980957
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_365
timestamp 1688980957
transform 1 0 34684 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_371
timestamp 1688980957
transform 1 0 35236 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_389
timestamp 1688980957
transform 1 0 36892 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_395
timestamp 1688980957
transform 1 0 37444 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_41
timestamp 1688980957
transform 1 0 4876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_53
timestamp 1688980957
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 1688980957
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_81
timestamp 1688980957
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_93
timestamp 1688980957
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_105
timestamp 1688980957
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1688980957
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 1688980957
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_137
timestamp 1688980957
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_149
timestamp 1688980957
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 1688980957
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1688980957
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 1688980957
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_193
timestamp 1688980957
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_205
timestamp 1688980957
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_217
timestamp 1688980957
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1688980957
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_237
timestamp 1688980957
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_249
timestamp 1688980957
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_261
timestamp 1688980957
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_273
timestamp 1688980957
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1688980957
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_293
timestamp 1688980957
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_305
timestamp 1688980957
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_317
timestamp 1688980957
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_329
timestamp 1688980957
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_335
timestamp 1688980957
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_337
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_349
timestamp 1688980957
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_361
timestamp 1688980957
transform 1 0 34316 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_389
timestamp 1688980957
transform 1 0 36892 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_393
timestamp 1688980957
transform 1 0 37260 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_25
timestamp 1688980957
transform 1 0 3404 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_37
timestamp 1688980957
transform 1 0 4508 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_49
timestamp 1688980957
transform 1 0 5612 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_61
timestamp 1688980957
transform 1 0 6716 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_73
timestamp 1688980957
transform 1 0 7820 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_81
timestamp 1688980957
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 1688980957
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 1688980957
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_121
timestamp 1688980957
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_133
timestamp 1688980957
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1688980957
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_153
timestamp 1688980957
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_165
timestamp 1688980957
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_177
timestamp 1688980957
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_189
timestamp 1688980957
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1688980957
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_209
timestamp 1688980957
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_221
timestamp 1688980957
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_233
timestamp 1688980957
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_245
timestamp 1688980957
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 1688980957
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_265
timestamp 1688980957
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_277
timestamp 1688980957
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_289
timestamp 1688980957
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_301
timestamp 1688980957
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_307
timestamp 1688980957
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 1688980957
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_321
timestamp 1688980957
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_333
timestamp 1688980957
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_345
timestamp 1688980957
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_357
timestamp 1688980957
transform 1 0 33948 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_361
timestamp 1688980957
transform 1 0 34316 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_365
timestamp 1688980957
transform 1 0 34684 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_19
timestamp 1688980957
transform 1 0 2852 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_25
timestamp 1688980957
transform 1 0 3404 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_41
timestamp 1688980957
transform 1 0 4876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_53
timestamp 1688980957
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 1688980957
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 1688980957
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_105
timestamp 1688980957
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_125
timestamp 1688980957
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_137
timestamp 1688980957
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_149
timestamp 1688980957
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_161
timestamp 1688980957
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1688980957
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_181
timestamp 1688980957
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_193
timestamp 1688980957
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_205
timestamp 1688980957
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_217
timestamp 1688980957
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1688980957
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 1688980957
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 1688980957
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_261
timestamp 1688980957
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_273
timestamp 1688980957
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 1688980957
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_293
timestamp 1688980957
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_305
timestamp 1688980957
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_317
timestamp 1688980957
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_329
timestamp 1688980957
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_335
timestamp 1688980957
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_349
timestamp 1688980957
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_361
timestamp 1688980957
transform 1 0 34316 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_367
timestamp 1688980957
transform 1 0 34868 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_385
timestamp 1688980957
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_391
timestamp 1688980957
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_393
timestamp 1688980957
transform 1 0 37260 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_25
timestamp 1688980957
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_37
timestamp 1688980957
transform 1 0 4508 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_49
timestamp 1688980957
transform 1 0 5612 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_61
timestamp 1688980957
transform 1 0 6716 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_73
timestamp 1688980957
transform 1 0 7820 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_81
timestamp 1688980957
transform 1 0 8556 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 1688980957
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_109
timestamp 1688980957
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_121
timestamp 1688980957
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_133
timestamp 1688980957
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1688980957
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_153
timestamp 1688980957
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_165
timestamp 1688980957
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_177
timestamp 1688980957
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_189
timestamp 1688980957
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1688980957
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_209
timestamp 1688980957
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_221
timestamp 1688980957
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_233
timestamp 1688980957
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_245
timestamp 1688980957
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1688980957
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 1688980957
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_277
timestamp 1688980957
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_289
timestamp 1688980957
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_301
timestamp 1688980957
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_307
timestamp 1688980957
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_309
timestamp 1688980957
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_321
timestamp 1688980957
transform 1 0 30636 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_332
timestamp 1688980957
transform 1 0 31648 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_344
timestamp 1688980957
transform 1 0 32752 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_356
timestamp 1688980957
transform 1 0 33856 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_389
timestamp 1688980957
transform 1 0 36892 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_395
timestamp 1688980957
transform 1 0 37444 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_47
timestamp 1688980957
transform 1 0 5428 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_93
timestamp 1688980957
transform 1 0 9660 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_97
timestamp 1688980957
transform 1 0 10028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_109
timestamp 1688980957
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 1688980957
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 1688980957
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 1688980957
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 1688980957
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_181
timestamp 1688980957
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_193
timestamp 1688980957
transform 1 0 18860 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_201
timestamp 1688980957
transform 1 0 19596 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_210
timestamp 1688980957
transform 1 0 20424 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_222
timestamp 1688980957
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 1688980957
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_249
timestamp 1688980957
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_261
timestamp 1688980957
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_273
timestamp 1688980957
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1688980957
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 1688980957
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_305
timestamp 1688980957
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_317
timestamp 1688980957
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_329
timestamp 1688980957
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_335
timestamp 1688980957
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_337
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_349
timestamp 1688980957
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_361
timestamp 1688980957
transform 1 0 34316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_393
timestamp 1688980957
transform 1 0 37260 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_25
timestamp 1688980957
transform 1 0 3404 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_42
timestamp 1688980957
transform 1 0 4968 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_65
timestamp 1688980957
transform 1 0 7084 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_69
timestamp 1688980957
transform 1 0 7452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_81
timestamp 1688980957
transform 1 0 8556 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1688980957
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_109
timestamp 1688980957
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_121
timestamp 1688980957
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_133
timestamp 1688980957
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 1688980957
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 1688980957
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_165
timestamp 1688980957
transform 1 0 16284 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_173
timestamp 1688980957
transform 1 0 17020 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_178
timestamp 1688980957
transform 1 0 17480 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_190
timestamp 1688980957
transform 1 0 18584 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_209
timestamp 1688980957
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_221
timestamp 1688980957
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_233
timestamp 1688980957
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_245
timestamp 1688980957
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 1688980957
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 1688980957
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 1688980957
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_289
timestamp 1688980957
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_301
timestamp 1688980957
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 1688980957
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_309
timestamp 1688980957
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_321
timestamp 1688980957
transform 1 0 30636 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_331
timestamp 1688980957
transform 1 0 31556 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_343
timestamp 1688980957
transform 1 0 32660 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_355
timestamp 1688980957
transform 1 0 33764 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_363
timestamp 1688980957
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_365
timestamp 1688980957
transform 1 0 34684 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_370
timestamp 1688980957
transform 1 0 35144 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_389
timestamp 1688980957
transform 1 0 36892 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_395
timestamp 1688980957
transform 1 0 37444 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_49
timestamp 1688980957
transform 1 0 5612 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 1688980957
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 1688980957
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_125
timestamp 1688980957
transform 1 0 12604 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_133
timestamp 1688980957
transform 1 0 13340 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_150
timestamp 1688980957
transform 1 0 14904 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_162
timestamp 1688980957
transform 1 0 16008 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_180
timestamp 1688980957
transform 1 0 17664 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_184
timestamp 1688980957
transform 1 0 18032 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_196
timestamp 1688980957
transform 1 0 19136 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_208
timestamp 1688980957
transform 1 0 20240 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_220
timestamp 1688980957
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 1688980957
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 1688980957
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 1688980957
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_273
timestamp 1688980957
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 1688980957
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_293
timestamp 1688980957
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_305
timestamp 1688980957
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_317
timestamp 1688980957
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_329
timestamp 1688980957
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 1688980957
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_337
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_349
timestamp 1688980957
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_361
timestamp 1688980957
transform 1 0 34316 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_389
timestamp 1688980957
transform 1 0 36892 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_393
timestamp 1688980957
transform 1 0 37260 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_9
timestamp 1688980957
transform 1 0 1932 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_43
timestamp 1688980957
transform 1 0 5060 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_55
timestamp 1688980957
transform 1 0 6164 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_67
timestamp 1688980957
transform 1 0 7268 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_79
timestamp 1688980957
transform 1 0 8372 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1688980957
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1688980957
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 1688980957
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_121
timestamp 1688980957
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 1688980957
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 1688980957
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_153
timestamp 1688980957
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_165
timestamp 1688980957
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_177
timestamp 1688980957
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_189
timestamp 1688980957
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 1688980957
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 1688980957
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_221
timestamp 1688980957
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_233
timestamp 1688980957
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_245
timestamp 1688980957
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 1688980957
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 1688980957
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_277
timestamp 1688980957
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_289
timestamp 1688980957
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_301
timestamp 1688980957
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_307
timestamp 1688980957
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 1688980957
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_321
timestamp 1688980957
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_333
timestamp 1688980957
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_345
timestamp 1688980957
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_357
timestamp 1688980957
transform 1 0 33948 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_361
timestamp 1688980957
transform 1 0 34316 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_365
timestamp 1688980957
transform 1 0 34684 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_19
timestamp 1688980957
transform 1 0 2852 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_25
timestamp 1688980957
transform 1 0 3404 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_35
timestamp 1688980957
transform 1 0 4324 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_47
timestamp 1688980957
transform 1 0 5428 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1688980957
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 1688980957
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_81
timestamp 1688980957
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_93
timestamp 1688980957
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_105
timestamp 1688980957
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1688980957
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_125
timestamp 1688980957
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_137
timestamp 1688980957
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_149
timestamp 1688980957
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_161
timestamp 1688980957
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1688980957
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_181
timestamp 1688980957
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_193
timestamp 1688980957
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_205
timestamp 1688980957
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_217
timestamp 1688980957
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 1688980957
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_225
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_237
timestamp 1688980957
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_249
timestamp 1688980957
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_261
timestamp 1688980957
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_273
timestamp 1688980957
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 1688980957
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 1688980957
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 1688980957
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_317
timestamp 1688980957
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_329
timestamp 1688980957
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_335
timestamp 1688980957
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_337
timestamp 1688980957
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_349
timestamp 1688980957
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_361
timestamp 1688980957
transform 1 0 34316 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_367
timestamp 1688980957
transform 1 0 34868 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_385
timestamp 1688980957
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_391
timestamp 1688980957
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_393
timestamp 1688980957
transform 1 0 37260 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_25
timestamp 1688980957
transform 1 0 3404 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_37
timestamp 1688980957
transform 1 0 4508 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_49
timestamp 1688980957
transform 1 0 5612 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_61
timestamp 1688980957
transform 1 0 6716 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_73
timestamp 1688980957
transform 1 0 7820 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_81
timestamp 1688980957
transform 1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_97
timestamp 1688980957
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_109
timestamp 1688980957
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_121
timestamp 1688980957
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_133
timestamp 1688980957
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1688980957
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 1688980957
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_165
timestamp 1688980957
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_177
timestamp 1688980957
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_189
timestamp 1688980957
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 1688980957
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_205
timestamp 1688980957
transform 1 0 19964 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_217
timestamp 1688980957
transform 1 0 21068 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_229
timestamp 1688980957
transform 1 0 22172 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_241
timestamp 1688980957
transform 1 0 23276 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_249
timestamp 1688980957
transform 1 0 24012 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 1688980957
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 1688980957
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_277
timestamp 1688980957
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_289
timestamp 1688980957
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_301
timestamp 1688980957
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 1688980957
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 1688980957
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_321
timestamp 1688980957
transform 1 0 30636 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_347
timestamp 1688980957
transform 1 0 33028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_359
timestamp 1688980957
transform 1 0 34132 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_363
timestamp 1688980957
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_389
timestamp 1688980957
transform 1 0 36892 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_395
timestamp 1688980957
transform 1 0 37444 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_47
timestamp 1688980957
transform 1 0 5428 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1688980957
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 1688980957
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_81
timestamp 1688980957
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_93
timestamp 1688980957
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_105
timestamp 1688980957
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_111
timestamp 1688980957
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_125
timestamp 1688980957
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_137
timestamp 1688980957
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_149
timestamp 1688980957
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_161
timestamp 1688980957
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 1688980957
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_181
timestamp 1688980957
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_193
timestamp 1688980957
transform 1 0 18860 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_201
timestamp 1688980957
transform 1 0 19596 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_212
timestamp 1688980957
transform 1 0 20608 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_225
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_237
timestamp 1688980957
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_249
timestamp 1688980957
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_261
timestamp 1688980957
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_273
timestamp 1688980957
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 1688980957
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_293
timestamp 1688980957
transform 1 0 28060 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_319
timestamp 1688980957
transform 1 0 30452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_331
timestamp 1688980957
transform 1 0 31556 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_335
timestamp 1688980957
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_345
timestamp 1688980957
transform 1 0 32844 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_357
timestamp 1688980957
transform 1 0 33948 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_361
timestamp 1688980957
transform 1 0 34316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_393
timestamp 1688980957
transform 1 0 37260 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_25
timestamp 1688980957
transform 1 0 3404 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_37
timestamp 1688980957
transform 1 0 4508 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_49
timestamp 1688980957
transform 1 0 5612 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_55
timestamp 1688980957
transform 1 0 6164 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_64
timestamp 1688980957
transform 1 0 6992 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_76
timestamp 1688980957
transform 1 0 8096 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_97
timestamp 1688980957
transform 1 0 10028 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_105
timestamp 1688980957
transform 1 0 10764 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_114
timestamp 1688980957
transform 1 0 11592 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_126
timestamp 1688980957
transform 1 0 12696 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_138
timestamp 1688980957
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_153
timestamp 1688980957
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_165
timestamp 1688980957
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_177
timestamp 1688980957
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_189
timestamp 1688980957
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 1688980957
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_209
timestamp 1688980957
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_221
timestamp 1688980957
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_233
timestamp 1688980957
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_245
timestamp 1688980957
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_251
timestamp 1688980957
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_265
timestamp 1688980957
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 1688980957
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_289
timestamp 1688980957
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_301
timestamp 1688980957
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 1688980957
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 1688980957
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_321
timestamp 1688980957
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_333
timestamp 1688980957
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_345
timestamp 1688980957
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_357
timestamp 1688980957
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_363
timestamp 1688980957
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_365
timestamp 1688980957
transform 1 0 34684 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_370
timestamp 1688980957
transform 1 0 35144 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_389
timestamp 1688980957
transform 1 0 36892 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_393
timestamp 1688980957
transform 1 0 37260 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_33
timestamp 1688980957
transform 1 0 4140 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_45
timestamp 1688980957
transform 1 0 5244 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_53
timestamp 1688980957
transform 1 0 5980 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 1688980957
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 1688980957
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_93
timestamp 1688980957
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_105
timestamp 1688980957
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 1688980957
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_125
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_137
timestamp 1688980957
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 1688980957
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_161
timestamp 1688980957
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 1688980957
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_181
timestamp 1688980957
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_193
timestamp 1688980957
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_205
timestamp 1688980957
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_217
timestamp 1688980957
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 1688980957
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_237
timestamp 1688980957
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_249
timestamp 1688980957
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_261
timestamp 1688980957
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_273
timestamp 1688980957
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 1688980957
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1688980957
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 1688980957
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_305
timestamp 1688980957
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_317
timestamp 1688980957
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_329
timestamp 1688980957
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 1688980957
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_337
timestamp 1688980957
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_349
timestamp 1688980957
transform 1 0 33212 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_389
timestamp 1688980957
transform 1 0 36892 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_393
timestamp 1688980957
transform 1 0 37260 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_3
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_9
timestamp 1688980957
transform 1 0 1932 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1688980957
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_43
timestamp 1688980957
transform 1 0 5060 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_55
timestamp 1688980957
transform 1 0 6164 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_67
timestamp 1688980957
transform 1 0 7268 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_79
timestamp 1688980957
transform 1 0 8372 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1688980957
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_97
timestamp 1688980957
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_109
timestamp 1688980957
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_121
timestamp 1688980957
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_133
timestamp 1688980957
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 1688980957
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_153
timestamp 1688980957
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_165
timestamp 1688980957
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_177
timestamp 1688980957
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_189
timestamp 1688980957
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_195
timestamp 1688980957
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_209
timestamp 1688980957
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_221
timestamp 1688980957
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_233
timestamp 1688980957
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_245
timestamp 1688980957
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 1688980957
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_253
timestamp 1688980957
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_265
timestamp 1688980957
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_277
timestamp 1688980957
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_289
timestamp 1688980957
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_301
timestamp 1688980957
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 1688980957
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 1688980957
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_321
timestamp 1688980957
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_333
timestamp 1688980957
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_345
timestamp 1688980957
transform 1 0 32844 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_365
timestamp 1688980957
transform 1 0 34684 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_35
timestamp 1688980957
transform 1 0 4324 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_47
timestamp 1688980957
transform 1 0 5428 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1688980957
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 1688980957
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_81
timestamp 1688980957
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_93
timestamp 1688980957
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_105
timestamp 1688980957
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 1688980957
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 1688980957
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_137
timestamp 1688980957
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_149
timestamp 1688980957
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_161
timestamp 1688980957
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 1688980957
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_181
timestamp 1688980957
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_193
timestamp 1688980957
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_205
timestamp 1688980957
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_217
timestamp 1688980957
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 1688980957
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_225
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_237
timestamp 1688980957
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_249
timestamp 1688980957
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_261
timestamp 1688980957
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_273
timestamp 1688980957
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 1688980957
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_281
timestamp 1688980957
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_293
timestamp 1688980957
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_305
timestamp 1688980957
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_317
timestamp 1688980957
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_329
timestamp 1688980957
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 1688980957
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_337
timestamp 1688980957
transform 1 0 32108 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_343
timestamp 1688980957
transform 1 0 32660 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_385
timestamp 1688980957
transform 1 0 36524 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_389
timestamp 1688980957
transform 1 0 36892 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_393
timestamp 1688980957
transform 1 0 37260 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_9
timestamp 1688980957
transform 1 0 1932 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_37
timestamp 1688980957
transform 1 0 4508 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_49
timestamp 1688980957
transform 1 0 5612 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_61
timestamp 1688980957
transform 1 0 6716 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_73
timestamp 1688980957
transform 1 0 7820 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_97
timestamp 1688980957
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_109
timestamp 1688980957
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_121
timestamp 1688980957
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_133
timestamp 1688980957
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 1688980957
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 1688980957
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_165
timestamp 1688980957
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_177
timestamp 1688980957
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_189
timestamp 1688980957
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 1688980957
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_209
timestamp 1688980957
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_221
timestamp 1688980957
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_233
timestamp 1688980957
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_245
timestamp 1688980957
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_251
timestamp 1688980957
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_253
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_265
timestamp 1688980957
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_277
timestamp 1688980957
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_289
timestamp 1688980957
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_301
timestamp 1688980957
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_307
timestamp 1688980957
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_309
timestamp 1688980957
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_321
timestamp 1688980957
transform 1 0 30636 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_346
timestamp 1688980957
transform 1 0 32936 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_395
timestamp 1688980957
transform 1 0 37444 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_43
timestamp 1688980957
transform 1 0 5060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1688980957
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 1688980957
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 1688980957
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_93
timestamp 1688980957
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_105
timestamp 1688980957
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 1688980957
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_125
timestamp 1688980957
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_137
timestamp 1688980957
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_149
timestamp 1688980957
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_161
timestamp 1688980957
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1688980957
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_181
timestamp 1688980957
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_193
timestamp 1688980957
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_205
timestamp 1688980957
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_217
timestamp 1688980957
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 1688980957
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_237
timestamp 1688980957
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_249
timestamp 1688980957
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_261
timestamp 1688980957
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_273
timestamp 1688980957
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 1688980957
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_281
timestamp 1688980957
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_293
timestamp 1688980957
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_305
timestamp 1688980957
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_317
timestamp 1688980957
transform 1 0 30268 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_337
timestamp 1688980957
transform 1 0 32108 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_385
timestamp 1688980957
transform 1 0 36524 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_389
timestamp 1688980957
transform 1 0 36892 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_393
timestamp 1688980957
transform 1 0 37260 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_35
timestamp 1688980957
transform 1 0 4324 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_45
timestamp 1688980957
transform 1 0 5244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_57
timestamp 1688980957
transform 1 0 6348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_69
timestamp 1688980957
transform 1 0 7452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_81
timestamp 1688980957
transform 1 0 8556 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1688980957
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 1688980957
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 1688980957
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 1688980957
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1688980957
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 1688980957
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_165
timestamp 1688980957
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_177
timestamp 1688980957
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_189
timestamp 1688980957
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 1688980957
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_209
timestamp 1688980957
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_221
timestamp 1688980957
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_233
timestamp 1688980957
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 1688980957
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 1688980957
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_265
timestamp 1688980957
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_277
timestamp 1688980957
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_289
timestamp 1688980957
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_301
timestamp 1688980957
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 1688980957
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_309
timestamp 1688980957
transform 1 0 29532 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_365
timestamp 1688980957
transform 1 0 34684 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_9
timestamp 1688980957
transform 1 0 1932 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_35
timestamp 1688980957
transform 1 0 4324 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1688980957
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_63
timestamp 1688980957
transform 1 0 6900 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_75
timestamp 1688980957
transform 1 0 8004 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_87
timestamp 1688980957
transform 1 0 9108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_99
timestamp 1688980957
transform 1 0 10212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 1688980957
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_125
timestamp 1688980957
transform 1 0 12604 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_131
timestamp 1688980957
transform 1 0 13156 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_134
timestamp 1688980957
transform 1 0 13432 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_138
timestamp 1688980957
transform 1 0 13800 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_153
timestamp 1688980957
transform 1 0 15180 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_157
timestamp 1688980957
transform 1 0 15548 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_165
timestamp 1688980957
transform 1 0 16284 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_181
timestamp 1688980957
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_193
timestamp 1688980957
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_205
timestamp 1688980957
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_217
timestamp 1688980957
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_223
timestamp 1688980957
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_225
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_237
timestamp 1688980957
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_249
timestamp 1688980957
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_261
timestamp 1688980957
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_273
timestamp 1688980957
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_279
timestamp 1688980957
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_281
timestamp 1688980957
transform 1 0 26956 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_289
timestamp 1688980957
transform 1 0 27692 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_294
timestamp 1688980957
transform 1 0 28152 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_310
timestamp 1688980957
transform 1 0 29624 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_337
timestamp 1688980957
transform 1 0 32108 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_350
timestamp 1688980957
transform 1 0 33304 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_354
timestamp 1688980957
transform 1 0 33672 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_389
timestamp 1688980957
transform 1 0 36892 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_393
timestamp 1688980957
transform 1 0 37260 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_9
timestamp 1688980957
transform 1 0 1932 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_19
timestamp 1688980957
transform 1 0 2852 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_53
timestamp 1688980957
transform 1 0 5980 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_64
timestamp 1688980957
transform 1 0 6992 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_72
timestamp 1688980957
transform 1 0 7728 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_82
timestamp 1688980957
transform 1 0 8648 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_93
timestamp 1688980957
transform 1 0 9660 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_104
timestamp 1688980957
transform 1 0 10672 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_116
timestamp 1688980957
transform 1 0 11776 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_121
timestamp 1688980957
transform 1 0 12236 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_125
timestamp 1688980957
transform 1 0 12604 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_149
timestamp 1688980957
transform 1 0 14812 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_160
timestamp 1688980957
transform 1 0 15824 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_172
timestamp 1688980957
transform 1 0 16928 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_184
timestamp 1688980957
transform 1 0 18032 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_189
timestamp 1688980957
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 1688980957
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_209
timestamp 1688980957
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_221
timestamp 1688980957
transform 1 0 21436 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_225
timestamp 1688980957
transform 1 0 21804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_232
timestamp 1688980957
transform 1 0 22448 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_236
timestamp 1688980957
transform 1 0 22816 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_240
timestamp 1688980957
transform 1 0 23184 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_253
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_261
timestamp 1688980957
transform 1 0 25116 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_266
timestamp 1688980957
transform 1 0 25576 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_270
timestamp 1688980957
transform 1 0 25944 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_279
timestamp 1688980957
transform 1 0 26772 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_283
timestamp 1688980957
transform 1 0 27140 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_309
timestamp 1688980957
transform 1 0 29532 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_341
timestamp 1688980957
transform 1 0 32476 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_345
timestamp 1688980957
transform 1 0 32844 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_357
timestamp 1688980957
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_363
timestamp 1688980957
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_379
timestamp 1688980957
transform 1 0 35972 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_389
timestamp 1688980957
transform 1 0 36892 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_393
timestamp 1688980957
transform 1 0 37260 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_34
timestamp 1688980957
transform 1 0 4232 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1688980957
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_65
timestamp 1688980957
transform 1 0 7084 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_84
timestamp 1688980957
transform 1 0 8832 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_91
timestamp 1688980957
transform 1 0 9476 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_95
timestamp 1688980957
transform 1 0 9844 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_105
timestamp 1688980957
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 1688980957
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_119
timestamp 1688980957
transform 1 0 12052 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_128
timestamp 1688980957
transform 1 0 12880 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_148
timestamp 1688980957
transform 1 0 14720 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_161
timestamp 1688980957
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 1688980957
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_195
timestamp 1688980957
transform 1 0 19044 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_211
timestamp 1688980957
transform 1 0 20516 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_215
timestamp 1688980957
transform 1 0 20884 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_223
timestamp 1688980957
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_241
timestamp 1688980957
transform 1 0 23276 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_264
timestamp 1688980957
transform 1 0 25392 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 1688980957
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_297
timestamp 1688980957
transform 1 0 28428 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_353
timestamp 1688980957
transform 1 0 33580 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_366
timestamp 1688980957
transform 1 0 34776 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_372
timestamp 1688980957
transform 1 0 35328 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_389
timestamp 1688980957
transform 1 0 36892 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_393
timestamp 1688980957
transform 1 0 37260 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_3
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_25
timestamp 1688980957
transform 1 0 3404 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_35
timestamp 1688980957
transform 1 0 4324 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_136
timestamp 1688980957
transform 1 0 13616 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_187
timestamp 1688980957
transform 1 0 18308 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_213
timestamp 1688980957
transform 1 0 20700 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_217
timestamp 1688980957
transform 1 0 21068 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_234
timestamp 1688980957
transform 1 0 22632 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_253
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_257
timestamp 1688980957
transform 1 0 24748 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_274
timestamp 1688980957
transform 1 0 26312 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_309
timestamp 1688980957
transform 1 0 29532 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_328
timestamp 1688980957
transform 1 0 31280 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_374
timestamp 1688980957
transform 1 0 35512 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_378
timestamp 1688980957
transform 1 0 35880 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_395
timestamp 1688980957
transform 1 0 37444 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_9
timestamp 1688980957
transform 1 0 1932 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_19
timestamp 1688980957
transform 1 0 2852 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_36
timestamp 1688980957
transform 1 0 4416 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_77
timestamp 1688980957
transform 1 0 8188 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_83
timestamp 1688980957
transform 1 0 8740 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_93
timestamp 1688980957
transform 1 0 9660 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_117
timestamp 1688980957
transform 1 0 11868 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_134
timestamp 1688980957
transform 1 0 13432 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_140
timestamp 1688980957
transform 1 0 13984 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_150
timestamp 1688980957
transform 1 0 14904 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_191
timestamp 1688980957
transform 1 0 18676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_197
timestamp 1688980957
transform 1 0 19228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_207
timestamp 1688980957
transform 1 0 20148 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_217
timestamp 1688980957
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1688980957
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_233
timestamp 1688980957
transform 1 0 22540 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_250
timestamp 1688980957
transform 1 0 24104 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_254
timestamp 1688980957
transform 1 0 24472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 1688980957
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_281
timestamp 1688980957
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_285
timestamp 1688980957
transform 1 0 27324 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_295
timestamp 1688980957
transform 1 0 28244 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_299
timestamp 1688980957
transform 1 0 28612 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_327
timestamp 1688980957
transform 1 0 31188 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_331
timestamp 1688980957
transform 1 0 31556 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_335
timestamp 1688980957
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_362
timestamp 1688980957
transform 1 0 34408 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_368
timestamp 1688980957
transform 1 0 34960 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_378
timestamp 1688980957
transform 1 0 35880 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_382
timestamp 1688980957
transform 1 0 36248 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_391
timestamp 1688980957
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_393
timestamp 1688980957
transform 1 0 37260 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_3
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_40
timestamp 1688980957
transform 1 0 4784 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_46
timestamp 1688980957
transform 1 0 5336 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_57
timestamp 1688980957
transform 1 0 6348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_66
timestamp 1688980957
transform 1 0 7176 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_96
timestamp 1688980957
transform 1 0 9936 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_102
timestamp 1688980957
transform 1 0 10488 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_113
timestamp 1688980957
transform 1 0 11500 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_152
timestamp 1688980957
transform 1 0 15088 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_158
timestamp 1688980957
transform 1 0 15640 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_169
timestamp 1688980957
transform 1 0 16652 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_205
timestamp 1688980957
transform 1 0 19964 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_225
timestamp 1688980957
transform 1 0 21804 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_238
timestamp 1688980957
transform 1 0 23000 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_250
timestamp 1688980957
transform 1 0 24104 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_262
timestamp 1688980957
transform 1 0 25208 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_268
timestamp 1688980957
transform 1 0 25760 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_277
timestamp 1688980957
transform 1 0 26588 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_305
timestamp 1688980957
transform 1 0 29164 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_318
timestamp 1688980957
transform 1 0 30360 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_324
timestamp 1688980957
transform 1 0 30912 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_333
timestamp 1688980957
transform 1 0 31740 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_361
timestamp 1688980957
transform 1 0 34316 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_389
timestamp 1688980957
transform 1 0 36892 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_393
timestamp 1688980957
transform 1 0 37260 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3588 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold2 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 2852 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform -1 0 4508 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold4
timestamp 1688980957
transform -1 0 2852 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform -1 0 4140 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold6
timestamp 1688980957
transform -1 0 2852 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform -1 0 4140 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold8
timestamp 1688980957
transform -1 0 2852 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform -1 0 4508 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold10
timestamp 1688980957
transform -1 0 2852 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold12
timestamp 1688980957
transform -1 0 2852 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform 1 0 11408 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold14
timestamp 1688980957
transform 1 0 11960 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform -1 0 18492 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold16
timestamp 1688980957
transform 1 0 17204 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform 1 0 4692 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold18
timestamp 1688980957
transform -1 0 6256 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform -1 0 19136 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold20
timestamp 1688980957
transform -1 0 19136 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform -1 0 9936 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold22
timestamp 1688980957
transform 1 0 9936 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform 1 0 7912 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold24
timestamp 1688980957
transform -1 0 8832 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform -1 0 15824 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold26
timestamp 1688980957
transform 1 0 15088 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform -1 0 26864 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold28
timestamp 1688980957
transform -1 0 26864 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform -1 0 6992 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold30
timestamp 1688980957
transform 1 0 6716 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform -1 0 29624 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold32
timestamp 1688980957
transform -1 0 30544 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform -1 0 14812 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold34
timestamp 1688980957
transform -1 0 13984 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform -1 0 29164 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold36
timestamp 1688980957
transform 1 0 28888 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform -1 0 17388 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold38
timestamp 1688980957
transform 1 0 17664 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform -1 0 15640 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold40
timestamp 1688980957
transform 1 0 15088 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform -1 0 12420 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold42
timestamp 1688980957
transform -1 0 11408 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform 1 0 11776 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold44
timestamp 1688980957
transform 1 0 12512 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1688980957
transform 1 0 36432 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold46
timestamp 1688980957
transform 1 0 36064 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform -1 0 35696 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold48
timestamp 1688980957
transform 1 0 35696 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform -1 0 17388 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold50
timestamp 1688980957
transform 1 0 15088 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform -1 0 29624 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold52
timestamp 1688980957
transform 1 0 32108 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform 1 0 32752 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold54
timestamp 1688980957
transform -1 0 34224 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform 1 0 34960 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold56
timestamp 1688980957
transform 1 0 35696 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform 1 0 10948 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold58
timestamp 1688980957
transform 1 0 9936 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform -1 0 35420 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold60
timestamp 1688980957
transform 1 0 36064 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform 1 0 9200 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold62
timestamp 1688980957
transform -1 0 8832 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform 1 0 29624 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold64
timestamp 1688980957
transform -1 0 32016 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1688980957
transform 1 0 34960 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold66
timestamp 1688980957
transform 1 0 35696 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1688980957
transform -1 0 35420 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold68
timestamp 1688980957
transform 1 0 36064 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform 1 0 33856 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold70
timestamp 1688980957
transform 1 0 36064 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1688980957
transform -1 0 34316 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold72
timestamp 1688980957
transform -1 0 32016 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1688980957
transform 1 0 31096 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold74
timestamp 1688980957
transform -1 0 35696 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1688980957
transform -1 0 35420 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold76
timestamp 1688980957
transform 1 0 35696 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1688980957
transform -1 0 23276 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold78
timestamp 1688980957
transform 1 0 22632 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform 1 0 34684 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold80
timestamp 1688980957
transform 1 0 36064 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1688980957
transform -1 0 19964 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold82
timestamp 1688980957
transform 1 0 19964 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform -1 0 35420 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold84
timestamp 1688980957
transform 1 0 35696 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold86
timestamp 1688980957
transform 1 0 36064 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform -1 0 26772 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold88
timestamp 1688980957
transform 1 0 24564 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform 1 0 34684 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold90
timestamp 1688980957
transform 1 0 36064 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1688980957
transform -1 0 35420 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold92
timestamp 1688980957
transform 1 0 35696 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1688980957
transform -1 0 33120 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold94
timestamp 1688980957
transform 1 0 33580 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1688980957
transform -1 0 35420 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold96
timestamp 1688980957
transform 1 0 36064 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1688980957
transform 1 0 34684 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold98
timestamp 1688980957
transform 1 0 36064 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1688980957
transform -1 0 36892 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold100
timestamp 1688980957
transform -1 0 33580 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1688980957
transform 1 0 33488 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold102
timestamp 1688980957
transform -1 0 33120 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1688980957
transform -1 0 26772 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold104
timestamp 1688980957
transform -1 0 28428 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1688980957
transform -1 0 31740 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold106
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1688980957
transform -1 0 34592 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold108
timestamp 1688980957
transform 1 0 36064 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1688980957
transform -1 0 33120 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold110
timestamp 1688980957
transform -1 0 31648 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1688980957
transform -1 0 35420 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold112
timestamp 1688980957
transform -1 0 34592 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1688980957
transform -1 0 36892 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold114
timestamp 1688980957
transform -1 0 36156 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1688980957
transform 1 0 30544 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold116
timestamp 1688980957
transform 1 0 33120 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1688980957
transform 1 0 2852 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold118
timestamp 1688980957
transform -1 0 2852 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1688980957
transform 1 0 2852 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold120
timestamp 1688980957
transform -1 0 2852 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1688980957
transform -1 0 4876 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold122
timestamp 1688980957
transform -1 0 2852 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1688980957
transform 1 0 33948 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold124
timestamp 1688980957
transform -1 0 31648 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1688980957
transform 1 0 2852 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold126
timestamp 1688980957
transform -1 0 2852 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 1688980957
transform 1 0 4876 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold128
timestamp 1688980957
transform -1 0 2852 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 1688980957
transform 1 0 2852 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold130
timestamp 1688980957
transform -1 0 2852 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 1688980957
transform 1 0 2852 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold132
timestamp 1688980957
transform -1 0 2852 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold134
timestamp 1688980957
transform -1 0 2852 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 1688980957
transform -1 0 33856 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold136
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 1688980957
transform 1 0 2024 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold138
timestamp 1688980957
transform -1 0 3680 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 1688980957
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold140
timestamp 1688980957
transform -1 0 2852 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 1688980957
transform 1 0 2852 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold142
timestamp 1688980957
transform -1 0 2852 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold144
timestamp 1688980957
transform -1 0 2852 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 1688980957
transform -1 0 27692 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold146
timestamp 1688980957
transform 1 0 35696 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold147
timestamp 1688980957
transform -1 0 29624 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold148
timestamp 1688980957
transform -1 0 34592 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold149
timestamp 1688980957
transform 1 0 30820 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold150
timestamp 1688980957
transform -1 0 30544 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  hold151 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  hold152
timestamp 1688980957
transform -1 0 8464 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold153
timestamp 1688980957
transform -1 0 6164 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold154
timestamp 1688980957
transform 1 0 2852 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold155
timestamp 1688980957
transform 1 0 6900 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold156
timestamp 1688980957
transform -1 0 6256 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold157
timestamp 1688980957
transform -1 0 29164 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold158
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold159
timestamp 1688980957
transform 1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold160
timestamp 1688980957
transform -1 0 2852 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold161
timestamp 1688980957
transform -1 0 20608 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold162
timestamp 1688980957
transform 1 0 20240 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold163
timestamp 1688980957
transform -1 0 19964 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold164
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold165
timestamp 1688980957
transform -1 0 8832 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold166
timestamp 1688980957
transform -1 0 4324 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold167
timestamp 1688980957
transform 1 0 4140 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold168
timestamp 1688980957
transform -1 0 2852 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold169
timestamp 1688980957
transform 1 0 32108 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold170
timestamp 1688980957
transform -1 0 35696 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold171
timestamp 1688980957
transform 1 0 2852 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold172
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold173
timestamp 1688980957
transform -1 0 23644 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold174
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold175
timestamp 1688980957
transform -1 0 3588 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold176
timestamp 1688980957
transform -1 0 2852 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold177
timestamp 1688980957
transform 1 0 4048 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold178
timestamp 1688980957
transform 1 0 5244 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold179
timestamp 1688980957
transform -1 0 19964 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold180
timestamp 1688980957
transform 1 0 19228 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold181
timestamp 1688980957
transform 1 0 34684 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold182
timestamp 1688980957
transform 1 0 34960 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold183
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold184
timestamp 1688980957
transform 1 0 23920 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold185
timestamp 1688980957
transform 1 0 34684 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold186
timestamp 1688980957
transform 1 0 31832 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold187
timestamp 1688980957
transform 1 0 28336 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold188
timestamp 1688980957
transform 1 0 33488 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold189
timestamp 1688980957
transform 1 0 17020 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold190
timestamp 1688980957
transform -1 0 17664 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold191
timestamp 1688980957
transform -1 0 12512 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold192
timestamp 1688980957
transform -1 0 12880 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold193
timestamp 1688980957
transform -1 0 34960 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold194
timestamp 1688980957
transform -1 0 36800 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold195
timestamp 1688980957
transform -1 0 35420 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold196
timestamp 1688980957
transform 1 0 34960 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold197
timestamp 1688980957
transform 1 0 30360 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold198
timestamp 1688980957
transform 1 0 33120 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold199
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold200
timestamp 1688980957
transform -1 0 3588 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold201
timestamp 1688980957
transform 1 0 2852 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold202
timestamp 1688980957
transform -1 0 3588 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold203
timestamp 1688980957
transform -1 0 4508 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold204
timestamp 1688980957
transform -1 0 3588 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold205
timestamp 1688980957
transform 1 0 26312 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold206
timestamp 1688980957
transform -1 0 27784 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold207
timestamp 1688980957
transform -1 0 9936 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold208
timestamp 1688980957
transform 1 0 9936 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold209
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold210
timestamp 1688980957
transform -1 0 3588 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold211
timestamp 1688980957
transform -1 0 13248 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold212
timestamp 1688980957
transform -1 0 14812 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold213
timestamp 1688980957
transform 1 0 14352 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold214
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold215
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold216
timestamp 1688980957
transform -1 0 4416 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold217
timestamp 1688980957
transform -1 0 18400 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold218
timestamp 1688980957
transform 1 0 16928 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold219
timestamp 1688980957
transform 1 0 28520 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold220
timestamp 1688980957
transform 1 0 28152 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold221
timestamp 1688980957
transform 1 0 27968 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold222
timestamp 1688980957
transform 1 0 30728 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold223
timestamp 1688980957
transform -1 0 35696 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold224
timestamp 1688980957
transform 1 0 34684 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold225
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold226
timestamp 1688980957
transform -1 0 7176 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold227
timestamp 1688980957
transform -1 0 35696 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold228
timestamp 1688980957
transform 1 0 34684 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold229
timestamp 1688980957
transform -1 0 35696 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold230
timestamp 1688980957
transform 1 0 34960 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold231
timestamp 1688980957
transform -1 0 36064 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold232
timestamp 1688980957
transform 1 0 34684 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold233
timestamp 1688980957
transform -1 0 35696 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold234
timestamp 1688980957
transform 1 0 33856 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold235
timestamp 1688980957
transform -1 0 35696 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold236
timestamp 1688980957
transform 1 0 34960 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold237
timestamp 1688980957
transform -1 0 35696 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold238
timestamp 1688980957
transform 1 0 34960 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold239
timestamp 1688980957
transform -1 0 34592 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold240
timestamp 1688980957
transform 1 0 33120 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold241
timestamp 1688980957
transform -1 0 36064 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold242
timestamp 1688980957
transform 1 0 35328 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold243
timestamp 1688980957
transform 1 0 7360 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold244
timestamp 1688980957
transform 1 0 8096 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold245
timestamp 1688980957
transform -1 0 36064 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold246
timestamp 1688980957
transform 1 0 35328 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold247
timestamp 1688980957
transform 1 0 32476 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold248
timestamp 1688980957
transform 1 0 31648 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold249
timestamp 1688980957
transform 1 0 14352 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold250
timestamp 1688980957
transform 1 0 14996 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold251
timestamp 1688980957
transform -1 0 36064 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold252
timestamp 1688980957
transform 1 0 35328 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold253
timestamp 1688980957
transform -1 0 36064 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold254
timestamp 1688980957
transform 1 0 35328 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold255
timestamp 1688980957
transform -1 0 36064 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold256
timestamp 1688980957
transform 1 0 35328 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold257
timestamp 1688980957
transform 1 0 9936 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold258
timestamp 1688980957
transform -1 0 11408 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold259
timestamp 1688980957
transform 1 0 27692 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold260
timestamp 1688980957
transform 1 0 26956 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold261
timestamp 1688980957
transform -1 0 3588 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold262
timestamp 1688980957
transform -1 0 4508 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold263
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold264
timestamp 1688980957
transform -1 0 3588 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold265
timestamp 1688980957
transform -1 0 34592 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold266
timestamp 1688980957
transform 1 0 30912 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold267
timestamp 1688980957
transform 1 0 16560 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold268
timestamp 1688980957
transform -1 0 16560 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold269
timestamp 1688980957
transform 1 0 13248 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold270
timestamp 1688980957
transform 1 0 13892 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold271
timestamp 1688980957
transform -1 0 4324 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold272
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold273
timestamp 1688980957
transform 1 0 19136 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold274
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold275
timestamp 1688980957
transform -1 0 3588 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold276
timestamp 1688980957
transform -1 0 5060 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold277
timestamp 1688980957
transform -1 0 36892 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold278
timestamp 1688980957
transform -1 0 36892 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold279
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold280
timestamp 1688980957
transform -1 0 3588 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold281
timestamp 1688980957
transform 1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold282
timestamp 1688980957
transform -1 0 5152 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold283
timestamp 1688980957
transform -1 0 3588 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold284
timestamp 1688980957
transform -1 0 4140 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold285
timestamp 1688980957
transform -1 0 12512 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold286
timestamp 1688980957
transform -1 0 13892 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold287
timestamp 1688980957
transform -1 0 4324 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold288
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold289
timestamp 1688980957
transform -1 0 36064 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold290
timestamp 1688980957
transform 1 0 35328 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold291
timestamp 1688980957
transform -1 0 14628 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold292
timestamp 1688980957
transform -1 0 13248 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold293
timestamp 1688980957
transform -1 0 31740 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold294
timestamp 1688980957
transform 1 0 28704 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold295
timestamp 1688980957
transform -1 0 2208 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold296
timestamp 1688980957
transform 1 0 2944 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold297
timestamp 1688980957
transform 1 0 24104 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold298
timestamp 1688980957
transform 1 0 23368 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold299
timestamp 1688980957
transform 1 0 2852 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold300
timestamp 1688980957
transform -1 0 4324 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold301
timestamp 1688980957
transform -1 0 4508 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold302
timestamp 1688980957
transform -1 0 4140 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold303
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold304
timestamp 1688980957
transform 1 0 21804 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold305
timestamp 1688980957
transform -1 0 35420 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold306
timestamp 1688980957
transform 1 0 31280 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold307
timestamp 1688980957
transform 1 0 25484 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold308
timestamp 1688980957
transform 1 0 25852 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold309
timestamp 1688980957
transform 1 0 31280 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold310
timestamp 1688980957
transform -1 0 34316 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold311
timestamp 1688980957
transform -1 0 36064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold312
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold313
timestamp 1688980957
transform -1 0 32200 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold314
timestamp 1688980957
transform 1 0 31280 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold315
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold316
timestamp 1688980957
transform 1 0 30360 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold317
timestamp 1688980957
transform 1 0 29808 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold318
timestamp 1688980957
transform 1 0 30544 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold319
timestamp 1688980957
transform 1 0 25300 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold320
timestamp 1688980957
transform 1 0 25760 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold321
timestamp 1688980957
transform 1 0 29624 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold322
timestamp 1688980957
transform 1 0 27784 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold323
timestamp 1688980957
transform -1 0 3588 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold324
timestamp 1688980957
transform -1 0 3588 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold325
timestamp 1688980957
transform -1 0 11592 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold326
timestamp 1688980957
transform -1 0 6992 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold327
timestamp 1688980957
transform 1 0 1472 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold328
timestamp 1688980957
transform -1 0 4508 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold329
timestamp 1688980957
transform -1 0 13156 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold330
timestamp 1688980957
transform -1 0 17388 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold331
timestamp 1688980957
transform 1 0 30912 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold332
timestamp 1688980957
transform 1 0 32200 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold333
timestamp 1688980957
transform 1 0 6532 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold334
timestamp 1688980957
transform -1 0 11132 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold335
timestamp 1688980957
transform 1 0 4324 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold336
timestamp 1688980957
transform -1 0 4508 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold337
timestamp 1688980957
transform 1 0 19688 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold338
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold339
timestamp 1688980957
transform -1 0 4508 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold340
timestamp 1688980957
transform -1 0 8280 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold341
timestamp 1688980957
transform 1 0 3404 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold342
timestamp 1688980957
transform -1 0 4508 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold343
timestamp 1688980957
transform 1 0 23092 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold344
timestamp 1688980957
transform 1 0 21988 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold345
timestamp 1688980957
transform 1 0 27140 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold346
timestamp 1688980957
transform -1 0 28060 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold347
timestamp 1688980957
transform 1 0 17204 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold348
timestamp 1688980957
transform 1 0 18492 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold349
timestamp 1688980957
transform -1 0 4508 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold350
timestamp 1688980957
transform -1 0 4140 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold351
timestamp 1688980957
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold352
timestamp 1688980957
transform -1 0 4508 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold353
timestamp 1688980957
transform -1 0 13984 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  output2 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 2852 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output3
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output4
timestamp 1688980957
transform -1 0 6164 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output5
timestamp 1688980957
transform -1 0 6256 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output6
timestamp 1688980957
transform 1 0 8832 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output7
timestamp 1688980957
transform -1 0 10764 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output8
timestamp 1688980957
transform -1 0 11408 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output9
timestamp 1688980957
transform -1 0 14904 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output10
timestamp 1688980957
transform 1 0 15088 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output11
timestamp 1688980957
transform -1 0 16560 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output12
timestamp 1688980957
transform -1 0 20148 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output13
timestamp 1688980957
transform -1 0 5244 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output14
timestamp 1688980957
transform 1 0 22172 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output15
timestamp 1688980957
transform 1 0 24380 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output16
timestamp 1688980957
transform 1 0 29532 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output17
timestamp 1688980957
transform 1 0 27416 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output18
timestamp 1688980957
transform 1 0 30360 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output19
timestamp 1688980957
transform 1 0 33580 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output20
timestamp 1688980957
transform 1 0 35052 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output21
timestamp 1688980957
transform 1 0 33120 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output22
timestamp 1688980957
transform 1 0 31648 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output23
timestamp 1688980957
transform 1 0 34684 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output24
timestamp 1688980957
transform 1 0 20240 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output25
timestamp 1688980957
transform -1 0 26220 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output26
timestamp 1688980957
transform -1 0 27600 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output27
timestamp 1688980957
transform 1 0 28428 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output28
timestamp 1688980957
transform 1 0 29900 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output29
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output30
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output31
timestamp 1688980957
transform -1 0 35420 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output32
timestamp 1688980957
transform -1 0 36064 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output33
timestamp 1688980957
transform 1 0 35696 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output34
timestamp 1688980957
transform 1 0 35696 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output35
timestamp 1688980957
transform 1 0 23276 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output36
timestamp 1688980957
transform 1 0 36064 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output37
timestamp 1688980957
transform 1 0 35696 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output38
timestamp 1688980957
transform 1 0 36064 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output39
timestamp 1688980957
transform 1 0 35696 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output40
timestamp 1688980957
transform 1 0 36064 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output41
timestamp 1688980957
transform 1 0 35696 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output42
timestamp 1688980957
transform 1 0 36064 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output43
timestamp 1688980957
transform 1 0 35696 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output44
timestamp 1688980957
transform 1 0 35696 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output45
timestamp 1688980957
transform 1 0 35696 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output46
timestamp 1688980957
transform 1 0 34224 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output47
timestamp 1688980957
transform 1 0 36064 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output48
timestamp 1688980957
transform 1 0 35696 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output49
timestamp 1688980957
transform 1 0 36064 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output50
timestamp 1688980957
transform 1 0 35696 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output51
timestamp 1688980957
transform 1 0 36064 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output52
timestamp 1688980957
transform 1 0 35696 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output53
timestamp 1688980957
transform 1 0 36064 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output54
timestamp 1688980957
transform 1 0 32476 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output55
timestamp 1688980957
transform 1 0 33948 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output56
timestamp 1688980957
transform 1 0 35696 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output57
timestamp 1688980957
transform 1 0 36064 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output58
timestamp 1688980957
transform -1 0 8832 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output59
timestamp 1688980957
transform -1 0 9936 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output60
timestamp 1688980957
transform -1 0 10764 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output61
timestamp 1688980957
transform -1 0 11408 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output62
timestamp 1688980957
transform -1 0 13616 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output63
timestamp 1688980957
transform -1 0 15916 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output64
timestamp 1688980957
transform -1 0 15088 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output65
timestamp 1688980957
transform 1 0 17664 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output66
timestamp 1688980957
transform 1 0 19504 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output67
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output68
timestamp 1688980957
transform -1 0 7360 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output69
timestamp 1688980957
transform -1 0 2852 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output70
timestamp 1688980957
transform -1 0 2852 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output71
timestamp 1688980957
transform -1 0 2852 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output72
timestamp 1688980957
transform -1 0 2852 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output73
timestamp 1688980957
transform -1 0 4324 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output74
timestamp 1688980957
transform -1 0 2852 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output75
timestamp 1688980957
transform -1 0 4324 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output76
timestamp 1688980957
transform -1 0 2852 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output77
timestamp 1688980957
transform -1 0 2852 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output78
timestamp 1688980957
transform -1 0 2852 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output79
timestamp 1688980957
transform -1 0 2852 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output80
timestamp 1688980957
transform -1 0 2852 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output81
timestamp 1688980957
transform -1 0 2852 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output82
timestamp 1688980957
transform -1 0 2852 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output83
timestamp 1688980957
transform -1 0 2852 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output84
timestamp 1688980957
transform -1 0 2852 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output85
timestamp 1688980957
transform -1 0 2852 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output86
timestamp 1688980957
transform -1 0 2852 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output87
timestamp 1688980957
transform -1 0 2852 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output88
timestamp 1688980957
transform -1 0 2852 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output89
timestamp 1688980957
transform -1 0 2852 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 37812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 37812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 37812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 37812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 37812 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 37812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 37812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 37812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 37812 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 37812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 37812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 37812 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 37812 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 37812 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 37812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 37812 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 37812 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 37812 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 37812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 37812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 37812 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 37812 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 37812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 37812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 37812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 37812 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 37812 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 37812 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 37812 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 37812 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 37812 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 37812 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 37812 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 37812 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 37812 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 37812 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 37812 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 37812 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 37812 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 37812 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 37812 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 37812 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 37812 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 37812 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 37812 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 37812 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 37812 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 37812 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 37812 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 37812 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 37812 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 37812 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 37812 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 37812 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 37812 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 37812 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 37812 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 37812 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 37812 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 37812 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 37812 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 37812 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 37812 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1688980957
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1688980957
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1688980957
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1688980957
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1688980957
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1688980957
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1688980957
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1688980957
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1688980957
transform 1 0 6256 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1688980957
transform 1 0 11408 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1688980957
transform 1 0 16560 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1688980957
transform 1 0 21712 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1688980957
transform 1 0 26864 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1688980957
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1688980957
transform 1 0 32016 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1688980957
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1688980957
transform 1 0 37168 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  unused_tie_97 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  unused_tie_98
timestamp 1688980957
transform -1 0 3588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  unused_tie_99
timestamp 1688980957
transform 1 0 4508 0 1 2176
box -38 -48 314 592
<< labels >>
flabel metal2 s 1766 0 1822 800 0 FreeSans 224 90 0 0 irq[0]
port 0 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 irq[1]
port 1 nsew signal tristate
flabel metal2 s 4710 0 4766 800 0 FreeSans 224 90 0 0 irq[2]
port 2 nsew signal tristate
flabel metal3 s 0 34824 800 34944 0 FreeSans 480 0 0 0 la_data_out[0]
port 3 nsew signal tristate
flabel metal2 s 2870 38200 2926 39000 0 FreeSans 224 90 0 0 la_data_out[10]
port 4 nsew signal tristate
flabel metal2 s 4618 38200 4674 39000 0 FreeSans 224 90 0 0 la_data_out[11]
port 5 nsew signal tristate
flabel metal2 s 6366 38200 6422 39000 0 FreeSans 224 90 0 0 la_data_out[12]
port 6 nsew signal tristate
flabel metal2 s 8114 38200 8170 39000 0 FreeSans 224 90 0 0 la_data_out[13]
port 7 nsew signal tristate
flabel metal2 s 9862 38200 9918 39000 0 FreeSans 224 90 0 0 la_data_out[14]
port 8 nsew signal tristate
flabel metal2 s 11610 38200 11666 39000 0 FreeSans 224 90 0 0 la_data_out[15]
port 9 nsew signal tristate
flabel metal2 s 13358 38200 13414 39000 0 FreeSans 224 90 0 0 la_data_out[16]
port 10 nsew signal tristate
flabel metal2 s 15106 38200 15162 39000 0 FreeSans 224 90 0 0 la_data_out[17]
port 11 nsew signal tristate
flabel metal2 s 16854 38200 16910 39000 0 FreeSans 224 90 0 0 la_data_out[18]
port 12 nsew signal tristate
flabel metal2 s 18602 38200 18658 39000 0 FreeSans 224 90 0 0 la_data_out[19]
port 13 nsew signal tristate
flabel metal2 s 1122 38200 1178 39000 0 FreeSans 224 90 0 0 la_data_out[1]
port 14 nsew signal tristate
flabel metal2 s 22098 38200 22154 39000 0 FreeSans 224 90 0 0 la_data_out[20]
port 15 nsew signal tristate
flabel metal2 s 23846 38200 23902 39000 0 FreeSans 224 90 0 0 la_data_out[21]
port 16 nsew signal tristate
flabel metal2 s 25594 38200 25650 39000 0 FreeSans 224 90 0 0 la_data_out[22]
port 17 nsew signal tristate
flabel metal2 s 27342 38200 27398 39000 0 FreeSans 224 90 0 0 la_data_out[23]
port 18 nsew signal tristate
flabel metal2 s 29090 38200 29146 39000 0 FreeSans 224 90 0 0 la_data_out[24]
port 19 nsew signal tristate
flabel metal2 s 30838 38200 30894 39000 0 FreeSans 224 90 0 0 la_data_out[25]
port 20 nsew signal tristate
flabel metal2 s 32586 38200 32642 39000 0 FreeSans 224 90 0 0 la_data_out[26]
port 21 nsew signal tristate
flabel metal2 s 34334 38200 34390 39000 0 FreeSans 224 90 0 0 la_data_out[27]
port 22 nsew signal tristate
flabel metal2 s 36082 38200 36138 39000 0 FreeSans 224 90 0 0 la_data_out[28]
port 23 nsew signal tristate
flabel metal2 s 37830 38200 37886 39000 0 FreeSans 224 90 0 0 la_data_out[29]
port 24 nsew signal tristate
flabel metal2 s 20350 38200 20406 39000 0 FreeSans 224 90 0 0 la_data_out[2]
port 25 nsew signal tristate
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 la_data_out[30]
port 26 nsew signal tristate
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 la_data_out[31]
port 27 nsew signal tristate
flabel metal2 s 26790 0 26846 800 0 FreeSans 224 90 0 0 la_data_out[32]
port 28 nsew signal tristate
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 la_data_out[33]
port 29 nsew signal tristate
flabel metal2 s 29734 0 29790 800 0 FreeSans 224 90 0 0 la_data_out[34]
port 30 nsew signal tristate
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 la_data_out[35]
port 31 nsew signal tristate
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 la_data_out[36]
port 32 nsew signal tristate
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 la_data_out[37]
port 33 nsew signal tristate
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 la_data_out[38]
port 34 nsew signal tristate
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 la_data_out[39]
port 35 nsew signal tristate
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 la_data_out[3]
port 36 nsew signal tristate
flabel metal3 s 38200 5448 39000 5568 0 FreeSans 480 0 0 0 la_data_out[40]
port 37 nsew signal tristate
flabel metal3 s 38200 7080 39000 7200 0 FreeSans 480 0 0 0 la_data_out[41]
port 38 nsew signal tristate
flabel metal3 s 38200 8712 39000 8832 0 FreeSans 480 0 0 0 la_data_out[42]
port 39 nsew signal tristate
flabel metal3 s 38200 10344 39000 10464 0 FreeSans 480 0 0 0 la_data_out[43]
port 40 nsew signal tristate
flabel metal3 s 38200 11976 39000 12096 0 FreeSans 480 0 0 0 la_data_out[44]
port 41 nsew signal tristate
flabel metal3 s 38200 13608 39000 13728 0 FreeSans 480 0 0 0 la_data_out[45]
port 42 nsew signal tristate
flabel metal3 s 38200 15240 39000 15360 0 FreeSans 480 0 0 0 la_data_out[46]
port 43 nsew signal tristate
flabel metal3 s 38200 16872 39000 16992 0 FreeSans 480 0 0 0 la_data_out[47]
port 44 nsew signal tristate
flabel metal3 s 38200 18504 39000 18624 0 FreeSans 480 0 0 0 la_data_out[48]
port 45 nsew signal tristate
flabel metal3 s 38200 20136 39000 20256 0 FreeSans 480 0 0 0 la_data_out[49]
port 46 nsew signal tristate
flabel metal3 s 38200 3816 39000 3936 0 FreeSans 480 0 0 0 la_data_out[4]
port 47 nsew signal tristate
flabel metal3 s 38200 23400 39000 23520 0 FreeSans 480 0 0 0 la_data_out[50]
port 48 nsew signal tristate
flabel metal3 s 38200 25032 39000 25152 0 FreeSans 480 0 0 0 la_data_out[51]
port 49 nsew signal tristate
flabel metal3 s 38200 26664 39000 26784 0 FreeSans 480 0 0 0 la_data_out[52]
port 50 nsew signal tristate
flabel metal3 s 38200 28296 39000 28416 0 FreeSans 480 0 0 0 la_data_out[53]
port 51 nsew signal tristate
flabel metal3 s 38200 29928 39000 30048 0 FreeSans 480 0 0 0 la_data_out[54]
port 52 nsew signal tristate
flabel metal3 s 38200 31560 39000 31680 0 FreeSans 480 0 0 0 la_data_out[55]
port 53 nsew signal tristate
flabel metal3 s 38200 33192 39000 33312 0 FreeSans 480 0 0 0 la_data_out[56]
port 54 nsew signal tristate
flabel metal3 s 38200 34824 39000 34944 0 FreeSans 480 0 0 0 la_data_out[57]
port 55 nsew signal tristate
flabel metal3 s 38200 36456 39000 36576 0 FreeSans 480 0 0 0 la_data_out[58]
port 56 nsew signal tristate
flabel metal3 s 38200 38088 39000 38208 0 FreeSans 480 0 0 0 la_data_out[59]
port 57 nsew signal tristate
flabel metal3 s 38200 21768 39000 21888 0 FreeSans 480 0 0 0 la_data_out[5]
port 58 nsew signal tristate
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 la_data_out[60]
port 59 nsew signal tristate
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 la_data_out[61]
port 60 nsew signal tristate
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 la_data_out[62]
port 61 nsew signal tristate
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 la_data_out[63]
port 62 nsew signal tristate
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 la_data_out[64]
port 63 nsew signal tristate
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 la_data_out[65]
port 64 nsew signal tristate
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 la_data_out[66]
port 65 nsew signal tristate
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 la_data_out[67]
port 66 nsew signal tristate
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 la_data_out[68]
port 67 nsew signal tristate
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 la_data_out[69]
port 68 nsew signal tristate
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 la_data_out[6]
port 69 nsew signal tristate
flabel metal3 s 0 18504 800 18624 0 FreeSans 480 0 0 0 la_data_out[70]
port 70 nsew signal tristate
flabel metal3 s 0 20136 800 20256 0 FreeSans 480 0 0 0 la_data_out[71]
port 71 nsew signal tristate
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 la_data_out[72]
port 72 nsew signal tristate
flabel metal3 s 0 23400 800 23520 0 FreeSans 480 0 0 0 la_data_out[73]
port 73 nsew signal tristate
flabel metal3 s 0 25032 800 25152 0 FreeSans 480 0 0 0 la_data_out[74]
port 74 nsew signal tristate
flabel metal3 s 0 26664 800 26784 0 FreeSans 480 0 0 0 la_data_out[75]
port 75 nsew signal tristate
flabel metal3 s 0 28296 800 28416 0 FreeSans 480 0 0 0 la_data_out[76]
port 76 nsew signal tristate
flabel metal3 s 0 29928 800 30048 0 FreeSans 480 0 0 0 la_data_out[77]
port 77 nsew signal tristate
flabel metal3 s 0 31560 800 31680 0 FreeSans 480 0 0 0 la_data_out[78]
port 78 nsew signal tristate
flabel metal3 s 0 33192 800 33312 0 FreeSans 480 0 0 0 la_data_out[79]
port 79 nsew signal tristate
flabel metal3 s 0 16872 800 16992 0 FreeSans 480 0 0 0 la_data_out[7]
port 80 nsew signal tristate
flabel metal3 s 0 3816 800 3936 0 FreeSans 480 0 0 0 la_data_out[80]
port 81 nsew signal tristate
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 la_data_out[81]
port 82 nsew signal tristate
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 la_data_out[82]
port 83 nsew signal tristate
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 la_data_out[83]
port 84 nsew signal tristate
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 la_data_out[84]
port 85 nsew signal tristate
flabel metal3 s 0 11976 800 12096 0 FreeSans 480 0 0 0 la_data_out[85]
port 86 nsew signal tristate
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 la_data_out[86]
port 87 nsew signal tristate
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 la_data_out[87]
port 88 nsew signal tristate
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 la_data_out[8]
port 89 nsew signal tristate
flabel metal3 s 0 36456 800 36576 0 FreeSans 480 0 0 0 la_data_out[9]
port 90 nsew signal tristate
flabel metal4 s 4208 2128 4528 36496 0 FreeSans 1920 90 0 0 vccd1
port 91 nsew power bidirectional
flabel metal4 s 34928 2128 35248 36496 0 FreeSans 1920 90 0 0 vccd1
port 91 nsew power bidirectional
flabel metal4 s 19568 2128 19888 36496 0 FreeSans 1920 90 0 0 vssd1
port 92 nsew ground bidirectional
flabel metal3 s 38200 552 39000 672 0 FreeSans 480 0 0 0 wb_clk_i
port 93 nsew signal input
flabel metal3 s 38200 2184 39000 2304 0 FreeSans 480 0 0 0 wb_rst_i
port 94 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 39000 39000
<< end >>
