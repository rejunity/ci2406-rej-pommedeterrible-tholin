// This is the unpowered netlist.
module scrapcpu (rst_n,
    wb_clk_i,
    io_in,
    io_oeb,
    io_out);
 input rst_n;
 input wb_clk_i;
 input [35:0] io_in;
 output [35:0] io_oeb;
 output [35:0] io_out;

 wire net158;
 wire net159;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net178;
 wire net160;
 wire net171;
 wire net161;
 wire net162;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire \A[0] ;
 wire \A[1] ;
 wire \A[2] ;
 wire \A[3] ;
 wire \A[4] ;
 wire \A[5] ;
 wire \B[0] ;
 wire \B[1] ;
 wire \B[2] ;
 wire \B[3] ;
 wire \B[4] ;
 wire \B[5] ;
 wire \MAR[0] ;
 wire \MAR[1] ;
 wire \MAR[2] ;
 wire \MAR[3] ;
 wire \MAR[4] ;
 wire \PC[0] ;
 wire \PC[1] ;
 wire \PC[2] ;
 wire \PC[3] ;
 wire \PC[4] ;
 wire \PC[5] ;
 wire \PC[6] ;
 wire \P[0] ;
 wire \P[1] ;
 wire \P[2] ;
 wire \P[3] ;
 wire \P[4] ;
 wire \P[5] ;
 wire \RAM[0][0] ;
 wire \RAM[0][1] ;
 wire \RAM[0][2] ;
 wire \RAM[0][3] ;
 wire \RAM[0][4] ;
 wire \RAM[0][5] ;
 wire \RAM[10][0] ;
 wire \RAM[10][1] ;
 wire \RAM[10][2] ;
 wire \RAM[10][3] ;
 wire \RAM[10][4] ;
 wire \RAM[10][5] ;
 wire \RAM[11][0] ;
 wire \RAM[11][1] ;
 wire \RAM[11][2] ;
 wire \RAM[11][3] ;
 wire \RAM[11][4] ;
 wire \RAM[11][5] ;
 wire \RAM[12][0] ;
 wire \RAM[12][1] ;
 wire \RAM[12][2] ;
 wire \RAM[12][3] ;
 wire \RAM[12][4] ;
 wire \RAM[12][5] ;
 wire \RAM[13][0] ;
 wire \RAM[13][1] ;
 wire \RAM[13][2] ;
 wire \RAM[13][3] ;
 wire \RAM[13][4] ;
 wire \RAM[13][5] ;
 wire \RAM[14][0] ;
 wire \RAM[14][1] ;
 wire \RAM[14][2] ;
 wire \RAM[14][3] ;
 wire \RAM[14][4] ;
 wire \RAM[14][5] ;
 wire \RAM[15][0] ;
 wire \RAM[15][1] ;
 wire \RAM[15][2] ;
 wire \RAM[15][3] ;
 wire \RAM[15][4] ;
 wire \RAM[15][5] ;
 wire \RAM[16][0] ;
 wire \RAM[16][1] ;
 wire \RAM[16][2] ;
 wire \RAM[16][3] ;
 wire \RAM[16][4] ;
 wire \RAM[16][5] ;
 wire \RAM[17][0] ;
 wire \RAM[17][1] ;
 wire \RAM[17][2] ;
 wire \RAM[17][3] ;
 wire \RAM[17][4] ;
 wire \RAM[17][5] ;
 wire \RAM[18][0] ;
 wire \RAM[18][1] ;
 wire \RAM[18][2] ;
 wire \RAM[18][3] ;
 wire \RAM[18][4] ;
 wire \RAM[18][5] ;
 wire \RAM[19][0] ;
 wire \RAM[19][1] ;
 wire \RAM[19][2] ;
 wire \RAM[19][3] ;
 wire \RAM[19][4] ;
 wire \RAM[19][5] ;
 wire \RAM[1][0] ;
 wire \RAM[1][1] ;
 wire \RAM[1][2] ;
 wire \RAM[1][3] ;
 wire \RAM[1][4] ;
 wire \RAM[1][5] ;
 wire \RAM[20][0] ;
 wire \RAM[20][1] ;
 wire \RAM[20][2] ;
 wire \RAM[20][3] ;
 wire \RAM[20][4] ;
 wire \RAM[20][5] ;
 wire \RAM[21][0] ;
 wire \RAM[21][1] ;
 wire \RAM[21][2] ;
 wire \RAM[21][3] ;
 wire \RAM[21][4] ;
 wire \RAM[21][5] ;
 wire \RAM[22][0] ;
 wire \RAM[22][1] ;
 wire \RAM[22][2] ;
 wire \RAM[22][3] ;
 wire \RAM[22][4] ;
 wire \RAM[22][5] ;
 wire \RAM[23][0] ;
 wire \RAM[23][1] ;
 wire \RAM[23][2] ;
 wire \RAM[23][3] ;
 wire \RAM[23][4] ;
 wire \RAM[23][5] ;
 wire \RAM[24][0] ;
 wire \RAM[24][1] ;
 wire \RAM[24][2] ;
 wire \RAM[24][3] ;
 wire \RAM[24][4] ;
 wire \RAM[24][5] ;
 wire \RAM[25][0] ;
 wire \RAM[25][1] ;
 wire \RAM[25][2] ;
 wire \RAM[25][3] ;
 wire \RAM[25][4] ;
 wire \RAM[25][5] ;
 wire \RAM[26][0] ;
 wire \RAM[26][1] ;
 wire \RAM[26][2] ;
 wire \RAM[26][3] ;
 wire \RAM[26][4] ;
 wire \RAM[26][5] ;
 wire \RAM[27][0] ;
 wire \RAM[27][1] ;
 wire \RAM[27][2] ;
 wire \RAM[27][3] ;
 wire \RAM[27][4] ;
 wire \RAM[27][5] ;
 wire \RAM[28][0] ;
 wire \RAM[28][1] ;
 wire \RAM[28][2] ;
 wire \RAM[28][3] ;
 wire \RAM[28][4] ;
 wire \RAM[28][5] ;
 wire \RAM[29][0] ;
 wire \RAM[29][1] ;
 wire \RAM[29][2] ;
 wire \RAM[29][3] ;
 wire \RAM[29][4] ;
 wire \RAM[29][5] ;
 wire \RAM[2][0] ;
 wire \RAM[2][1] ;
 wire \RAM[2][2] ;
 wire \RAM[2][3] ;
 wire \RAM[2][4] ;
 wire \RAM[2][5] ;
 wire \RAM[30][0] ;
 wire \RAM[30][1] ;
 wire \RAM[30][2] ;
 wire \RAM[30][3] ;
 wire \RAM[30][4] ;
 wire \RAM[30][5] ;
 wire \RAM[31][0] ;
 wire \RAM[31][1] ;
 wire \RAM[31][2] ;
 wire \RAM[31][3] ;
 wire \RAM[31][4] ;
 wire \RAM[31][5] ;
 wire \RAM[32][0] ;
 wire \RAM[32][1] ;
 wire \RAM[32][2] ;
 wire \RAM[32][3] ;
 wire \RAM[32][4] ;
 wire \RAM[32][5] ;
 wire \RAM[33][0] ;
 wire \RAM[33][1] ;
 wire \RAM[33][2] ;
 wire \RAM[33][3] ;
 wire \RAM[33][4] ;
 wire \RAM[33][5] ;
 wire \RAM[34][0] ;
 wire \RAM[34][1] ;
 wire \RAM[34][2] ;
 wire \RAM[34][3] ;
 wire \RAM[34][4] ;
 wire \RAM[34][5] ;
 wire \RAM[35][0] ;
 wire \RAM[35][1] ;
 wire \RAM[35][2] ;
 wire \RAM[35][3] ;
 wire \RAM[35][4] ;
 wire \RAM[35][5] ;
 wire \RAM[36][0] ;
 wire \RAM[36][1] ;
 wire \RAM[36][2] ;
 wire \RAM[36][3] ;
 wire \RAM[36][4] ;
 wire \RAM[36][5] ;
 wire \RAM[37][0] ;
 wire \RAM[37][1] ;
 wire \RAM[37][2] ;
 wire \RAM[37][3] ;
 wire \RAM[37][4] ;
 wire \RAM[37][5] ;
 wire \RAM[38][0] ;
 wire \RAM[38][1] ;
 wire \RAM[38][2] ;
 wire \RAM[38][3] ;
 wire \RAM[38][4] ;
 wire \RAM[38][5] ;
 wire \RAM[39][0] ;
 wire \RAM[39][1] ;
 wire \RAM[39][2] ;
 wire \RAM[39][3] ;
 wire \RAM[39][4] ;
 wire \RAM[39][5] ;
 wire \RAM[3][0] ;
 wire \RAM[3][1] ;
 wire \RAM[3][2] ;
 wire \RAM[3][3] ;
 wire \RAM[3][4] ;
 wire \RAM[3][5] ;
 wire \RAM[40][0] ;
 wire \RAM[40][1] ;
 wire \RAM[40][2] ;
 wire \RAM[40][3] ;
 wire \RAM[40][4] ;
 wire \RAM[40][5] ;
 wire \RAM[41][0] ;
 wire \RAM[41][1] ;
 wire \RAM[41][2] ;
 wire \RAM[41][3] ;
 wire \RAM[41][4] ;
 wire \RAM[41][5] ;
 wire \RAM[42][0] ;
 wire \RAM[42][1] ;
 wire \RAM[42][2] ;
 wire \RAM[42][3] ;
 wire \RAM[42][4] ;
 wire \RAM[42][5] ;
 wire \RAM[43][0] ;
 wire \RAM[43][1] ;
 wire \RAM[43][2] ;
 wire \RAM[43][3] ;
 wire \RAM[43][4] ;
 wire \RAM[43][5] ;
 wire \RAM[44][0] ;
 wire \RAM[44][1] ;
 wire \RAM[44][2] ;
 wire \RAM[44][3] ;
 wire \RAM[44][4] ;
 wire \RAM[44][5] ;
 wire \RAM[45][0] ;
 wire \RAM[45][1] ;
 wire \RAM[45][2] ;
 wire \RAM[45][3] ;
 wire \RAM[45][4] ;
 wire \RAM[45][5] ;
 wire \RAM[46][0] ;
 wire \RAM[46][1] ;
 wire \RAM[46][2] ;
 wire \RAM[46][3] ;
 wire \RAM[46][4] ;
 wire \RAM[46][5] ;
 wire \RAM[47][0] ;
 wire \RAM[47][1] ;
 wire \RAM[47][2] ;
 wire \RAM[47][3] ;
 wire \RAM[47][4] ;
 wire \RAM[47][5] ;
 wire \RAM[48][0] ;
 wire \RAM[48][1] ;
 wire \RAM[48][2] ;
 wire \RAM[48][3] ;
 wire \RAM[48][4] ;
 wire \RAM[48][5] ;
 wire \RAM[49][0] ;
 wire \RAM[49][1] ;
 wire \RAM[49][2] ;
 wire \RAM[49][3] ;
 wire \RAM[49][4] ;
 wire \RAM[49][5] ;
 wire \RAM[4][0] ;
 wire \RAM[4][1] ;
 wire \RAM[4][2] ;
 wire \RAM[4][3] ;
 wire \RAM[4][4] ;
 wire \RAM[4][5] ;
 wire \RAM[50][0] ;
 wire \RAM[50][1] ;
 wire \RAM[50][2] ;
 wire \RAM[50][3] ;
 wire \RAM[50][4] ;
 wire \RAM[50][5] ;
 wire \RAM[51][0] ;
 wire \RAM[51][1] ;
 wire \RAM[51][2] ;
 wire \RAM[51][3] ;
 wire \RAM[51][4] ;
 wire \RAM[51][5] ;
 wire \RAM[52][0] ;
 wire \RAM[52][1] ;
 wire \RAM[52][2] ;
 wire \RAM[52][3] ;
 wire \RAM[52][4] ;
 wire \RAM[52][5] ;
 wire \RAM[53][0] ;
 wire \RAM[53][1] ;
 wire \RAM[53][2] ;
 wire \RAM[53][3] ;
 wire \RAM[53][4] ;
 wire \RAM[53][5] ;
 wire \RAM[54][0] ;
 wire \RAM[54][1] ;
 wire \RAM[54][2] ;
 wire \RAM[54][3] ;
 wire \RAM[54][4] ;
 wire \RAM[54][5] ;
 wire \RAM[55][0] ;
 wire \RAM[55][1] ;
 wire \RAM[55][2] ;
 wire \RAM[55][3] ;
 wire \RAM[55][4] ;
 wire \RAM[55][5] ;
 wire \RAM[56][0] ;
 wire \RAM[56][1] ;
 wire \RAM[56][2] ;
 wire \RAM[56][3] ;
 wire \RAM[56][4] ;
 wire \RAM[56][5] ;
 wire \RAM[57][0] ;
 wire \RAM[57][1] ;
 wire \RAM[57][2] ;
 wire \RAM[57][3] ;
 wire \RAM[57][4] ;
 wire \RAM[57][5] ;
 wire \RAM[59][0] ;
 wire \RAM[59][1] ;
 wire \RAM[59][2] ;
 wire \RAM[59][3] ;
 wire \RAM[59][4] ;
 wire \RAM[59][5] ;
 wire \RAM[5][0] ;
 wire \RAM[5][1] ;
 wire \RAM[5][2] ;
 wire \RAM[5][3] ;
 wire \RAM[5][4] ;
 wire \RAM[5][5] ;
 wire \RAM[61][0] ;
 wire \RAM[61][1] ;
 wire \RAM[61][2] ;
 wire \RAM[61][3] ;
 wire \RAM[61][4] ;
 wire \RAM[61][5] ;
 wire \RAM[62][0] ;
 wire \RAM[62][1] ;
 wire \RAM[62][2] ;
 wire \RAM[62][3] ;
 wire \RAM[62][4] ;
 wire \RAM[62][5] ;
 wire \RAM[6][0] ;
 wire \RAM[6][1] ;
 wire \RAM[6][2] ;
 wire \RAM[6][3] ;
 wire \RAM[6][4] ;
 wire \RAM[6][5] ;
 wire \RAM[7][0] ;
 wire \RAM[7][1] ;
 wire \RAM[7][2] ;
 wire \RAM[7][3] ;
 wire \RAM[7][4] ;
 wire \RAM[7][5] ;
 wire \RAM[8][0] ;
 wire \RAM[8][1] ;
 wire \RAM[8][2] ;
 wire \RAM[8][3] ;
 wire \RAM[8][4] ;
 wire \RAM[8][5] ;
 wire \RAM[9][0] ;
 wire \RAM[9][1] ;
 wire \RAM[9][2] ;
 wire \RAM[9][3] ;
 wire \RAM[9][4] ;
 wire \RAM[9][5] ;
 wire ROM_OEB;
 wire \ROM_addr_buff[0] ;
 wire \ROM_addr_buff[10] ;
 wire \ROM_addr_buff[11] ;
 wire \ROM_addr_buff[1] ;
 wire \ROM_addr_buff[2] ;
 wire \ROM_addr_buff[3] ;
 wire \ROM_addr_buff[4] ;
 wire \ROM_addr_buff[5] ;
 wire \ROM_addr_buff[6] ;
 wire \ROM_addr_buff[7] ;
 wire \ROM_addr_buff[8] ;
 wire \ROM_addr_buff[9] ;
 wire \ROM_dest[0] ;
 wire \ROM_dest[1] ;
 wire \ROM_dest[2] ;
 wire \ROM_spi_cycle[0] ;
 wire \ROM_spi_cycle[1] ;
 wire \ROM_spi_cycle[2] ;
 wire \ROM_spi_cycle[3] ;
 wire \ROM_spi_cycle[4] ;
 wire \ROM_spi_dat_out[0] ;
 wire \ROM_spi_dat_out[1] ;
 wire \ROM_spi_dat_out[2] ;
 wire \ROM_spi_dat_out[3] ;
 wire \ROM_spi_dat_out[4] ;
 wire \ROM_spi_dat_out[5] ;
 wire \ROM_spi_dat_out[6] ;
 wire \ROM_spi_dat_out[7] ;
 wire ROM_spi_mode;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0__leaf_wb_clk_i;
 wire clknet_3_1__leaf_wb_clk_i;
 wire clknet_3_2__leaf_wb_clk_i;
 wire clknet_3_3__leaf_wb_clk_i;
 wire clknet_3_4__leaf_wb_clk_i;
 wire clknet_3_5__leaf_wb_clk_i;
 wire clknet_3_6__leaf_wb_clk_i;
 wire clknet_3_7__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire \imm_buff[0] ;
 wire \imm_buff[1] ;
 wire \imm_buff[2] ;
 wire \imm_buff[3] ;
 wire \imm_buff[4] ;
 wire \imm_buff[5] ;
 wire \insin[0] ;
 wire \insin[1] ;
 wire \insin[2] ;
 wire \insin[3] ;
 wire \insin[4] ;
 wire \insin[5] ;
 wire \instr_cycle[1] ;
 wire \instr_cycle[2] ;
 wire \last_A[0] ;
 wire \last_A[1] ;
 wire \last_A[2] ;
 wire \last_A[3] ;
 wire \last_A[4] ;
 wire \last_A[5] ;
 wire \last_B[0] ;
 wire \last_B[1] ;
 wire \last_B[2] ;
 wire \last_B[3] ;
 wire \last_B[4] ;
 wire \last_B[5] ;
 wire \last_MAR[0] ;
 wire \last_MAR[1] ;
 wire \last_MAR[2] ;
 wire \last_MAR[3] ;
 wire \last_MAR[4] ;
 wire \last_MAR[5] ;
 wire \last_PC[0] ;
 wire \last_PC[10] ;
 wire \last_PC[11] ;
 wire \last_PC[1] ;
 wire \last_PC[2] ;
 wire \last_PC[3] ;
 wire \last_PC[4] ;
 wire \last_PC[5] ;
 wire \last_PC[6] ;
 wire \last_PC[7] ;
 wire \last_PC[8] ;
 wire \last_PC[9] ;
 wire \last_P[0] ;
 wire \last_P[1] ;
 wire \last_P[2] ;
 wire \last_P[3] ;
 wire \last_P[4] ;
 wire \last_P[5] ;
 wire \last_addr[0] ;
 wire \last_addr[10] ;
 wire \last_addr[11] ;
 wire \last_addr[1] ;
 wire \last_addr[2] ;
 wire \last_addr[3] ;
 wire \last_addr[4] ;
 wire \last_addr[5] ;
 wire \last_addr[6] ;
 wire \last_addr[7] ;
 wire \last_addr[8] ;
 wire \last_addr[9] ;
 wire \last_flags[0] ;
 wire \last_flags[1] ;
 wire last_inter;
 wire \mem_cycle[0] ;
 wire \mem_cycle[1] ;
 wire \mem_cycle[2] ;
 wire \mem_cycle[3] ;
 wire \mem_cycle[4] ;
 wire needs_irupt;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net109;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net110;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net111;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net112;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net113;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net114;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net115;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net116;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net117;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net118;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net119;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net12;
 wire net120;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net121;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net122;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net123;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net124;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net125;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net126;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net16;
 wire net17;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire spi_clkdiv;
 wire \startup_cycle[0] ;
 wire \startup_cycle[1] ;
 wire \startup_cycle[2] ;
 wire \startup_cycle[3] ;
 wire \startup_cycle[4] ;
 wire \startup_cycle[5] ;
 wire \startup_cycle[6] ;

 sky130_fd_sc_hd__diode_2 ANTENNA__1604__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__1616__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__1620__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__1622__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__1623__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__1624__A (.DIODE(\MAR[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1625__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__1640__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1640__B (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1641__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1641__B (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1642__A (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1642__B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__1642__C (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__1669__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__1670__A (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1670__B (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1671__B (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__1678__B (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1681__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__1682__A1 (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1684__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__1685__A (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1686__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__1687__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__1687__A2 (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1687__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__1687__C1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__1693__A2 (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1693__C1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__1694__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__1697__B1 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1698__B (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__1698__C (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1699__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__1700__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__1702__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__1703__B2 (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1703__C1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__1708__B (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1710__C (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1712__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__1714__B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__1715__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__1715__B (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__1716__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__1716__B (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__1717__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__1717__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__1718__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__1718__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__1719__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__1719__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__1720__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__1720__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__1721__S0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__1721__S1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__1722__S0 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__1722__S1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__1723__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__1724__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1725__S (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__1726__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__1727__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1727__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__1728__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1729__S0 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__1729__S1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__1730__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1732__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__1733__S (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__1734__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1735__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1735__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1736__S0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__1736__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__1737__S0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__1737__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__1738__S0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__1738__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__1740__S0 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__1740__S1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__1741__S1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__1742__S (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__1743__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1744__B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__1745__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__1745__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1746__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__1746__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__1747__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__1748__S0 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1748__S1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__1749__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__1750__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__1751__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__1752__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__1753__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1754__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__1754__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__1755__A (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1756__A1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1756__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__1757__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__1757__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__1759__C1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1760__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__1760__B (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__1763__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1764__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__1765__A2 (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1768__A2 (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1768__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__1769__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__1769__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__1770__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__1771__A0 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__1772__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__1773__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__1773__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__1774__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__1774__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__1775__S0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__1775__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__1776__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__1776__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__1777__S0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__1777__S1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__1778__S0 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__1778__S1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__1779__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__1780__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__1781__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__1781__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__1782__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1783__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1783__C1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__1784__S0 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__1784__S1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__1787__S (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__1788__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1788__B1 (.DIODE(\MAR[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1789__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__1790__S0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__1790__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__1791__S0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__1791__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__1792__S0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__1792__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__1794__S0 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__1794__S1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__1795__S1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__1797__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1799__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__1799__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1800__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__1800__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__1801__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__1802__S0 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1802__S1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__1803__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__1804__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__1805__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__1806__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__1807__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1808__A1 (.DIODE(\MAR[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1808__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1809__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__1809__C1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1810__A1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1811__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__1813__C1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1814__A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__1814__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1815__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__1816__A2 (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1817__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__1817__B1 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1818__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__1820__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__1820__C1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__1823__B (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1824__C (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1825__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__1825__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__1826__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__1826__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__1827__S0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__1827__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__1828__S0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__1828__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__1829__S0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__1829__S1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__1830__S0 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__1830__S1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__1831__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__1832__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1833__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__1834__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__1835__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1835__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__1836__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1837__S0 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__1837__S1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__1838__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1839__S (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__1840__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__1841__S (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__1842__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1843__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1844__S0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__1844__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__1845__S0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__1845__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__1848__S0 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__1848__S1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__1849__S0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__1849__S1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__1850__S (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__1851__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1853__A1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__1853__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1854__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__1854__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__1855__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__1856__S0 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1856__S1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__1857__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__1858__S (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1859__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__1860__S (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1861__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1862__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__1862__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__1863__A1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1864__A1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1865__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__1867__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1868__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1869__A1 (.DIODE(_0561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1869__C1 (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1870__B (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1872__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__1872__B1 (.DIODE(_0796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1873__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__1874__A0 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__1875__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__1876__S0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__1876__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__1877__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__1877__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__1878__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__1878__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__1879__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__1879__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__1880__S0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__1880__S1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__1881__S0 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__1881__S1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__1882__S (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__1883__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1884__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__1885__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__1886__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1886__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__1887__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1888__S1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__1889__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1890__S (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__1891__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__1893__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1894__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1894__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1895__S0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__1895__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__1896__S0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__1896__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__1897__S0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__1897__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__1899__S0 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__1899__S1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__1900__S0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__1900__S1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__1902__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1904__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__1904__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1905__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__1905__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__1906__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__1907__S0 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1907__S1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__1908__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__1909__S (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1910__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__1911__S (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1912__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1913__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__1913__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__1914__A1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1915__A1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1916__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__1918__B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1919__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1920__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__1921__C1 (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1922__B (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1925__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__1925__B1 (.DIODE(_0848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1926__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__1928__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__1928__C1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__1929__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__1929__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__1930__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__1930__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__1931__S0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__1931__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__1932__S0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__1932__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__1933__S0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__1933__S1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__1934__S0 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__1934__S1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__1935__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__1936__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1937__S (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__1938__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__1939__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1939__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1940__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1941__S1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__1942__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__1943__S (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__1944__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__1945__S (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__1946__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1947__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1949__S0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__1949__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__1952__S0 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__1952__S1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__1953__S1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__1954__S (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__1955__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1957__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__1957__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1958__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__1958__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__1959__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__1960__S0 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1960__S1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__1961__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__1962__S (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1963__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__1964__S (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1965__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1966__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__1966__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__1967__A1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1968__A1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1969__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__1971__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1972__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1973__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__1974__A2 (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1975__A (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1976__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__1976__B1 (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1977__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__1978__A0 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__1979__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__1980__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__1980__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__1981__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__1981__S1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__1982__S0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__1982__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__1983__S0 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__1983__S1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__1984__S0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__1984__S1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__1985__S0 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__1985__S1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__1986__S (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__1987__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1988__S (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__1989__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__1990__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1990__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1991__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1992__S1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__1995__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__1997__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1998__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1999__S0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2000__S0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2000__S1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__2003__S0 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2003__S1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2004__S0 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2004__S1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__2006__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__2007__B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2008__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__2008__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__2009__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2009__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__2010__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2011__S0 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2011__S1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__2012__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2013__S (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2014__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__2015__S (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2016__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__2017__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2017__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__2018__A1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2019__A1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2020__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2022__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__2023__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__2024__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__2025__A2 (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2026__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__2026__B1 (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2027__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__2028__A0 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__2029__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__2030__B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2035__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__2035__B1 (.DIODE(_0796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2036__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__2037__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__2037__B2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2038__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__2039__C1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2040__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__2040__B1 (.DIODE(_0848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2041__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__2041__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__2042__B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2042__C (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2043__C1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__2044__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__2044__B1 (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2045__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__2046__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__2047__C1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2048__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__2048__B1 (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2049__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2050__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__2051__C1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2052__B (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2054__B (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2055__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2057__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__2057__A2 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2057__C1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__2059__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2059__A2 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2059__C1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__2061__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__2061__A2 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2061__C1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__2063__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__2063__A2 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2063__C1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__2064__B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2065__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__2065__B2 (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2066__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2067__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__2068__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2069__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__2069__B1 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2070__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2070__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__2071__B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2071__C (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2072__C1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2074__A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__2075__C1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2076__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2077__C1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2082__B (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2084__A (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2084__B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__2085__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__2085__B (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2085__C (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__2085__D (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__2086__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__2086__C (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__2087__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__2087__C (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__2088__A (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2089__A1 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA__2089__A2 (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2090__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__2091__A1 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA__2091__A2 (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2092__A1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2093__A2 (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2094__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2095__A2 (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2096__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__2097__A2 (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2098__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2099__A2 (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2100__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2101__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2101__B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__2102__A (.DIODE(\MAR[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2102__B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2103__A1 (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2103__A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__2103__B1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2103__C1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2103__D1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2105__A (.DIODE(_1005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2106__A0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__2108__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__2109__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__2110__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2111__A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2112__A1 (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2112__A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__2112__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2112__C1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2112__D1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__2113__B (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2114__A0 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__2115__A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2116__A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2117__A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__2118__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2119__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2160__B1 (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2167__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2168__C1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__2171__C1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__2175__A1 (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2175__C1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__2180__A2 (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2180__C1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__2184__A2 (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2184__C1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__2185__B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2185__C (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__2185__D (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__2186__B (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2187__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__2188__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2189__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__2190__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__2191__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2192__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2193__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2193__B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__2194__A_N (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2195__A (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2195__B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2195__C (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2195__D (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__2196__A (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2197__A0 (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2198__A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2200__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2201__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2202__A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2203__B (.DIODE(_1005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2204__A0 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__2205__A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2206__A0 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__2207__A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__2208__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2209__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2210__B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2212__A (.DIODE(_1005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2213__A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2214__A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2215__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__2216__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2217__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2218__A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2219__A_N (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2219__B_N (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__2219__C (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__2219__D (.DIODE(\MAR[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2220__B (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2221__A0 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__2222__A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2223__A0 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__2224__A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__2225__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2226__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2227__C (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2227__D (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__2228__C (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2228__D (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__2229__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2229__A2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2229__A3 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__2229__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__2230__B (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2231__A0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__2233__A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__2234__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__2235__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2236__A0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2237__B (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2238__A0 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__2239__A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2240__A0 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__2241__A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__2242__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2243__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2244__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__2244__B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2245__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2245__B (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2245__C (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2245__D_N (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2246__B (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2247__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__2248__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2249__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2250__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__2251__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2252__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2253__A (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2254__A1 (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2254__S (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2255__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2255__S (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2256__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__2256__S (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2257__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2257__S (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2258__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2258__S (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2259__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2259__S (.DIODE(_1091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2260__B (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2261__A0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__2263__A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__2264__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__2265__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2266__A0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2267__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2267__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2267__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__2269__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__2269__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2269__A3 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__2269__C1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2271__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__2271__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2271__A3 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2271__C1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2273__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__2273__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2273__A3 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2273__C1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2275__A1 (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2275__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2275__A3 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__2275__C1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2277__A1 (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2277__A2 (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2277__A3 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2277__C1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2279__A1 (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2279__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__2279__A3 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2279__C1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2280__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2280__A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__2280__A3 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__2280__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__2283__A0 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__2284__A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2285__A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2286__A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__2287__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2288__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2289__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2289__D (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__2290__B (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2291__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__2292__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2293__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2294__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__2295__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2296__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2297__A1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2320__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__2325__C1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__2330__C1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__2331__B (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2332__A0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__2334__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__2335__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__2336__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2337__A0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2338__A (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2339__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__2339__A2 (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2339__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__2341__A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2342__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__2343__A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2344__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__2345__A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__2346__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__2347__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2348__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__2349__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2350__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__2351__A (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2352__A (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2353__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__2354__C1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2355__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2356__C1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2357__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__2358__C1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__2359__A (.DIODE(_1001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2360__C1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__2361__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2362__C1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__2363__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2364__C1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__2365__B (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2366__A0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__2368__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__2369__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__2370__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2371__A0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2372__B (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2373__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__2374__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2375__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2376__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__2377__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2378__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2379__A (.DIODE(_1005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2380__A0 (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2381__A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2382__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__2383__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2384__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2385__A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2386__A (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2387__A0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__2389__A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__2390__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__2391__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2392__A0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2393__B (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2394__A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2395__A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2397__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2398__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2399__A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2400__B (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2401__A0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__2403__A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__2404__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__2405__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2406__A0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2407__B (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2408__A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2409__A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2411__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2412__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2413__A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2414__B (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2415__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__2417__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__2418__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__2419__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2420__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2421__B (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2422__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2423__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2424__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__2425__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2426__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2427__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2428__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2428__B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__2428__C (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__2428__D (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__2430__A (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2431__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__2432__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__2433__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__2434__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__2435__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2436__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2437__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__2437__A2 (.DIODE(_0989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2437__A3 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__2437__B1 (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2438__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__2439__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2440__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2441__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__2442__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2443__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2444__A (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2445__A0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__2447__A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__2448__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__2449__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2450__A0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2451__A (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2452__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__2453__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__2454__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2455__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__2456__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2457__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2458__A (.DIODE(_1005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2459__A0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__2461__A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__2462__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__2463__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2464__A0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2465__A (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2466__A0 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__2467__A0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__2468__A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2469__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__2470__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2471__A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2472__A (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2473__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__2475__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__2476__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__2477__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2478__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2479__A (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2479__B (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2480__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2480__B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__2480__C (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__2480__D_N (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__2481__A (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2482__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__2483__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2484__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__2485__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__2486__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2487__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2488__A (.DIODE(_1005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2489__A0 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__2490__A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2491__A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2492__A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__2493__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2494__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2495__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2496__B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2498__A0 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__2499__A0 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2500__A (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2501__A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2504__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__2505__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2506__A0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2507__A (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2508__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__2509__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__2510__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__2511__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__2512__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2513__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2514__A (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2515__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2518__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__2519__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2520__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2521__A (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2522__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__2523__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__2524__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__2525__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__2526__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2527__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2528__A (.DIODE(_1005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2529__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__2530__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__2531__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__2532__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__2533__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2534__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2535__B (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2536__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2539__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2540__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2541__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2542__A (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2543__A0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__2544__A0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__2545__A0 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__2546__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__2547__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2548__A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2549__B (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2550__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2553__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__2554__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2555__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2556__A (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2557__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__2558__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__2559__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__2560__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__2561__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2562__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2563__B (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2564__A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2565__A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2566__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__2567__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2568__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2569__A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2570__A (.DIODE(_1005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2571__A0 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__2572__A0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__2573__A0 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__2574__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__2575__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2576__A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2577__B (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2578__A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2579__A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2580__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__2581__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2582__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2583__A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2584__A (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2585__A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2586__A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2587__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__2588__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__2589__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2590__A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2591__A (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2592__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__2593__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__2594__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2595__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__2596__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2597__A1 (.DIODE(_1003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2598__A (.DIODE(_1085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2599__A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2600__A0 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__2601__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__2602__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__2603__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2604__A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2605__A (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2606__A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2607__A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2608__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__2609__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2610__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2611__A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2612__B (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2613__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__2614__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2616__A1 (.DIODE(_1001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2617__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2618__A1 (.DIODE(_1003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2619__A (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2620__A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2621__A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2622__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__2623__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2624__A0 (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2625__A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2626__B (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2627__A1 (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2628__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2630__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2631__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2632__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2633__A (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2634__A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2635__A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2636__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__2637__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2638__A0 (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2639__A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2640__A (.DIODE(_0994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2641__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__2642__A1 (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2644__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2645__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2646__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2647__A (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2648__A0 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__2649__A0 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__2650__A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2651__A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__2652__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__2653__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2655__A0 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__2656__A0 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2657__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__2658__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2659__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2660__A0 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2661__A (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2662__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__2663__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__2664__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__2665__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__2666__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2667__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__2671__B (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2672__B (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2674__A_N (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2675__B (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2676__B (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2678__A_N (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2679__B (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2680__B (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2681__B (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2682__A (.DIODE(\A[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2683__B1 (.DIODE(\A[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2685__B1_N (.DIODE(\A[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2687__A (.DIODE(\A[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2690__B (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2691__B (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2692__B (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2701__A (.DIODE(\A[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2701__B (.DIODE(_0796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2711__A2 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2715__A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__2716__A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__2720__A (.DIODE(\A[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2728__A0 (.DIODE(_0796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2728__A1 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA__2730__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__2730__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__2731__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__2731__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__2732__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2732__B1 (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2733__A1 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA__2733__C1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2747__A0 (.DIODE(_0848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2747__A1 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA__2749__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2749__B1 (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2750__A1 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA__2750__C1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2751__A0 (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2765__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2766__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2766__B1 (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2767__C1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2768__A0 (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2782__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2783__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2783__B1 (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2784__C1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2785__A0 (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2797__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2798__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2798__B1 (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2799__C1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2812__A0 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2814__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2814__B1 (.DIODE(_1264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2815__C1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2817__A1 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA__2826__A1 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA__2826__A2 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2826__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2827__C1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2828__A1 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA__2829__A2 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2829__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2830__C1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2833__A2 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2833__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2834__C1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2837__A2 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2837__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2838__C1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2841__A2 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2841__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2842__C1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2847__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2848__C1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2854__B (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__2855__A1 (.DIODE(net1086));
 sky130_fd_sc_hd__diode_2 ANTENNA__2855__C1 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2856__A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2859__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2860__C (.DIODE(\A[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2862__C1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2864__A1 (.DIODE(\A[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2865__A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__2866__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__2867__A (.DIODE(_0848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2867__B (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2867__C (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2868__C (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2868__D (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2869__A1 (.DIODE(_0796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2873__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2875__C1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2876__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2877__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2877__C1 (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2879__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__2881__A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__2882__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2884__A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2884__B1 (.DIODE(_0796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2884__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2885__B (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2887__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2887__A2 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2888__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2888__A2 (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2889__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2890__C1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__2891__A2_N (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2893__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2894__C1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2895__A2 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2895__B1 (.DIODE(_0897_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2899__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2901__C1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__2902__A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2902__B1 (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2902__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2906__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2908__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2908__A2 (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2908__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2910__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2912__A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2912__B1 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2912__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2916__A1 (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2918__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2918__B2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2921__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2922__C1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__2923__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2923__B2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2927__C1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__2928__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2928__B2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2930__B2 (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2933__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__2934__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2934__B2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2936__A1_N (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2939__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__2940__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2940__B2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__2943__A1 (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2946__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__2947__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2949__B2 (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2951__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__2953__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__2955__A (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2956__A0 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__2957__A0 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2958__A0 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__2959__A0 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__2960__A (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2961__A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2974__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__2974__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__2975__A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__2975__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__2976__A1 (.DIODE(\A[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2976__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__2977__A1 (.DIODE(\A[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2977__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__2978__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__2979__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__2980__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__2981__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__2982__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__2983__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__2984__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__2985__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__2986__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__2987__S (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__2988__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2989__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__2990__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__2991__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__2992__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2993__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3000__B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__3002__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3002__A2 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3003__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__3004__B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3020__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3022__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3041__B1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3042__B1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3044__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3045__B (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3046__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3048__B (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3049__D1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3050__C1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3055__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3057__C1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3058__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3058__B (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__3070__A2 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3071__C1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3073__B1 (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3076__B1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3082__D1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3091__B1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3095__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3099__A2 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3101__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3102__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3103__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3108__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3111__C1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3114__C1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3117__C1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3121__C1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3123__C1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3127__C1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3129__C1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3148__C1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3150__C1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3152__C1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3154__C1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3156__C1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3157__B (.DIODE(_0969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3168__C1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3170__C1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3172__C1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3174__C1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3176__C1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3178__C1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3180__C1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3184__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__3185__A (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3186__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3187__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3188__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3189__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3190__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3191__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3192__B (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3193__A0 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3195__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3196__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3197__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3198__A0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3199__A (.DIODE(_1089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3200__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3201__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3202__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3203__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3204__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3205__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3767__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__3768__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__3773__A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_wb_clk_i_A (.DIODE(clknet_3_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_wb_clk_i_A (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_wb_clk_i_A (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_wb_clk_i_A (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_wb_clk_i_A (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_wb_clk_i_A (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_wb_clk_i_A (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_wb_clk_i_A (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_wb_clk_i_A (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_wb_clk_i_A (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_wb_clk_i_A (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_wb_clk_i_A (.DIODE(clknet_3_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_wb_clk_i_A (.DIODE(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_wb_clk_i_A (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_wb_clk_i_A (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_wb_clk_i_A (.DIODE(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_wb_clk_i_A (.DIODE(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_wb_clk_i_A (.DIODE(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_wb_clk_i_A (.DIODE(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_wb_clk_i_A (.DIODE(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_wb_clk_i_A (.DIODE(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_wb_clk_i_A (.DIODE(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_wb_clk_i_A (.DIODE(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_wb_clk_i_A (.DIODE(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_wb_clk_i_A (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_wb_clk_i_A (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_wb_clk_i_A (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_wb_clk_i_A (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_wb_clk_i_A (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_wb_clk_i_A (.DIODE(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_wb_clk_i_A (.DIODE(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_wb_clk_i_A (.DIODE(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_wb_clk_i_A (.DIODE(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_wb_clk_i_A (.DIODE(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_wb_clk_i_A (.DIODE(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_wb_clk_i_A (.DIODE(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_wb_clk_i_A (.DIODE(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_wb_clk_i_A (.DIODE(clknet_3_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_wb_clk_i_A (.DIODE(clknet_3_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_wb_clk_i_A (.DIODE(clknet_3_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_wb_clk_i_A (.DIODE(clknet_3_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_wb_clk_i_A (.DIODE(clknet_3_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_wb_clk_i_A (.DIODE(clknet_3_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_wb_clk_i_A (.DIODE(clknet_3_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_wb_clk_i_A (.DIODE(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_wb_clk_i_A (.DIODE(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_wb_clk_i_A (.DIODE(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_wb_clk_i_A (.DIODE(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_wb_clk_i_A (.DIODE(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_wb_clk_i_A (.DIODE(clknet_3_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_wb_clk_i_A (.DIODE(clknet_3_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_wb_clk_i_A (.DIODE(clknet_3_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_57_wb_clk_i_A (.DIODE(clknet_3_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_wb_clk_i_A (.DIODE(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_wb_clk_i_A (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_wb_clk_i_A (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_wb_clk_i_A (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_wb_clk_i_A (.DIODE(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout103_A (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(\MAR[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(\MAR[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(\MAR[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(\MAR[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(\MAR[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(\MAR[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(\MAR[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(\MAR[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout71_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_A (.DIODE(_1003_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout73_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout74_A (.DIODE(_1003_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout76_A (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout78_A (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_A (.DIODE(_1001_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_A (.DIODE(_1001_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_A (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout87_A (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_A (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout89_A (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_A (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout91_A (.DIODE(_0999_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout93_A (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout94_A (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout95_A (.DIODE(_0998_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_A (.DIODE(_0993_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout97_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1021_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1033_A (.DIODE(\MAR[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1050_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold1062_A (.DIODE(\MAR[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold860_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold908_A (.DIODE(\A[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold918_A (.DIODE(\A[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold938_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold992_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold996_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_output19_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_output21_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_output23_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_output25_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_output27_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_output29_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_output36_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_output38_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_output40_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_output51_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_output53_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_output54_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_output61_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_output62_A (.DIODE(net62));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_90 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _1599_ (.A(net1191),
    .Y(_0540_));
 sky130_fd_sc_hd__inv_2 _1600_ (.A(net1147),
    .Y(_0541_));
 sky130_fd_sc_hd__inv_2 _1601_ (.A(net1090),
    .Y(_0542_));
 sky130_fd_sc_hd__inv_2 _1602_ (.A(net1088),
    .Y(_0543_));
 sky130_fd_sc_hd__inv_2 _1603_ (.A(net1234),
    .Y(_0544_));
 sky130_fd_sc_hd__clkinv_4 _1604_ (.A(net146),
    .Y(_0545_));
 sky130_fd_sc_hd__inv_2 _1605_ (.A(net1245),
    .Y(_0546_));
 sky130_fd_sc_hd__inv_2 _1606_ (.A(\A[5] ),
    .Y(_0547_));
 sky130_fd_sc_hd__inv_2 _1607_ (.A(\RAM[59][5] ),
    .Y(net29));
 sky130_fd_sc_hd__inv_2 _1608_ (.A(\RAM[59][4] ),
    .Y(net27));
 sky130_fd_sc_hd__inv_2 _1609_ (.A(\RAM[59][3] ),
    .Y(net25));
 sky130_fd_sc_hd__inv_2 _1610_ (.A(\RAM[59][2] ),
    .Y(net23));
 sky130_fd_sc_hd__inv_2 _1611_ (.A(\RAM[59][1] ),
    .Y(net21));
 sky130_fd_sc_hd__inv_2 _1612_ (.A(\RAM[59][0] ),
    .Y(net19));
 sky130_fd_sc_hd__inv_2 _1613_ (.A(\insin[0] ),
    .Y(_0548_));
 sky130_fd_sc_hd__inv_2 _1614_ (.A(net1160),
    .Y(_0549_));
 sky130_fd_sc_hd__inv_2 _1615_ (.A(net1184),
    .Y(_0550_));
 sky130_fd_sc_hd__inv_2 _1616_ (.A(net144),
    .Y(_0551_));
 sky130_fd_sc_hd__inv_2 _1617_ (.A(net1168),
    .Y(_0552_));
 sky130_fd_sc_hd__inv_2 _1618_ (.A(net1182),
    .Y(_0553_));
 sky130_fd_sc_hd__inv_2 _1619_ (.A(net1205),
    .Y(_0554_));
 sky130_fd_sc_hd__inv_2 _1620_ (.A(net156),
    .Y(_0555_));
 sky130_fd_sc_hd__inv_2 _1621_ (.A(net1094),
    .Y(_0556_));
 sky130_fd_sc_hd__inv_4 _1622_ (.A(net118),
    .Y(_0557_));
 sky130_fd_sc_hd__inv_2 _1623_ (.A(net116),
    .Y(_0558_));
 sky130_fd_sc_hd__inv_2 _1624_ (.A(\MAR[2] ),
    .Y(_0559_));
 sky130_fd_sc_hd__inv_2 _1625_ (.A(net131),
    .Y(_0560_));
 sky130_fd_sc_hd__inv_2 _1626_ (.A(net17),
    .Y(_0561_));
 sky130_fd_sc_hd__inv_2 _1627_ (.A(net997),
    .Y(_0562_));
 sky130_fd_sc_hd__or2_1 _1628_ (.A(net1107),
    .B(net1098),
    .X(_0563_));
 sky130_fd_sc_hd__nor4_1 _1629_ (.A(\ROM_spi_cycle[4] ),
    .B(\ROM_spi_cycle[1] ),
    .C(\ROM_spi_cycle[0] ),
    .D(_0563_),
    .Y(_0564_));
 sky130_fd_sc_hd__or4_1 _1630_ (.A(net1224),
    .B(net1231),
    .C(\ROM_spi_cycle[0] ),
    .D(_0563_),
    .X(_0565_));
 sky130_fd_sc_hd__or2_2 _1631_ (.A(net1234),
    .B(net1123),
    .X(_0566_));
 sky130_fd_sc_hd__or2_2 _1632_ (.A(net1007),
    .B(\startup_cycle[0] ),
    .X(_0567_));
 sky130_fd_sc_hd__or2_2 _1633_ (.A(_0566_),
    .B(_0567_),
    .X(_0568_));
 sky130_fd_sc_hd__or3_4 _1634_ (.A(net1090),
    .B(\startup_cycle[5] ),
    .C(net1088),
    .X(_0569_));
 sky130_fd_sc_hd__nor2_4 _1635_ (.A(_0568_),
    .B(_0569_),
    .Y(_0570_));
 sky130_fd_sc_hd__or2_4 _1636_ (.A(_0568_),
    .B(_0569_),
    .X(_0571_));
 sky130_fd_sc_hd__or3_2 _1637_ (.A(\mem_cycle[4] ),
    .B(\mem_cycle[3] ),
    .C(\mem_cycle[2] ),
    .X(_0572_));
 sky130_fd_sc_hd__or2_1 _1638_ (.A(net1195),
    .B(net1182),
    .X(_0573_));
 sky130_fd_sc_hd__or2_4 _1639_ (.A(_0572_),
    .B(_0573_),
    .X(_0574_));
 sky130_fd_sc_hd__nor3_4 _1640_ (.A(net106),
    .B(_0571_),
    .C(net1196),
    .Y(_0575_));
 sky130_fd_sc_hd__or3_4 _1641_ (.A(net106),
    .B(_0571_),
    .C(_0574_),
    .X(_0576_));
 sky130_fd_sc_hd__and3_1 _1642_ (.A(_0545_),
    .B(net144),
    .C(net149),
    .X(_0577_));
 sky130_fd_sc_hd__or2_2 _1643_ (.A(\insin[2] ),
    .B(net1239),
    .X(_0578_));
 sky130_fd_sc_hd__or3_2 _1644_ (.A(_0548_),
    .B(\insin[1] ),
    .C(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__or2_2 _1645_ (.A(_0550_),
    .B(net1080),
    .X(_0580_));
 sky130_fd_sc_hd__inv_2 _1646_ (.A(_0580_),
    .Y(_0581_));
 sky130_fd_sc_hd__nor2_1 _1647_ (.A(_0579_),
    .B(_0580_),
    .Y(_0582_));
 sky130_fd_sc_hd__or3_2 _1648_ (.A(\insin[0] ),
    .B(\insin[1] ),
    .C(_0578_),
    .X(_0583_));
 sky130_fd_sc_hd__nor3_1 _1649_ (.A(\insin[4] ),
    .B(net1080),
    .C(_0583_),
    .Y(_0584_));
 sky130_fd_sc_hd__nor2_1 _1650_ (.A(_0582_),
    .B(_0584_),
    .Y(_0585_));
 sky130_fd_sc_hd__and3b_1 _1651_ (.A_N(_0583_),
    .B(_0550_),
    .C(net1080),
    .X(_0586_));
 sky130_fd_sc_hd__or3b_2 _1652_ (.A(_0583_),
    .B(net1184),
    .C_N(net1080),
    .X(_0587_));
 sky130_fd_sc_hd__or4b_2 _1653_ (.A(\insin[2] ),
    .B(\insin[3] ),
    .C(_0580_),
    .D_N(\insin[1] ),
    .X(_0588_));
 sky130_fd_sc_hd__and3_1 _1654_ (.A(_0585_),
    .B(_0587_),
    .C(_0588_),
    .X(_0589_));
 sky130_fd_sc_hd__nor2_1 _1655_ (.A(_0550_),
    .B(_0583_),
    .Y(_0590_));
 sky130_fd_sc_hd__nand2_1 _1656_ (.A(net1160),
    .B(net1150),
    .Y(_0591_));
 sky130_fd_sc_hd__nand2_2 _1657_ (.A(_0548_),
    .B(\insin[1] ),
    .Y(_0592_));
 sky130_fd_sc_hd__a21oi_1 _1658_ (.A1(\insin[4] ),
    .A2(_0592_),
    .B1(_0591_),
    .Y(_0593_));
 sky130_fd_sc_hd__or3_1 _1659_ (.A(net1080),
    .B(_0590_),
    .C(_0593_),
    .X(_0594_));
 sky130_fd_sc_hd__nand2_2 _1660_ (.A(\insin[0] ),
    .B(\insin[1] ),
    .Y(_0595_));
 sky130_fd_sc_hd__or4_1 _1661_ (.A(\insin[4] ),
    .B(net1080),
    .C(_0591_),
    .D(_0595_),
    .X(_0596_));
 sky130_fd_sc_hd__nand2_1 _1662_ (.A(_0594_),
    .B(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__nand2_2 _1663_ (.A(\insin[4] ),
    .B(net1080),
    .Y(_0598_));
 sky130_fd_sc_hd__nor3_4 _1664_ (.A(_0578_),
    .B(_0592_),
    .C(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hd__or3_4 _1665_ (.A(_0578_),
    .B(_0592_),
    .C(_0598_),
    .X(_0600_));
 sky130_fd_sc_hd__or2_1 _1666_ (.A(_0579_),
    .B(_0598_),
    .X(_0601_));
 sky130_fd_sc_hd__nand3_1 _1667_ (.A(_0589_),
    .B(_0600_),
    .C(_0601_),
    .Y(_0602_));
 sky130_fd_sc_hd__a22o_1 _1668_ (.A1(_0589_),
    .A2(_0597_),
    .B1(_0602_),
    .B2(net1094),
    .X(_0603_));
 sky130_fd_sc_hd__nor2_1 _1669_ (.A(net146),
    .B(_0576_),
    .Y(_0604_));
 sky130_fd_sc_hd__nand2_4 _1670_ (.A(_0545_),
    .B(_0575_),
    .Y(_0605_));
 sky130_fd_sc_hd__and3_1 _1671_ (.A(net114),
    .B(net149),
    .C(_0604_),
    .X(_0606_));
 sky130_fd_sc_hd__and2b_1 _1672_ (.A_N(\insin[5] ),
    .B(_0593_),
    .X(_0607_));
 sky130_fd_sc_hd__nor3_1 _1673_ (.A(_0591_),
    .B(_0595_),
    .C(_0598_),
    .Y(_0608_));
 sky130_fd_sc_hd__inv_2 _1674_ (.A(_0608_),
    .Y(_0609_));
 sky130_fd_sc_hd__o21a_1 _1675_ (.A1(_0580_),
    .A2(_0583_),
    .B1(_0596_),
    .X(_0610_));
 sky130_fd_sc_hd__and3b_4 _1676_ (.A_N(_0607_),
    .B(_0609_),
    .C(_0610_),
    .X(_0611_));
 sky130_fd_sc_hd__or3b_4 _1677_ (.A(_0607_),
    .B(_0608_),
    .C_N(_0610_),
    .X(_0612_));
 sky130_fd_sc_hd__and2_1 _1678_ (.A(_0594_),
    .B(_0611_),
    .X(_0613_));
 sky130_fd_sc_hd__and3_1 _1679_ (.A(_0600_),
    .B(_0601_),
    .C(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__a31o_1 _1680_ (.A1(_0577_),
    .A2(_0587_),
    .A3(_0614_),
    .B1(_0576_),
    .X(_0615_));
 sky130_fd_sc_hd__a21o_1 _1681_ (.A1(net149),
    .A2(_0615_),
    .B1(_0606_),
    .X(_0616_));
 sky130_fd_sc_hd__a32o_1 _1682_ (.A1(_0575_),
    .A2(_0577_),
    .A3(_0603_),
    .B1(_0616_),
    .B2(net1094),
    .X(_0020_));
 sky130_fd_sc_hd__nand2b_1 _1683_ (.A_N(_0602_),
    .B(_0610_),
    .Y(_0617_));
 sky130_fd_sc_hd__a211o_1 _1684_ (.A1(net144),
    .A2(_0617_),
    .B1(_0576_),
    .C1(net1110),
    .X(_0618_));
 sky130_fd_sc_hd__nand2_1 _1685_ (.A(_0545_),
    .B(_0576_),
    .Y(_0619_));
 sky130_fd_sc_hd__a21o_1 _1686_ (.A1(_0618_),
    .A2(_0619_),
    .B1(net148),
    .X(_0021_));
 sky130_fd_sc_hd__o211a_1 _1687_ (.A1(net144),
    .A2(_0575_),
    .B1(net102),
    .C1(net149),
    .X(_0023_));
 sky130_fd_sc_hd__nand2_1 _1688_ (.A(net145),
    .B(_0588_),
    .Y(_0620_));
 sky130_fd_sc_hd__o2111a_1 _1689_ (.A1(_0550_),
    .A2(_0579_),
    .B1(_0587_),
    .C1(_0588_),
    .D1(net145),
    .X(_0621_));
 sky130_fd_sc_hd__nand2_1 _1690_ (.A(_0600_),
    .B(_0621_),
    .Y(_0622_));
 sky130_fd_sc_hd__nor2_1 _1691_ (.A(_0584_),
    .B(_0622_),
    .Y(_0623_));
 sky130_fd_sc_hd__a21o_1 _1692_ (.A1(_0610_),
    .A2(_0623_),
    .B1(_0576_),
    .X(_0624_));
 sky130_fd_sc_hd__o211a_1 _1693_ (.A1(net1110),
    .A2(_0575_),
    .B1(_0624_),
    .C1(net149),
    .X(_0022_));
 sky130_fd_sc_hd__nor2_1 _1694_ (.A(net146),
    .B(_0623_),
    .Y(_0625_));
 sky130_fd_sc_hd__o21ai_1 _1695_ (.A1(_0615_),
    .A2(_0625_),
    .B1(net1013),
    .Y(_0626_));
 sky130_fd_sc_hd__nor2_4 _1696_ (.A(net114),
    .B(_0599_),
    .Y(_0627_));
 sky130_fd_sc_hd__o21ai_1 _1697_ (.A1(_0580_),
    .A2(_0583_),
    .B1(_0627_),
    .Y(_0628_));
 sky130_fd_sc_hd__or4_1 _1698_ (.A(_0597_),
    .B(net102),
    .C(_0611_),
    .D(_0628_),
    .X(_0629_));
 sky130_fd_sc_hd__a21oi_1 _1699_ (.A1(net1014),
    .A2(_0629_),
    .B1(net148),
    .Y(_0019_));
 sky130_fd_sc_hd__o21bai_1 _1700_ (.A1(net146),
    .A2(_0621_),
    .B1_N(_0615_),
    .Y(_0630_));
 sky130_fd_sc_hd__or2_1 _1701_ (.A(_0584_),
    .B(_0599_),
    .X(_0631_));
 sky130_fd_sc_hd__a31o_1 _1702_ (.A1(net145),
    .A2(net1034),
    .A3(_0631_),
    .B1(net146),
    .X(_0632_));
 sky130_fd_sc_hd__a221o_1 _1703_ (.A1(net1034),
    .A2(_0630_),
    .B1(_0632_),
    .B2(_0575_),
    .C1(net148),
    .X(_0018_));
 sky130_fd_sc_hd__nor2_2 _1704_ (.A(ROM_spi_mode),
    .B(_0540_),
    .Y(net38));
 sky130_fd_sc_hd__or2_2 _1705_ (.A(ROM_spi_mode),
    .B(ROM_OEB),
    .X(net36));
 sky130_fd_sc_hd__nand2_1 _1706_ (.A(net1188),
    .B(net1182),
    .Y(_0633_));
 sky130_fd_sc_hd__or4b_4 _1707_ (.A(_0552_),
    .B(net1242),
    .C(_0633_),
    .D_N(net1178),
    .X(_0634_));
 sky130_fd_sc_hd__or2_1 _1708_ (.A(net1034),
    .B(_0571_),
    .X(_0635_));
 sky130_fd_sc_hd__or2_1 _1709_ (.A(_0634_),
    .B(_0635_),
    .X(_0636_));
 sky130_fd_sc_hd__or4_2 _1710_ (.A(net1094),
    .B(net1013),
    .C(net106),
    .D(_0636_),
    .X(_0637_));
 sky130_fd_sc_hd__and2_1 _1711_ (.A(net114),
    .B(\instr_cycle[1] ),
    .X(_0638_));
 sky130_fd_sc_hd__nand2_4 _1712_ (.A(net115),
    .B(net1110),
    .Y(_0639_));
 sky130_fd_sc_hd__or3_4 _1713_ (.A(_0550_),
    .B(_0583_),
    .C(_0639_),
    .X(_0640_));
 sky130_fd_sc_hd__nand2_4 _1714_ (.A(net117),
    .B(net116),
    .Y(_0641_));
 sky130_fd_sc_hd__nand2_2 _1715_ (.A(net123),
    .B(net119),
    .Y(_0642_));
 sky130_fd_sc_hd__or4_4 _1716_ (.A(net134),
    .B(net126),
    .C(_0641_),
    .D(_0642_),
    .X(_0643_));
 sky130_fd_sc_hd__mux4_1 _1717_ (.A0(\RAM[44][4] ),
    .A1(\RAM[45][4] ),
    .A2(\RAM[46][4] ),
    .A3(\RAM[47][4] ),
    .S0(net133),
    .S1(net125),
    .X(_0644_));
 sky130_fd_sc_hd__mux4_1 _1718_ (.A0(\RAM[40][4] ),
    .A1(\RAM[41][4] ),
    .A2(\RAM[42][4] ),
    .A3(\RAM[43][4] ),
    .S0(net133),
    .S1(net125),
    .X(_0645_));
 sky130_fd_sc_hd__mux4_1 _1719_ (.A0(\RAM[32][4] ),
    .A1(\RAM[33][4] ),
    .A2(\RAM[34][4] ),
    .A3(\RAM[35][4] ),
    .S0(net133),
    .S1(net125),
    .X(_0646_));
 sky130_fd_sc_hd__mux4_1 _1720_ (.A0(\RAM[36][4] ),
    .A1(\RAM[37][4] ),
    .A2(\RAM[38][4] ),
    .A3(\RAM[39][4] ),
    .S0(net133),
    .S1(net125),
    .X(_0647_));
 sky130_fd_sc_hd__mux4_2 _1721_ (.A0(_0646_),
    .A1(_0647_),
    .A2(_0645_),
    .A3(_0644_),
    .S0(net123),
    .S1(net119),
    .X(_0648_));
 sky130_fd_sc_hd__mux4_1 _1722_ (.A0(\RAM[12][4] ),
    .A1(\RAM[13][4] ),
    .A2(\RAM[14][4] ),
    .A3(\RAM[15][4] ),
    .S0(net140),
    .S1(net130),
    .X(_0649_));
 sky130_fd_sc_hd__mux2_1 _1723_ (.A0(\RAM[8][4] ),
    .A1(\RAM[9][4] ),
    .S(net140),
    .X(_0650_));
 sky130_fd_sc_hd__nand2_1 _1724_ (.A(net111),
    .B(_0650_),
    .Y(_0651_));
 sky130_fd_sc_hd__mux2_1 _1725_ (.A0(\RAM[10][4] ),
    .A1(\RAM[11][4] ),
    .S(net143),
    .X(_0652_));
 sky130_fd_sc_hd__nand2_1 _1726_ (.A(net130),
    .B(_0652_),
    .Y(_0653_));
 sky130_fd_sc_hd__o21ai_1 _1727_ (.A1(net112),
    .A2(_0649_),
    .B1(net121),
    .Y(_0654_));
 sky130_fd_sc_hd__a31o_1 _1728_ (.A1(net112),
    .A2(_0651_),
    .A3(_0653_),
    .B1(_0654_),
    .X(_0655_));
 sky130_fd_sc_hd__mux4_1 _1729_ (.A0(\RAM[4][4] ),
    .A1(\RAM[5][4] ),
    .A2(\RAM[6][4] ),
    .A3(\RAM[7][4] ),
    .S0(net141),
    .S1(net131),
    .X(_0656_));
 sky130_fd_sc_hd__nor2_1 _1730_ (.A(net112),
    .B(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__mux2_1 _1731_ (.A0(\RAM[2][4] ),
    .A1(\RAM[3][4] ),
    .S(net142),
    .X(_0658_));
 sky130_fd_sc_hd__nand2_1 _1732_ (.A(net131),
    .B(_0658_),
    .Y(_0659_));
 sky130_fd_sc_hd__mux2_1 _1733_ (.A0(\RAM[0][4] ),
    .A1(\RAM[1][4] ),
    .S(net141),
    .X(_0660_));
 sky130_fd_sc_hd__nand2_1 _1734_ (.A(net111),
    .B(_0660_),
    .Y(_0661_));
 sky130_fd_sc_hd__a311o_1 _1735_ (.A1(net112),
    .A2(_0659_),
    .A3(_0661_),
    .B1(net122),
    .C1(_0657_),
    .X(_0662_));
 sky130_fd_sc_hd__mux4_1 _1736_ (.A0(\RAM[24][4] ),
    .A1(\RAM[25][4] ),
    .A2(\RAM[26][4] ),
    .A3(\RAM[27][4] ),
    .S0(net135),
    .S1(net127),
    .X(_0663_));
 sky130_fd_sc_hd__mux4_1 _1737_ (.A0(\RAM[28][4] ),
    .A1(\RAM[29][4] ),
    .A2(\RAM[30][4] ),
    .A3(\RAM[31][4] ),
    .S0(net135),
    .S1(net127),
    .X(_0664_));
 sky130_fd_sc_hd__mux4_1 _1738_ (.A0(\RAM[20][4] ),
    .A1(\RAM[21][4] ),
    .A2(\RAM[22][4] ),
    .A3(\RAM[23][4] ),
    .S0(net135),
    .S1(net127),
    .X(_0665_));
 sky130_fd_sc_hd__mux4_1 _1739_ (.A0(\RAM[16][4] ),
    .A1(\RAM[17][4] ),
    .A2(\RAM[18][4] ),
    .A3(\RAM[19][4] ),
    .S0(net136),
    .S1(net128),
    .X(_0666_));
 sky130_fd_sc_hd__mux4_2 _1740_ (.A0(_0666_),
    .A1(_0665_),
    .A2(_0663_),
    .A3(_0664_),
    .S0(net124),
    .S1(net120),
    .X(_0667_));
 sky130_fd_sc_hd__mux4_1 _1741_ (.A0(net50),
    .A1(\RAM[61][4] ),
    .A2(\RAM[62][4] ),
    .A3(net44),
    .S0(net138),
    .S1(net129),
    .X(_0668_));
 sky130_fd_sc_hd__mux2_1 _1742_ (.A0(\RAM[56][4] ),
    .A1(\RAM[57][4] ),
    .S(net141),
    .X(_0669_));
 sky130_fd_sc_hd__nand2_1 _1743_ (.A(net110),
    .B(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__nor2_1 _1744_ (.A(net59),
    .B(net141),
    .Y(_0671_));
 sky130_fd_sc_hd__a211o_1 _1745_ (.A1(net27),
    .A2(net138),
    .B1(net110),
    .C1(_0671_),
    .X(_0672_));
 sky130_fd_sc_hd__o21ai_1 _1746_ (.A1(net113),
    .A2(_0668_),
    .B1(net121),
    .Y(_0673_));
 sky130_fd_sc_hd__a31o_1 _1747_ (.A1(net113),
    .A2(_0670_),
    .A3(_0672_),
    .B1(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__mux4_1 _1748_ (.A0(\RAM[48][4] ),
    .A1(\RAM[49][4] ),
    .A2(\RAM[50][4] ),
    .A3(\RAM[51][4] ),
    .S0(net137),
    .S1(net129),
    .X(_0675_));
 sky130_fd_sc_hd__nor2_1 _1749_ (.A(net123),
    .B(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__mux2_1 _1750_ (.A0(\RAM[54][4] ),
    .A1(\RAM[55][4] ),
    .S(net140),
    .X(_0677_));
 sky130_fd_sc_hd__nand2_1 _1751_ (.A(net130),
    .B(_0677_),
    .Y(_0678_));
 sky130_fd_sc_hd__mux2_1 _1752_ (.A0(\RAM[52][4] ),
    .A1(\RAM[53][4] ),
    .S(net140),
    .X(_0679_));
 sky130_fd_sc_hd__nand2_1 _1753_ (.A(net110),
    .B(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__a311o_1 _1754_ (.A1(net124),
    .A2(_0678_),
    .A3(_0680_),
    .B1(net119),
    .C1(_0676_),
    .X(_0681_));
 sky130_fd_sc_hd__nor2_1 _1755_ (.A(_0557_),
    .B(_0667_),
    .Y(_0682_));
 sky130_fd_sc_hd__a31o_1 _1756_ (.A1(_0557_),
    .A2(_0655_),
    .A3(_0662_),
    .B1(net116),
    .X(_0683_));
 sky130_fd_sc_hd__o21ai_1 _1757_ (.A1(net118),
    .A2(_0648_),
    .B1(net116),
    .Y(_0684_));
 sky130_fd_sc_hd__a31o_1 _1758_ (.A1(net117),
    .A2(_0674_),
    .A3(_0681_),
    .B1(_0684_),
    .X(_0685_));
 sky130_fd_sc_hd__o211ai_1 _1759_ (.A1(_0682_),
    .A2(_0683_),
    .B1(_0685_),
    .C1(net105),
    .Y(_0686_));
 sky130_fd_sc_hd__nand2_1 _1760_ (.A(net134),
    .B(net126),
    .Y(_0687_));
 sky130_fd_sc_hd__nor3_4 _1761_ (.A(_0641_),
    .B(_0642_),
    .C(_0687_),
    .Y(_0688_));
 sky130_fd_sc_hd__or3_4 _1762_ (.A(_0641_),
    .B(_0642_),
    .C(_0687_),
    .X(_0689_));
 sky130_fd_sc_hd__o211a_1 _1763_ (.A1(net10),
    .A2(net105),
    .B1(_0686_),
    .C1(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__a21o_1 _1764_ (.A1(net4),
    .A2(_0688_),
    .B1(_0612_),
    .X(_0691_));
 sky130_fd_sc_hd__o22a_4 _1765_ (.A1(net1001),
    .A2(_0611_),
    .B1(_0690_),
    .B2(_0691_),
    .X(_0692_));
 sky130_fd_sc_hd__nor2_2 _1766_ (.A(net114),
    .B(_0600_),
    .Y(_0693_));
 sky130_fd_sc_hd__nand2_2 _1767_ (.A(net145),
    .B(_0599_),
    .Y(_0694_));
 sky130_fd_sc_hd__o22a_1 _1768_ (.A1(_0640_),
    .A2(_0692_),
    .B1(net103),
    .B2(net945),
    .X(_0695_));
 sky130_fd_sc_hd__a21oi_4 _1769_ (.A1(_0640_),
    .A2(net103),
    .B1(net102),
    .Y(_0696_));
 sky130_fd_sc_hd__o22a_1 _1770_ (.A1(net102),
    .A2(_0695_),
    .B1(_0696_),
    .B2(net1241),
    .X(_0697_));
 sky130_fd_sc_hd__mux2_1 _1771_ (.A0(net13),
    .A1(_0697_),
    .S(_0637_),
    .X(_0698_));
 sky130_fd_sc_hd__and2_1 _1772_ (.A(net149),
    .B(_0698_),
    .X(_0010_));
 sky130_fd_sc_hd__mux4_1 _1773_ (.A0(\RAM[44][5] ),
    .A1(\RAM[45][5] ),
    .A2(\RAM[46][5] ),
    .A3(\RAM[47][5] ),
    .S0(net133),
    .S1(net127),
    .X(_0699_));
 sky130_fd_sc_hd__mux4_2 _1774_ (.A0(\RAM[40][5] ),
    .A1(\RAM[41][5] ),
    .A2(\RAM[42][5] ),
    .A3(\RAM[43][5] ),
    .S0(net133),
    .S1(net125),
    .X(_0700_));
 sky130_fd_sc_hd__mux4_1 _1775_ (.A0(\RAM[32][5] ),
    .A1(\RAM[33][5] ),
    .A2(\RAM[34][5] ),
    .A3(\RAM[35][5] ),
    .S0(net135),
    .S1(net127),
    .X(_0701_));
 sky130_fd_sc_hd__mux4_1 _1776_ (.A0(\RAM[36][5] ),
    .A1(\RAM[37][5] ),
    .A2(\RAM[38][5] ),
    .A3(\RAM[39][5] ),
    .S0(net133),
    .S1(net125),
    .X(_0702_));
 sky130_fd_sc_hd__mux4_1 _1777_ (.A0(_0701_),
    .A1(_0702_),
    .A2(_0700_),
    .A3(_0699_),
    .S0(net123),
    .S1(net119),
    .X(_0703_));
 sky130_fd_sc_hd__mux4_1 _1778_ (.A0(\RAM[12][5] ),
    .A1(\RAM[13][5] ),
    .A2(\RAM[14][5] ),
    .A3(\RAM[15][5] ),
    .S0(net143),
    .S1(net130),
    .X(_0704_));
 sky130_fd_sc_hd__mux2_1 _1779_ (.A0(\RAM[8][5] ),
    .A1(\RAM[9][5] ),
    .S(net140),
    .X(_0705_));
 sky130_fd_sc_hd__mux2_1 _1780_ (.A0(\RAM[10][5] ),
    .A1(\RAM[11][5] ),
    .S(net140),
    .X(_0706_));
 sky130_fd_sc_hd__a21o_1 _1781_ (.A1(net130),
    .A2(_0706_),
    .B1(net124),
    .X(_0707_));
 sky130_fd_sc_hd__a21o_1 _1782_ (.A1(net111),
    .A2(_0705_),
    .B1(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__o211ai_1 _1783_ (.A1(net112),
    .A2(_0704_),
    .B1(_0708_),
    .C1(net121),
    .Y(_0709_));
 sky130_fd_sc_hd__mux4_1 _1784_ (.A0(\RAM[4][5] ),
    .A1(\RAM[5][5] ),
    .A2(\RAM[6][5] ),
    .A3(\RAM[7][5] ),
    .S0(net141),
    .S1(net131),
    .X(_0710_));
 sky130_fd_sc_hd__nor2_1 _1785_ (.A(_0559_),
    .B(_0710_),
    .Y(_0711_));
 sky130_fd_sc_hd__mux2_1 _1786_ (.A0(\RAM[2][5] ),
    .A1(\RAM[3][5] ),
    .S(net142),
    .X(_0712_));
 sky130_fd_sc_hd__mux2_1 _1787_ (.A0(\RAM[0][5] ),
    .A1(\RAM[1][5] ),
    .S(net141),
    .X(_0713_));
 sky130_fd_sc_hd__a21o_1 _1788_ (.A1(net111),
    .A2(_0713_),
    .B1(\MAR[2] ),
    .X(_0714_));
 sky130_fd_sc_hd__a21oi_1 _1789_ (.A1(net130),
    .A2(_0712_),
    .B1(_0714_),
    .Y(_0715_));
 sky130_fd_sc_hd__mux4_1 _1790_ (.A0(\RAM[24][5] ),
    .A1(\RAM[25][5] ),
    .A2(\RAM[26][5] ),
    .A3(\RAM[27][5] ),
    .S0(net135),
    .S1(net127),
    .X(_0716_));
 sky130_fd_sc_hd__mux4_1 _1791_ (.A0(\RAM[28][5] ),
    .A1(\RAM[29][5] ),
    .A2(\RAM[30][5] ),
    .A3(\RAM[31][5] ),
    .S0(net135),
    .S1(net127),
    .X(_0717_));
 sky130_fd_sc_hd__mux4_1 _1792_ (.A0(\RAM[20][5] ),
    .A1(\RAM[21][5] ),
    .A2(\RAM[22][5] ),
    .A3(\RAM[23][5] ),
    .S0(net135),
    .S1(net127),
    .X(_0718_));
 sky130_fd_sc_hd__mux4_1 _1793_ (.A0(\RAM[16][5] ),
    .A1(\RAM[17][5] ),
    .A2(\RAM[18][5] ),
    .A3(\RAM[19][5] ),
    .S0(net136),
    .S1(net128),
    .X(_0719_));
 sky130_fd_sc_hd__mux4_1 _1794_ (.A0(_0719_),
    .A1(_0718_),
    .A2(_0716_),
    .A3(_0717_),
    .S0(net124),
    .S1(net120),
    .X(_0720_));
 sky130_fd_sc_hd__mux4_1 _1795_ (.A0(net52),
    .A1(\RAM[61][5] ),
    .A2(\RAM[62][5] ),
    .A3(net45),
    .S0(net138),
    .S1(net132),
    .X(_0721_));
 sky130_fd_sc_hd__mux2_1 _1796_ (.A0(\RAM[56][5] ),
    .A1(\RAM[57][5] ),
    .S(net138),
    .X(_0722_));
 sky130_fd_sc_hd__nand2_1 _1797_ (.A(net110),
    .B(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__nor2_1 _1798_ (.A(net60),
    .B(net138),
    .Y(_0724_));
 sky130_fd_sc_hd__a211o_1 _1799_ (.A1(net29),
    .A2(net138),
    .B1(net110),
    .C1(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__o21ai_1 _1800_ (.A1(net113),
    .A2(_0721_),
    .B1(net121),
    .Y(_0726_));
 sky130_fd_sc_hd__a31o_1 _1801_ (.A1(net113),
    .A2(_0723_),
    .A3(_0725_),
    .B1(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__mux4_1 _1802_ (.A0(\RAM[48][5] ),
    .A1(\RAM[49][5] ),
    .A2(\RAM[50][5] ),
    .A3(\RAM[51][5] ),
    .S0(net137),
    .S1(net129),
    .X(_0728_));
 sky130_fd_sc_hd__nor2_1 _1803_ (.A(net123),
    .B(_0728_),
    .Y(_0729_));
 sky130_fd_sc_hd__mux2_1 _1804_ (.A0(\RAM[54][5] ),
    .A1(\RAM[55][5] ),
    .S(net140),
    .X(_0730_));
 sky130_fd_sc_hd__nand2_1 _1805_ (.A(net130),
    .B(_0730_),
    .Y(_0731_));
 sky130_fd_sc_hd__mux2_1 _1806_ (.A0(\RAM[52][5] ),
    .A1(\RAM[53][5] ),
    .S(net140),
    .X(_0732_));
 sky130_fd_sc_hd__nand2_1 _1807_ (.A(net110),
    .B(_0732_),
    .Y(_0733_));
 sky130_fd_sc_hd__a311o_1 _1808_ (.A1(\MAR[2] ),
    .A2(_0731_),
    .A3(_0733_),
    .B1(net122),
    .C1(_0729_),
    .X(_0734_));
 sky130_fd_sc_hd__o311a_1 _1809_ (.A1(net121),
    .A2(_0711_),
    .A3(_0715_),
    .B1(_0709_),
    .C1(_0557_),
    .X(_0735_));
 sky130_fd_sc_hd__o21ai_1 _1810_ (.A1(_0557_),
    .A2(_0720_),
    .B1(_0558_),
    .Y(_0736_));
 sky130_fd_sc_hd__o21ai_1 _1811_ (.A1(net117),
    .A2(_0703_),
    .B1(net116),
    .Y(_0737_));
 sky130_fd_sc_hd__a31o_1 _1812_ (.A1(net117),
    .A2(_0727_),
    .A3(_0734_),
    .B1(_0737_),
    .X(_0738_));
 sky130_fd_sc_hd__o211ai_1 _1813_ (.A1(_0735_),
    .A2(_0736_),
    .B1(_0738_),
    .C1(net105),
    .Y(_0739_));
 sky130_fd_sc_hd__o211a_1 _1814_ (.A1(net11),
    .A2(net105),
    .B1(_0689_),
    .C1(_0739_),
    .X(_0740_));
 sky130_fd_sc_hd__a21o_1 _1815_ (.A1(net5),
    .A2(_0688_),
    .B1(_0612_),
    .X(_0741_));
 sky130_fd_sc_hd__o22a_4 _1816_ (.A1(net1011),
    .A2(_0611_),
    .B1(_0740_),
    .B2(_0741_),
    .X(_0742_));
 sky130_fd_sc_hd__o22a_1 _1817_ (.A1(net553),
    .A2(net103),
    .B1(_0742_),
    .B2(_0640_),
    .X(_0743_));
 sky130_fd_sc_hd__o22ai_1 _1818_ (.A1(net1186),
    .A2(_0696_),
    .B1(_0743_),
    .B2(net102),
    .Y(_0744_));
 sky130_fd_sc_hd__nand2_1 _1819_ (.A(_0637_),
    .B(_0744_),
    .Y(_0745_));
 sky130_fd_sc_hd__o211a_1 _1820_ (.A1(net14),
    .A2(_0637_),
    .B1(_0745_),
    .C1(net149),
    .X(_0011_));
 sky130_fd_sc_hd__and3_2 _1821_ (.A(net1168),
    .B(net1178),
    .C(net1205),
    .X(_0746_));
 sky130_fd_sc_hd__or3b_4 _1822_ (.A(net1188),
    .B(_0553_),
    .C_N(_0746_),
    .X(_0747_));
 sky130_fd_sc_hd__or2_1 _1823_ (.A(_0635_),
    .B(_0747_),
    .X(_0748_));
 sky130_fd_sc_hd__or4_4 _1824_ (.A(net1094),
    .B(net1013),
    .C(net106),
    .D(_0748_),
    .X(_0749_));
 sky130_fd_sc_hd__mux4_1 _1825_ (.A0(\RAM[44][0] ),
    .A1(\RAM[45][0] ),
    .A2(\RAM[46][0] ),
    .A3(\RAM[47][0] ),
    .S0(net133),
    .S1(net125),
    .X(_0750_));
 sky130_fd_sc_hd__mux4_1 _1826_ (.A0(\RAM[40][0] ),
    .A1(\RAM[41][0] ),
    .A2(\RAM[42][0] ),
    .A3(\RAM[43][0] ),
    .S0(net133),
    .S1(net125),
    .X(_0751_));
 sky130_fd_sc_hd__mux4_1 _1827_ (.A0(\RAM[32][0] ),
    .A1(\RAM[33][0] ),
    .A2(\RAM[34][0] ),
    .A3(\RAM[35][0] ),
    .S0(net134),
    .S1(net126),
    .X(_0752_));
 sky130_fd_sc_hd__mux4_1 _1828_ (.A0(\RAM[36][0] ),
    .A1(\RAM[37][0] ),
    .A2(\RAM[38][0] ),
    .A3(\RAM[39][0] ),
    .S0(net134),
    .S1(net126),
    .X(_0753_));
 sky130_fd_sc_hd__mux4_1 _1829_ (.A0(_0752_),
    .A1(_0753_),
    .A2(_0751_),
    .A3(_0750_),
    .S0(net123),
    .S1(net119),
    .X(_0754_));
 sky130_fd_sc_hd__mux4_1 _1830_ (.A0(\RAM[12][0] ),
    .A1(\RAM[13][0] ),
    .A2(\RAM[14][0] ),
    .A3(\RAM[15][0] ),
    .S0(net140),
    .S1(net130),
    .X(_0755_));
 sky130_fd_sc_hd__mux2_1 _1831_ (.A0(\RAM[8][0] ),
    .A1(\RAM[9][0] ),
    .S(net140),
    .X(_0756_));
 sky130_fd_sc_hd__nand2_1 _1832_ (.A(net110),
    .B(_0756_),
    .Y(_0757_));
 sky130_fd_sc_hd__mux2_1 _1833_ (.A0(\RAM[10][0] ),
    .A1(\RAM[11][0] ),
    .S(net140),
    .X(_0758_));
 sky130_fd_sc_hd__nand2_1 _1834_ (.A(net130),
    .B(_0758_),
    .Y(_0759_));
 sky130_fd_sc_hd__o21ai_1 _1835_ (.A1(net112),
    .A2(_0755_),
    .B1(net121),
    .Y(_0760_));
 sky130_fd_sc_hd__a31o_1 _1836_ (.A1(net112),
    .A2(_0757_),
    .A3(_0759_),
    .B1(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__mux4_1 _1837_ (.A0(\RAM[4][0] ),
    .A1(\RAM[5][0] ),
    .A2(\RAM[6][0] ),
    .A3(\RAM[7][0] ),
    .S0(net141),
    .S1(net131),
    .X(_0762_));
 sky130_fd_sc_hd__nor2_1 _1838_ (.A(net112),
    .B(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__mux2_1 _1839_ (.A0(\RAM[2][0] ),
    .A1(\RAM[3][0] ),
    .S(net141),
    .X(_0764_));
 sky130_fd_sc_hd__nand2_1 _1840_ (.A(net131),
    .B(_0764_),
    .Y(_0765_));
 sky130_fd_sc_hd__mux2_1 _1841_ (.A0(\RAM[0][0] ),
    .A1(\RAM[1][0] ),
    .S(net141),
    .X(_0766_));
 sky130_fd_sc_hd__nand2_1 _1842_ (.A(net111),
    .B(_0766_),
    .Y(_0767_));
 sky130_fd_sc_hd__a311o_1 _1843_ (.A1(_0559_),
    .A2(_0765_),
    .A3(_0767_),
    .B1(net122),
    .C1(_0763_),
    .X(_0768_));
 sky130_fd_sc_hd__mux4_1 _1844_ (.A0(\RAM[24][0] ),
    .A1(\RAM[25][0] ),
    .A2(\RAM[26][0] ),
    .A3(\RAM[27][0] ),
    .S0(net135),
    .S1(net127),
    .X(_0769_));
 sky130_fd_sc_hd__mux4_1 _1845_ (.A0(\RAM[28][0] ),
    .A1(\RAM[29][0] ),
    .A2(\RAM[30][0] ),
    .A3(\RAM[31][0] ),
    .S0(net135),
    .S1(net127),
    .X(_0770_));
 sky130_fd_sc_hd__mux4_1 _1846_ (.A0(\RAM[20][0] ),
    .A1(\RAM[21][0] ),
    .A2(\RAM[22][0] ),
    .A3(\RAM[23][0] ),
    .S0(net136),
    .S1(net128),
    .X(_0771_));
 sky130_fd_sc_hd__mux4_1 _1847_ (.A0(\RAM[16][0] ),
    .A1(\RAM[17][0] ),
    .A2(\RAM[18][0] ),
    .A3(\RAM[19][0] ),
    .S0(net136),
    .S1(net128),
    .X(_0772_));
 sky130_fd_sc_hd__mux4_1 _1848_ (.A0(_0772_),
    .A1(_0771_),
    .A2(_0769_),
    .A3(_0770_),
    .S0(net124),
    .S1(net120),
    .X(_0773_));
 sky130_fd_sc_hd__mux4_1 _1849_ (.A0(net46),
    .A1(\RAM[61][0] ),
    .A2(\RAM[62][0] ),
    .A3(net69),
    .S0(net139),
    .S1(net132),
    .X(_0774_));
 sky130_fd_sc_hd__mux2_1 _1850_ (.A0(\RAM[56][0] ),
    .A1(\RAM[57][0] ),
    .S(net139),
    .X(_0775_));
 sky130_fd_sc_hd__nand2_1 _1851_ (.A(net110),
    .B(_0775_),
    .Y(_0776_));
 sky130_fd_sc_hd__nor2_1 _1852_ (.A(net55),
    .B(net138),
    .Y(_0777_));
 sky130_fd_sc_hd__a211o_1 _1853_ (.A1(net19),
    .A2(net138),
    .B1(net110),
    .C1(_0777_),
    .X(_0778_));
 sky130_fd_sc_hd__o21ai_1 _1854_ (.A1(net113),
    .A2(_0774_),
    .B1(net121),
    .Y(_0779_));
 sky130_fd_sc_hd__a31o_1 _1855_ (.A1(net113),
    .A2(_0776_),
    .A3(_0778_),
    .B1(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__mux4_1 _1856_ (.A0(\RAM[48][0] ),
    .A1(\RAM[49][0] ),
    .A2(\RAM[50][0] ),
    .A3(\RAM[51][0] ),
    .S0(net137),
    .S1(net129),
    .X(_0781_));
 sky130_fd_sc_hd__nor2_1 _1857_ (.A(net124),
    .B(_0781_),
    .Y(_0782_));
 sky130_fd_sc_hd__mux2_1 _1858_ (.A0(\RAM[54][0] ),
    .A1(\RAM[55][0] ),
    .S(net137),
    .X(_0783_));
 sky130_fd_sc_hd__nand2_1 _1859_ (.A(net129),
    .B(_0783_),
    .Y(_0784_));
 sky130_fd_sc_hd__mux2_1 _1860_ (.A0(\RAM[52][0] ),
    .A1(\RAM[53][0] ),
    .S(net137),
    .X(_0785_));
 sky130_fd_sc_hd__nand2_1 _1861_ (.A(net110),
    .B(_0785_),
    .Y(_0786_));
 sky130_fd_sc_hd__a311o_1 _1862_ (.A1(net124),
    .A2(_0784_),
    .A3(_0786_),
    .B1(net119),
    .C1(_0782_),
    .X(_0787_));
 sky130_fd_sc_hd__o21ai_1 _1863_ (.A1(_0557_),
    .A2(_0773_),
    .B1(_0558_),
    .Y(_0788_));
 sky130_fd_sc_hd__a31o_1 _1864_ (.A1(_0557_),
    .A2(_0761_),
    .A3(_0768_),
    .B1(_0788_),
    .X(_0789_));
 sky130_fd_sc_hd__o21ai_1 _1865_ (.A1(net117),
    .A2(_0754_),
    .B1(net116),
    .Y(_0790_));
 sky130_fd_sc_hd__a31o_1 _1866_ (.A1(net117),
    .A2(_0780_),
    .A3(_0787_),
    .B1(_0790_),
    .X(_0791_));
 sky130_fd_sc_hd__and3_1 _1867_ (.A(net105),
    .B(_0789_),
    .C(_0791_),
    .X(_0792_));
 sky130_fd_sc_hd__o21ai_2 _1868_ (.A1(net6),
    .A2(net105),
    .B1(_0689_),
    .Y(_0793_));
 sky130_fd_sc_hd__o221ai_4 _1869_ (.A1(_0561_),
    .A2(_0689_),
    .B1(_0792_),
    .B2(_0793_),
    .C1(_0611_),
    .Y(_0794_));
 sky130_fd_sc_hd__or2_1 _1870_ (.A(net601),
    .B(_0611_),
    .X(_0795_));
 sky130_fd_sc_hd__and2_4 _1871_ (.A(_0794_),
    .B(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__o22a_1 _1872_ (.A1(net417),
    .A2(net103),
    .B1(_0796_),
    .B2(_0640_),
    .X(_0797_));
 sky130_fd_sc_hd__o22a_1 _1873_ (.A1(net1247),
    .A2(_0696_),
    .B1(_0797_),
    .B2(net102),
    .X(_0798_));
 sky130_fd_sc_hd__mux2_1 _1874_ (.A0(net13),
    .A1(_0798_),
    .S(_0749_),
    .X(_0799_));
 sky130_fd_sc_hd__and2_1 _1875_ (.A(net149),
    .B(_0799_),
    .X(_0006_));
 sky130_fd_sc_hd__mux4_1 _1876_ (.A0(\RAM[44][1] ),
    .A1(\RAM[45][1] ),
    .A2(\RAM[46][1] ),
    .A3(\RAM[47][1] ),
    .S0(net134),
    .S1(net125),
    .X(_0800_));
 sky130_fd_sc_hd__mux4_1 _1877_ (.A0(\RAM[40][1] ),
    .A1(\RAM[41][1] ),
    .A2(\RAM[42][1] ),
    .A3(\RAM[43][1] ),
    .S0(net133),
    .S1(net125),
    .X(_0801_));
 sky130_fd_sc_hd__mux4_1 _1878_ (.A0(\RAM[32][1] ),
    .A1(\RAM[33][1] ),
    .A2(\RAM[34][1] ),
    .A3(\RAM[35][1] ),
    .S0(net133),
    .S1(net125),
    .X(_0802_));
 sky130_fd_sc_hd__mux4_1 _1879_ (.A0(\RAM[36][1] ),
    .A1(\RAM[37][1] ),
    .A2(\RAM[38][1] ),
    .A3(\RAM[39][1] ),
    .S0(net133),
    .S1(net125),
    .X(_0803_));
 sky130_fd_sc_hd__mux4_1 _1880_ (.A0(_0802_),
    .A1(_0803_),
    .A2(_0801_),
    .A3(_0800_),
    .S0(net123),
    .S1(net119),
    .X(_0804_));
 sky130_fd_sc_hd__mux4_1 _1881_ (.A0(\RAM[12][1] ),
    .A1(\RAM[13][1] ),
    .A2(\RAM[14][1] ),
    .A3(\RAM[15][1] ),
    .S0(net143),
    .S1(net130),
    .X(_0805_));
 sky130_fd_sc_hd__mux2_1 _1882_ (.A0(\RAM[8][1] ),
    .A1(\RAM[9][1] ),
    .S(net143),
    .X(_0806_));
 sky130_fd_sc_hd__nand2_1 _1883_ (.A(net111),
    .B(_0806_),
    .Y(_0807_));
 sky130_fd_sc_hd__mux2_1 _1884_ (.A0(\RAM[10][1] ),
    .A1(\RAM[11][1] ),
    .S(net140),
    .X(_0808_));
 sky130_fd_sc_hd__nand2_1 _1885_ (.A(net130),
    .B(_0808_),
    .Y(_0809_));
 sky130_fd_sc_hd__o21ai_1 _1886_ (.A1(net112),
    .A2(_0805_),
    .B1(net121),
    .Y(_0810_));
 sky130_fd_sc_hd__a31o_1 _1887_ (.A1(net112),
    .A2(_0807_),
    .A3(_0809_),
    .B1(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__mux4_1 _1888_ (.A0(\RAM[4][1] ),
    .A1(\RAM[5][1] ),
    .A2(\RAM[6][1] ),
    .A3(\RAM[7][1] ),
    .S0(net142),
    .S1(net131),
    .X(_0812_));
 sky130_fd_sc_hd__nor2_1 _1889_ (.A(net112),
    .B(_0812_),
    .Y(_0813_));
 sky130_fd_sc_hd__mux2_1 _1890_ (.A0(\RAM[2][1] ),
    .A1(\RAM[3][1] ),
    .S(net141),
    .X(_0814_));
 sky130_fd_sc_hd__nand2_1 _1891_ (.A(net131),
    .B(_0814_),
    .Y(_0815_));
 sky130_fd_sc_hd__mux2_1 _1892_ (.A0(\RAM[0][1] ),
    .A1(\RAM[1][1] ),
    .S(net142),
    .X(_0816_));
 sky130_fd_sc_hd__nand2_1 _1893_ (.A(net111),
    .B(_0816_),
    .Y(_0817_));
 sky130_fd_sc_hd__a311o_1 _1894_ (.A1(net112),
    .A2(_0815_),
    .A3(_0817_),
    .B1(net122),
    .C1(_0813_),
    .X(_0818_));
 sky130_fd_sc_hd__mux4_1 _1895_ (.A0(\RAM[24][1] ),
    .A1(\RAM[25][1] ),
    .A2(\RAM[26][1] ),
    .A3(\RAM[27][1] ),
    .S0(net135),
    .S1(net127),
    .X(_0819_));
 sky130_fd_sc_hd__mux4_1 _1896_ (.A0(\RAM[28][1] ),
    .A1(\RAM[29][1] ),
    .A2(\RAM[30][1] ),
    .A3(\RAM[31][1] ),
    .S0(net135),
    .S1(net127),
    .X(_0820_));
 sky130_fd_sc_hd__mux4_1 _1897_ (.A0(\RAM[20][1] ),
    .A1(\RAM[21][1] ),
    .A2(\RAM[22][1] ),
    .A3(\RAM[23][1] ),
    .S0(net135),
    .S1(net127),
    .X(_0821_));
 sky130_fd_sc_hd__mux4_1 _1898_ (.A0(\RAM[16][1] ),
    .A1(\RAM[17][1] ),
    .A2(\RAM[18][1] ),
    .A3(\RAM[19][1] ),
    .S0(net136),
    .S1(net128),
    .X(_0822_));
 sky130_fd_sc_hd__mux4_1 _1899_ (.A0(_0822_),
    .A1(_0821_),
    .A2(_0819_),
    .A3(_0820_),
    .S0(net124),
    .S1(net120),
    .X(_0823_));
 sky130_fd_sc_hd__mux4_1 _1900_ (.A0(net47),
    .A1(\RAM[61][1] ),
    .A2(\RAM[62][1] ),
    .A3(net41),
    .S0(net139),
    .S1(net129),
    .X(_0824_));
 sky130_fd_sc_hd__mux2_1 _1901_ (.A0(\RAM[56][1] ),
    .A1(\RAM[57][1] ),
    .S(net138),
    .X(_0825_));
 sky130_fd_sc_hd__nand2_1 _1902_ (.A(net110),
    .B(_0825_),
    .Y(_0826_));
 sky130_fd_sc_hd__nor2_1 _1903_ (.A(net56),
    .B(net138),
    .Y(_0827_));
 sky130_fd_sc_hd__a211o_1 _1904_ (.A1(net21),
    .A2(net138),
    .B1(net110),
    .C1(_0827_),
    .X(_0828_));
 sky130_fd_sc_hd__o21ai_1 _1905_ (.A1(net113),
    .A2(_0824_),
    .B1(net121),
    .Y(_0829_));
 sky130_fd_sc_hd__a31o_1 _1906_ (.A1(net113),
    .A2(_0826_),
    .A3(_0828_),
    .B1(_0829_),
    .X(_0830_));
 sky130_fd_sc_hd__mux4_1 _1907_ (.A0(\RAM[48][1] ),
    .A1(\RAM[49][1] ),
    .A2(\RAM[50][1] ),
    .A3(\RAM[51][1] ),
    .S0(net137),
    .S1(net129),
    .X(_0831_));
 sky130_fd_sc_hd__nor2_1 _1908_ (.A(net123),
    .B(_0831_),
    .Y(_0832_));
 sky130_fd_sc_hd__mux2_1 _1909_ (.A0(\RAM[54][1] ),
    .A1(\RAM[55][1] ),
    .S(net137),
    .X(_0833_));
 sky130_fd_sc_hd__nand2_1 _1910_ (.A(net129),
    .B(_0833_),
    .Y(_0834_));
 sky130_fd_sc_hd__mux2_1 _1911_ (.A0(\RAM[52][1] ),
    .A1(\RAM[53][1] ),
    .S(net137),
    .X(_0835_));
 sky130_fd_sc_hd__nand2_1 _1912_ (.A(net110),
    .B(_0835_),
    .Y(_0836_));
 sky130_fd_sc_hd__a311o_1 _1913_ (.A1(net123),
    .A2(_0834_),
    .A3(_0836_),
    .B1(net119),
    .C1(_0832_),
    .X(_0837_));
 sky130_fd_sc_hd__o21ai_1 _1914_ (.A1(_0557_),
    .A2(_0823_),
    .B1(_0558_),
    .Y(_0838_));
 sky130_fd_sc_hd__a31o_1 _1915_ (.A1(_0557_),
    .A2(_0811_),
    .A3(_0818_),
    .B1(_0838_),
    .X(_0839_));
 sky130_fd_sc_hd__o21ai_1 _1916_ (.A1(net117),
    .A2(_0804_),
    .B1(net116),
    .Y(_0840_));
 sky130_fd_sc_hd__a31o_1 _1917_ (.A1(net117),
    .A2(_0830_),
    .A3(_0837_),
    .B1(_0840_),
    .X(_0841_));
 sky130_fd_sc_hd__nor2_1 _1918_ (.A(net7),
    .B(net105),
    .Y(_0842_));
 sky130_fd_sc_hd__a31o_1 _1919_ (.A1(net105),
    .A2(_0839_),
    .A3(_0841_),
    .B1(_0842_),
    .X(_0843_));
 sky130_fd_sc_hd__nand2_1 _1920_ (.A(net1),
    .B(_0688_),
    .Y(_0844_));
 sky130_fd_sc_hd__o211ai_4 _1921_ (.A1(_0688_),
    .A2(_0843_),
    .B1(_0844_),
    .C1(_0611_),
    .Y(_0845_));
 sky130_fd_sc_hd__or2_1 _1922_ (.A(net795),
    .B(_0611_),
    .X(_0846_));
 sky130_fd_sc_hd__nand2_1 _1923_ (.A(_0845_),
    .B(_0846_),
    .Y(_0847_));
 sky130_fd_sc_hd__inv_2 _1924_ (.A(_0847_),
    .Y(_0848_));
 sky130_fd_sc_hd__o22a_1 _1925_ (.A1(net983),
    .A2(net103),
    .B1(_0848_),
    .B2(_0640_),
    .X(_0849_));
 sky130_fd_sc_hd__o22ai_1 _1926_ (.A1(net1197),
    .A2(_0696_),
    .B1(_0849_),
    .B2(net102),
    .Y(_0850_));
 sky130_fd_sc_hd__nand2_1 _1927_ (.A(_0749_),
    .B(_0850_),
    .Y(_0851_));
 sky130_fd_sc_hd__o211a_1 _1928_ (.A1(net14),
    .A2(_0749_),
    .B1(_0851_),
    .C1(net149),
    .X(_0007_));
 sky130_fd_sc_hd__mux4_1 _1929_ (.A0(\RAM[44][2] ),
    .A1(\RAM[45][2] ),
    .A2(\RAM[46][2] ),
    .A3(\RAM[47][2] ),
    .S0(net133),
    .S1(net125),
    .X(_0852_));
 sky130_fd_sc_hd__mux4_2 _1930_ (.A0(\RAM[40][2] ),
    .A1(\RAM[41][2] ),
    .A2(\RAM[42][2] ),
    .A3(\RAM[43][2] ),
    .S0(net133),
    .S1(net125),
    .X(_0853_));
 sky130_fd_sc_hd__mux4_1 _1931_ (.A0(\RAM[32][2] ),
    .A1(\RAM[33][2] ),
    .A2(\RAM[34][2] ),
    .A3(\RAM[35][2] ),
    .S0(net134),
    .S1(net126),
    .X(_0854_));
 sky130_fd_sc_hd__mux4_1 _1932_ (.A0(\RAM[36][2] ),
    .A1(\RAM[37][2] ),
    .A2(\RAM[38][2] ),
    .A3(\RAM[39][2] ),
    .S0(net134),
    .S1(net126),
    .X(_0855_));
 sky130_fd_sc_hd__mux4_1 _1933_ (.A0(_0854_),
    .A1(_0855_),
    .A2(_0853_),
    .A3(_0852_),
    .S0(net123),
    .S1(net119),
    .X(_0856_));
 sky130_fd_sc_hd__mux4_1 _1934_ (.A0(\RAM[12][2] ),
    .A1(\RAM[13][2] ),
    .A2(\RAM[14][2] ),
    .A3(\RAM[15][2] ),
    .S0(net140),
    .S1(net130),
    .X(_0857_));
 sky130_fd_sc_hd__mux2_1 _1935_ (.A0(\RAM[8][2] ),
    .A1(\RAM[9][2] ),
    .S(net140),
    .X(_0858_));
 sky130_fd_sc_hd__nand2_1 _1936_ (.A(net111),
    .B(_0858_),
    .Y(_0859_));
 sky130_fd_sc_hd__mux2_1 _1937_ (.A0(\RAM[10][2] ),
    .A1(\RAM[11][2] ),
    .S(net140),
    .X(_0860_));
 sky130_fd_sc_hd__nand2_1 _1938_ (.A(net130),
    .B(_0860_),
    .Y(_0861_));
 sky130_fd_sc_hd__o21ai_1 _1939_ (.A1(net112),
    .A2(_0857_),
    .B1(net122),
    .Y(_0862_));
 sky130_fd_sc_hd__a31o_1 _1940_ (.A1(net112),
    .A2(_0859_),
    .A3(_0861_),
    .B1(_0862_),
    .X(_0863_));
 sky130_fd_sc_hd__mux4_1 _1941_ (.A0(\RAM[4][2] ),
    .A1(\RAM[5][2] ),
    .A2(\RAM[6][2] ),
    .A3(\RAM[7][2] ),
    .S0(net142),
    .S1(net131),
    .X(_0864_));
 sky130_fd_sc_hd__nor2_1 _1942_ (.A(net113),
    .B(_0864_),
    .Y(_0865_));
 sky130_fd_sc_hd__mux2_1 _1943_ (.A0(\RAM[2][2] ),
    .A1(\RAM[3][2] ),
    .S(net141),
    .X(_0866_));
 sky130_fd_sc_hd__nand2_1 _1944_ (.A(net131),
    .B(_0866_),
    .Y(_0867_));
 sky130_fd_sc_hd__mux2_1 _1945_ (.A0(\RAM[0][2] ),
    .A1(\RAM[1][2] ),
    .S(net141),
    .X(_0868_));
 sky130_fd_sc_hd__nand2_1 _1946_ (.A(net111),
    .B(_0868_),
    .Y(_0869_));
 sky130_fd_sc_hd__a311o_1 _1947_ (.A1(_0559_),
    .A2(_0867_),
    .A3(_0869_),
    .B1(net122),
    .C1(_0865_),
    .X(_0870_));
 sky130_fd_sc_hd__mux4_1 _1948_ (.A0(\RAM[24][2] ),
    .A1(\RAM[25][2] ),
    .A2(\RAM[26][2] ),
    .A3(\RAM[27][2] ),
    .S0(net136),
    .S1(net128),
    .X(_0871_));
 sky130_fd_sc_hd__mux4_1 _1949_ (.A0(\RAM[28][2] ),
    .A1(\RAM[29][2] ),
    .A2(\RAM[30][2] ),
    .A3(\RAM[31][2] ),
    .S0(net135),
    .S1(net127),
    .X(_0872_));
 sky130_fd_sc_hd__mux4_1 _1950_ (.A0(\RAM[20][2] ),
    .A1(\RAM[21][2] ),
    .A2(\RAM[22][2] ),
    .A3(\RAM[23][2] ),
    .S0(net136),
    .S1(net128),
    .X(_0873_));
 sky130_fd_sc_hd__mux4_1 _1951_ (.A0(\RAM[16][2] ),
    .A1(\RAM[17][2] ),
    .A2(\RAM[18][2] ),
    .A3(\RAM[19][2] ),
    .S0(net136),
    .S1(net128),
    .X(_0874_));
 sky130_fd_sc_hd__mux4_1 _1952_ (.A0(_0874_),
    .A1(_0873_),
    .A2(_0871_),
    .A3(_0872_),
    .S0(net124),
    .S1(net120),
    .X(_0875_));
 sky130_fd_sc_hd__mux4_1 _1953_ (.A0(net48),
    .A1(\RAM[61][2] ),
    .A2(\RAM[62][2] ),
    .A3(net42),
    .S0(net138),
    .S1(net129),
    .X(_0876_));
 sky130_fd_sc_hd__mux2_1 _1954_ (.A0(\RAM[56][2] ),
    .A1(\RAM[57][2] ),
    .S(net139),
    .X(_0877_));
 sky130_fd_sc_hd__nand2_1 _1955_ (.A(net111),
    .B(_0877_),
    .Y(_0878_));
 sky130_fd_sc_hd__nor2_1 _1956_ (.A(net57),
    .B(net138),
    .Y(_0879_));
 sky130_fd_sc_hd__a211o_1 _1957_ (.A1(net23),
    .A2(net138),
    .B1(net111),
    .C1(_0879_),
    .X(_0880_));
 sky130_fd_sc_hd__o21ai_1 _1958_ (.A1(net113),
    .A2(_0876_),
    .B1(net121),
    .Y(_0881_));
 sky130_fd_sc_hd__a31o_1 _1959_ (.A1(net113),
    .A2(_0878_),
    .A3(_0880_),
    .B1(_0881_),
    .X(_0882_));
 sky130_fd_sc_hd__mux4_1 _1960_ (.A0(\RAM[48][2] ),
    .A1(\RAM[49][2] ),
    .A2(\RAM[50][2] ),
    .A3(\RAM[51][2] ),
    .S0(net137),
    .S1(net129),
    .X(_0883_));
 sky130_fd_sc_hd__nor2_1 _1961_ (.A(net123),
    .B(_0883_),
    .Y(_0884_));
 sky130_fd_sc_hd__mux2_1 _1962_ (.A0(\RAM[54][2] ),
    .A1(\RAM[55][2] ),
    .S(net137),
    .X(_0885_));
 sky130_fd_sc_hd__nand2_1 _1963_ (.A(net129),
    .B(_0885_),
    .Y(_0886_));
 sky130_fd_sc_hd__mux2_1 _1964_ (.A0(\RAM[52][2] ),
    .A1(\RAM[53][2] ),
    .S(net137),
    .X(_0887_));
 sky130_fd_sc_hd__nand2_1 _1965_ (.A(net110),
    .B(_0887_),
    .Y(_0888_));
 sky130_fd_sc_hd__a311o_1 _1966_ (.A1(net123),
    .A2(_0886_),
    .A3(_0888_),
    .B1(net121),
    .C1(_0884_),
    .X(_0889_));
 sky130_fd_sc_hd__o21ai_1 _1967_ (.A1(_0557_),
    .A2(_0875_),
    .B1(_0558_),
    .Y(_0890_));
 sky130_fd_sc_hd__a31o_1 _1968_ (.A1(_0557_),
    .A2(_0863_),
    .A3(_0870_),
    .B1(_0890_),
    .X(_0891_));
 sky130_fd_sc_hd__o21ai_1 _1969_ (.A1(net117),
    .A2(_0856_),
    .B1(net116),
    .Y(_0892_));
 sky130_fd_sc_hd__a31o_1 _1970_ (.A1(net117),
    .A2(_0882_),
    .A3(_0889_),
    .B1(_0892_),
    .X(_0893_));
 sky130_fd_sc_hd__nand3_1 _1971_ (.A(net105),
    .B(_0891_),
    .C(_0893_),
    .Y(_0894_));
 sky130_fd_sc_hd__o211a_1 _1972_ (.A1(net8),
    .A2(net105),
    .B1(_0689_),
    .C1(_0894_),
    .X(_0895_));
 sky130_fd_sc_hd__a21o_1 _1973_ (.A1(net2),
    .A2(_0688_),
    .B1(_0612_),
    .X(_0896_));
 sky130_fd_sc_hd__o22a_4 _1974_ (.A1(net993),
    .A2(_0611_),
    .B1(_0895_),
    .B2(_0896_),
    .X(_0897_));
 sky130_fd_sc_hd__inv_2 _1975_ (.A(_0897_),
    .Y(_0898_));
 sky130_fd_sc_hd__o22a_1 _1976_ (.A1(net563),
    .A2(net103),
    .B1(_0897_),
    .B2(_0640_),
    .X(_0899_));
 sky130_fd_sc_hd__o22a_1 _1977_ (.A1(net1248),
    .A2(_0696_),
    .B1(_0899_),
    .B2(net102),
    .X(_0900_));
 sky130_fd_sc_hd__mux2_1 _1978_ (.A0(net15),
    .A1(_0900_),
    .S(_0749_),
    .X(_0901_));
 sky130_fd_sc_hd__and2_1 _1979_ (.A(net149),
    .B(_0901_),
    .X(_0008_));
 sky130_fd_sc_hd__mux4_1 _1980_ (.A0(\RAM[44][3] ),
    .A1(\RAM[45][3] ),
    .A2(\RAM[46][3] ),
    .A3(\RAM[47][3] ),
    .S0(net133),
    .S1(net125),
    .X(_0902_));
 sky130_fd_sc_hd__mux4_2 _1981_ (.A0(\RAM[40][3] ),
    .A1(\RAM[41][3] ),
    .A2(\RAM[42][3] ),
    .A3(\RAM[43][3] ),
    .S0(net133),
    .S1(net125),
    .X(_0903_));
 sky130_fd_sc_hd__mux4_1 _1982_ (.A0(\RAM[32][3] ),
    .A1(\RAM[33][3] ),
    .A2(\RAM[34][3] ),
    .A3(\RAM[35][3] ),
    .S0(net134),
    .S1(net126),
    .X(_0904_));
 sky130_fd_sc_hd__mux4_1 _1983_ (.A0(\RAM[36][3] ),
    .A1(\RAM[37][3] ),
    .A2(\RAM[38][3] ),
    .A3(\RAM[39][3] ),
    .S0(net134),
    .S1(net126),
    .X(_0905_));
 sky130_fd_sc_hd__mux4_1 _1984_ (.A0(_0904_),
    .A1(_0905_),
    .A2(_0903_),
    .A3(_0902_),
    .S0(net123),
    .S1(net119),
    .X(_0906_));
 sky130_fd_sc_hd__mux4_1 _1985_ (.A0(\RAM[12][3] ),
    .A1(\RAM[13][3] ),
    .A2(\RAM[14][3] ),
    .A3(\RAM[15][3] ),
    .S0(net143),
    .S1(net131),
    .X(_0907_));
 sky130_fd_sc_hd__mux2_1 _1986_ (.A0(\RAM[8][3] ),
    .A1(\RAM[9][3] ),
    .S(net143),
    .X(_0908_));
 sky130_fd_sc_hd__nand2_1 _1987_ (.A(net111),
    .B(_0908_),
    .Y(_0909_));
 sky130_fd_sc_hd__mux2_1 _1988_ (.A0(\RAM[10][3] ),
    .A1(\RAM[11][3] ),
    .S(net143),
    .X(_0910_));
 sky130_fd_sc_hd__nand2_1 _1989_ (.A(net130),
    .B(_0910_),
    .Y(_0911_));
 sky130_fd_sc_hd__o21ai_1 _1990_ (.A1(net112),
    .A2(_0907_),
    .B1(net122),
    .Y(_0912_));
 sky130_fd_sc_hd__a31o_1 _1991_ (.A1(net112),
    .A2(_0909_),
    .A3(_0911_),
    .B1(_0912_),
    .X(_0913_));
 sky130_fd_sc_hd__mux4_1 _1992_ (.A0(\RAM[4][3] ),
    .A1(\RAM[5][3] ),
    .A2(\RAM[6][3] ),
    .A3(\RAM[7][3] ),
    .S0(net142),
    .S1(net131),
    .X(_0914_));
 sky130_fd_sc_hd__nor2_1 _1993_ (.A(_0559_),
    .B(_0914_),
    .Y(_0915_));
 sky130_fd_sc_hd__mux2_1 _1994_ (.A0(\RAM[2][3] ),
    .A1(\RAM[3][3] ),
    .S(net142),
    .X(_0916_));
 sky130_fd_sc_hd__nand2_1 _1995_ (.A(net131),
    .B(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__mux2_1 _1996_ (.A0(\RAM[0][3] ),
    .A1(\RAM[1][3] ),
    .S(net142),
    .X(_0918_));
 sky130_fd_sc_hd__nand2_1 _1997_ (.A(net111),
    .B(_0918_),
    .Y(_0919_));
 sky130_fd_sc_hd__a311o_1 _1998_ (.A1(_0559_),
    .A2(_0917_),
    .A3(_0919_),
    .B1(net122),
    .C1(_0915_),
    .X(_0920_));
 sky130_fd_sc_hd__mux4_1 _1999_ (.A0(\RAM[24][3] ),
    .A1(\RAM[25][3] ),
    .A2(\RAM[26][3] ),
    .A3(\RAM[27][3] ),
    .S0(net135),
    .S1(net128),
    .X(_0921_));
 sky130_fd_sc_hd__mux4_1 _2000_ (.A0(\RAM[28][3] ),
    .A1(\RAM[29][3] ),
    .A2(\RAM[30][3] ),
    .A3(\RAM[31][3] ),
    .S0(net135),
    .S1(net127),
    .X(_0922_));
 sky130_fd_sc_hd__mux4_1 _2001_ (.A0(\RAM[20][3] ),
    .A1(\RAM[21][3] ),
    .A2(\RAM[22][3] ),
    .A3(\RAM[23][3] ),
    .S0(net136),
    .S1(net128),
    .X(_0923_));
 sky130_fd_sc_hd__mux4_1 _2002_ (.A0(\RAM[16][3] ),
    .A1(\RAM[17][3] ),
    .A2(\RAM[18][3] ),
    .A3(\RAM[19][3] ),
    .S0(net136),
    .S1(net128),
    .X(_0924_));
 sky130_fd_sc_hd__mux4_1 _2003_ (.A0(_0924_),
    .A1(_0923_),
    .A2(_0921_),
    .A3(_0922_),
    .S0(net124),
    .S1(net119),
    .X(_0925_));
 sky130_fd_sc_hd__mux4_1 _2004_ (.A0(net49),
    .A1(\RAM[61][3] ),
    .A2(\RAM[62][3] ),
    .A3(net43),
    .S0(net139),
    .S1(net129),
    .X(_0926_));
 sky130_fd_sc_hd__mux2_1 _2005_ (.A0(\RAM[56][3] ),
    .A1(\RAM[57][3] ),
    .S(net138),
    .X(_0927_));
 sky130_fd_sc_hd__nand2_1 _2006_ (.A(net111),
    .B(_0927_),
    .Y(_0928_));
 sky130_fd_sc_hd__nor2_1 _2007_ (.A(net58),
    .B(net141),
    .Y(_0929_));
 sky130_fd_sc_hd__a211o_1 _2008_ (.A1(net25),
    .A2(net138),
    .B1(net111),
    .C1(_0929_),
    .X(_0930_));
 sky130_fd_sc_hd__o21ai_1 _2009_ (.A1(net113),
    .A2(_0926_),
    .B1(net121),
    .Y(_0931_));
 sky130_fd_sc_hd__a31o_1 _2010_ (.A1(net113),
    .A2(_0928_),
    .A3(_0930_),
    .B1(_0931_),
    .X(_0932_));
 sky130_fd_sc_hd__mux4_1 _2011_ (.A0(\RAM[48][3] ),
    .A1(\RAM[49][3] ),
    .A2(\RAM[50][3] ),
    .A3(\RAM[51][3] ),
    .S0(net137),
    .S1(net129),
    .X(_0933_));
 sky130_fd_sc_hd__nor2_1 _2012_ (.A(net124),
    .B(_0933_),
    .Y(_0934_));
 sky130_fd_sc_hd__mux2_1 _2013_ (.A0(\RAM[54][3] ),
    .A1(\RAM[55][3] ),
    .S(net137),
    .X(_0935_));
 sky130_fd_sc_hd__nand2_1 _2014_ (.A(net129),
    .B(_0935_),
    .Y(_0936_));
 sky130_fd_sc_hd__mux2_1 _2015_ (.A0(\RAM[52][3] ),
    .A1(\RAM[53][3] ),
    .S(net137),
    .X(_0937_));
 sky130_fd_sc_hd__nand2_1 _2016_ (.A(net110),
    .B(_0937_),
    .Y(_0938_));
 sky130_fd_sc_hd__a311o_1 _2017_ (.A1(net124),
    .A2(_0936_),
    .A3(_0938_),
    .B1(net121),
    .C1(_0934_),
    .X(_0939_));
 sky130_fd_sc_hd__o21ai_1 _2018_ (.A1(_0557_),
    .A2(_0925_),
    .B1(_0558_),
    .Y(_0940_));
 sky130_fd_sc_hd__a31o_1 _2019_ (.A1(_0557_),
    .A2(_0913_),
    .A3(_0920_),
    .B1(_0940_),
    .X(_0941_));
 sky130_fd_sc_hd__o21ai_1 _2020_ (.A1(net117),
    .A2(_0906_),
    .B1(net116),
    .Y(_0942_));
 sky130_fd_sc_hd__a31o_1 _2021_ (.A1(net117),
    .A2(_0932_),
    .A3(_0939_),
    .B1(_0942_),
    .X(_0943_));
 sky130_fd_sc_hd__nand3_1 _2022_ (.A(net105),
    .B(_0941_),
    .C(_0943_),
    .Y(_0944_));
 sky130_fd_sc_hd__o211a_1 _2023_ (.A1(net9),
    .A2(net105),
    .B1(_0689_),
    .C1(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__a21o_1 _2024_ (.A1(net3),
    .A2(_0688_),
    .B1(_0612_),
    .X(_0946_));
 sky130_fd_sc_hd__o22a_4 _2025_ (.A1(net1005),
    .A2(_0611_),
    .B1(_0945_),
    .B2(_0946_),
    .X(_0947_));
 sky130_fd_sc_hd__o22a_1 _2026_ (.A1(net463),
    .A2(net103),
    .B1(_0947_),
    .B2(_0640_),
    .X(_0948_));
 sky130_fd_sc_hd__o22a_1 _2027_ (.A1(net1243),
    .A2(_0696_),
    .B1(_0948_),
    .B2(net102),
    .X(_0949_));
 sky130_fd_sc_hd__mux2_1 _2028_ (.A0(net16),
    .A1(_0949_),
    .S(_0749_),
    .X(_0950_));
 sky130_fd_sc_hd__and2_1 _2029_ (.A(net152),
    .B(_0950_),
    .X(_0009_));
 sky130_fd_sc_hd__or3_2 _2030_ (.A(_0556_),
    .B(net106),
    .C(_0748_),
    .X(_0951_));
 sky130_fd_sc_hd__inv_2 _2031_ (.A(_0951_),
    .Y(_0952_));
 sky130_fd_sc_hd__nor2_2 _2032_ (.A(_0549_),
    .B(_0595_),
    .Y(_0953_));
 sky130_fd_sc_hd__or2_2 _2033_ (.A(_0549_),
    .B(_0595_),
    .X(_0954_));
 sky130_fd_sc_hd__or4_4 _2034_ (.A(net1150),
    .B(net1184),
    .C(_0639_),
    .D(_0954_),
    .X(_0955_));
 sky130_fd_sc_hd__o22a_1 _2035_ (.A1(net697),
    .A2(net103),
    .B1(_0796_),
    .B2(_0955_),
    .X(_0956_));
 sky130_fd_sc_hd__a21oi_4 _2036_ (.A1(net103),
    .A2(_0955_),
    .B1(_0605_),
    .Y(_0957_));
 sky130_fd_sc_hd__o22a_1 _2037_ (.A1(net102),
    .A2(_0956_),
    .B1(_0957_),
    .B2(net134),
    .X(_0958_));
 sky130_fd_sc_hd__or2_1 _2038_ (.A(net13),
    .B(_0951_),
    .X(_0959_));
 sky130_fd_sc_hd__o211a_1 _2039_ (.A1(_0952_),
    .A2(_0958_),
    .B1(_0959_),
    .C1(net151),
    .X(_0000_));
 sky130_fd_sc_hd__o22a_1 _2040_ (.A1(net667),
    .A2(net103),
    .B1(_0848_),
    .B2(_0955_),
    .X(_0960_));
 sky130_fd_sc_hd__o22a_1 _2041_ (.A1(net126),
    .A2(_0957_),
    .B1(_0960_),
    .B2(net102),
    .X(_0961_));
 sky130_fd_sc_hd__or4_1 _2042_ (.A(_0556_),
    .B(net14),
    .C(net106),
    .D(_0748_),
    .X(_0962_));
 sky130_fd_sc_hd__o211a_1 _2043_ (.A1(_0952_),
    .A2(_0961_),
    .B1(_0962_),
    .C1(net149),
    .X(_0001_));
 sky130_fd_sc_hd__o22a_1 _2044_ (.A1(net767),
    .A2(net103),
    .B1(_0897_),
    .B2(_0955_),
    .X(_0963_));
 sky130_fd_sc_hd__o22a_1 _2045_ (.A1(net123),
    .A2(_0957_),
    .B1(_0963_),
    .B2(_0605_),
    .X(_0964_));
 sky130_fd_sc_hd__or2_1 _2046_ (.A(net15),
    .B(_0951_),
    .X(_0965_));
 sky130_fd_sc_hd__o211a_1 _2047_ (.A1(_0952_),
    .A2(_0964_),
    .B1(_0965_),
    .C1(net151),
    .X(_0002_));
 sky130_fd_sc_hd__o22a_1 _2048_ (.A1(net613),
    .A2(net103),
    .B1(_0947_),
    .B2(_0955_),
    .X(_0966_));
 sky130_fd_sc_hd__o22a_1 _2049_ (.A1(net119),
    .A2(_0957_),
    .B1(_0966_),
    .B2(_0605_),
    .X(_0967_));
 sky130_fd_sc_hd__or2_1 _2050_ (.A(net16),
    .B(_0951_),
    .X(_0968_));
 sky130_fd_sc_hd__o211a_1 _2051_ (.A1(_0952_),
    .A2(_0967_),
    .B1(_0968_),
    .C1(net151),
    .X(_0003_));
 sky130_fd_sc_hd__nor2_4 _2052_ (.A(net107),
    .B(_0571_),
    .Y(_0969_));
 sky130_fd_sc_hd__nand2_2 _2053_ (.A(net108),
    .B(_0570_),
    .Y(_0970_));
 sky130_fd_sc_hd__nand2_2 _2054_ (.A(net1034),
    .B(_0969_),
    .Y(_0971_));
 sky130_fd_sc_hd__nor2_1 _2055_ (.A(_0747_),
    .B(_0971_),
    .Y(_0972_));
 sky130_fd_sc_hd__or2_1 _2056_ (.A(net1223),
    .B(_0972_),
    .X(_0973_));
 sky130_fd_sc_hd__o311a_1 _2057_ (.A1(net13),
    .A2(_0747_),
    .A3(_0971_),
    .B1(_0973_),
    .C1(net149),
    .X(_0012_));
 sky130_fd_sc_hd__or2_1 _2058_ (.A(net1226),
    .B(_0972_),
    .X(_0974_));
 sky130_fd_sc_hd__o311a_1 _2059_ (.A1(net14),
    .A2(_0747_),
    .A3(_0971_),
    .B1(_0974_),
    .C1(net149),
    .X(_0013_));
 sky130_fd_sc_hd__or2_1 _2060_ (.A(net1160),
    .B(_0972_),
    .X(_0975_));
 sky130_fd_sc_hd__o311a_1 _2061_ (.A1(net15),
    .A2(_0747_),
    .A3(_0971_),
    .B1(net1161),
    .C1(net149),
    .X(_0014_));
 sky130_fd_sc_hd__or2_1 _2062_ (.A(net1150),
    .B(_0972_),
    .X(_0976_));
 sky130_fd_sc_hd__o311a_1 _2063_ (.A1(net16),
    .A2(_0747_),
    .A3(_0971_),
    .B1(net1151),
    .C1(net149),
    .X(_0015_));
 sky130_fd_sc_hd__nor3_1 _2064_ (.A(_0556_),
    .B(net106),
    .C(_0636_),
    .Y(_0977_));
 sky130_fd_sc_hd__o22a_1 _2065_ (.A1(net595),
    .A2(net103),
    .B1(_0955_),
    .B2(_0692_),
    .X(_0978_));
 sky130_fd_sc_hd__o22a_1 _2066_ (.A1(net118),
    .A2(_0957_),
    .B1(_0978_),
    .B2(_0605_),
    .X(_0979_));
 sky130_fd_sc_hd__mux2_1 _2067_ (.A0(_0979_),
    .A1(net13),
    .S(_0977_),
    .X(_0980_));
 sky130_fd_sc_hd__and2_1 _2068_ (.A(net151),
    .B(_0980_),
    .X(_0004_));
 sky130_fd_sc_hd__o22a_1 _2069_ (.A1(net651),
    .A2(net103),
    .B1(_0742_),
    .B2(_0955_),
    .X(_0981_));
 sky130_fd_sc_hd__o22a_1 _2070_ (.A1(net116),
    .A2(_0957_),
    .B1(_0981_),
    .B2(net102),
    .X(_0982_));
 sky130_fd_sc_hd__or4_1 _2071_ (.A(_0556_),
    .B(net14),
    .C(net106),
    .D(_0636_),
    .X(_0983_));
 sky130_fd_sc_hd__o211a_1 _2072_ (.A1(_0977_),
    .A2(_0982_),
    .B1(_0983_),
    .C1(net151),
    .X(_0005_));
 sky130_fd_sc_hd__nor2_1 _2073_ (.A(_0634_),
    .B(_0971_),
    .Y(_0984_));
 sky130_fd_sc_hd__or3_1 _2074_ (.A(net13),
    .B(_0634_),
    .C(_0971_),
    .X(_0985_));
 sky130_fd_sc_hd__o211a_1 _2075_ (.A1(net1184),
    .A2(_0984_),
    .B1(_0985_),
    .C1(net151),
    .X(_0016_));
 sky130_fd_sc_hd__or3_1 _2076_ (.A(net14),
    .B(_0634_),
    .C(_0971_),
    .X(_0986_));
 sky130_fd_sc_hd__o211a_1 _2077_ (.A1(net1080),
    .A2(_0984_),
    .B1(_0986_),
    .C1(net151),
    .X(_0017_));
 sky130_fd_sc_hd__nor2_1 _2078_ (.A(_0578_),
    .B(_0595_),
    .Y(_0987_));
 sky130_fd_sc_hd__and2_1 _2079_ (.A(_0550_),
    .B(_0987_),
    .X(_0988_));
 sky130_fd_sc_hd__and3_4 _2080_ (.A(net1110),
    .B(_0606_),
    .C(_0988_),
    .X(_0989_));
 sky130_fd_sc_hd__or2_2 _2081_ (.A(\insin[2] ),
    .B(_0592_),
    .X(_0990_));
 sky130_fd_sc_hd__or4_1 _2082_ (.A(\insin[4] ),
    .B(net148),
    .C(_0639_),
    .D(_0990_),
    .X(_0991_));
 sky130_fd_sc_hd__nor3_1 _2083_ (.A(net1150),
    .B(_0605_),
    .C(_0991_),
    .Y(_0992_));
 sky130_fd_sc_hd__nor2_4 _2084_ (.A(_0989_),
    .B(net101),
    .Y(_0993_));
 sky130_fd_sc_hd__or4_4 _2085_ (.A(net123),
    .B(net137),
    .C(net110),
    .D(net96),
    .X(_0994_));
 sky130_fd_sc_hd__nor3_4 _2086_ (.A(net121),
    .B(_0641_),
    .C(net96),
    .Y(_0995_));
 sky130_fd_sc_hd__or3_4 _2087_ (.A(net121),
    .B(_0641_),
    .C(net96),
    .X(_0996_));
 sky130_fd_sc_hd__nor2_2 _2088_ (.A(_0994_),
    .B(_0996_),
    .Y(_0997_));
 sky130_fd_sc_hd__a22o_4 _2089_ (.A1(net1086),
    .A2(_0989_),
    .B1(net100),
    .B2(net1156),
    .X(_0998_));
 sky130_fd_sc_hd__mux2_1 _2090_ (.A0(net569),
    .A1(net93),
    .S(_0997_),
    .X(_0024_));
 sky130_fd_sc_hd__a22o_4 _2091_ (.A1(net1096),
    .A2(_0989_),
    .B1(net100),
    .B2(net1121),
    .X(_0999_));
 sky130_fd_sc_hd__mux2_1 _2092_ (.A0(net343),
    .A1(_0999_),
    .S(_0997_),
    .X(_0025_));
 sky130_fd_sc_hd__a22o_2 _2093_ (.A1(net1101),
    .A2(_0989_),
    .B1(net100),
    .B2(net1028),
    .X(_1000_));
 sky130_fd_sc_hd__mux2_1 _2094_ (.A0(net269),
    .A1(net87),
    .S(_0997_),
    .X(_0026_));
 sky130_fd_sc_hd__a22o_4 _2095_ (.A1(net1071),
    .A2(_0989_),
    .B1(net100),
    .B2(net1128),
    .X(_1001_));
 sky130_fd_sc_hd__mux2_1 _2096_ (.A0(net263),
    .A1(net82),
    .S(_0997_),
    .X(_0027_));
 sky130_fd_sc_hd__a22o_2 _2097_ (.A1(net1082),
    .A2(_0989_),
    .B1(net100),
    .B2(net1030),
    .X(_1002_));
 sky130_fd_sc_hd__mux2_1 _2098_ (.A0(net489),
    .A1(net75),
    .S(_0997_),
    .X(_0028_));
 sky130_fd_sc_hd__a22o_4 _2099_ (.A1(net1112),
    .A2(_0989_),
    .B1(net100),
    .B2(net1103),
    .X(_1003_));
 sky130_fd_sc_hd__mux2_1 _2100_ (.A0(net203),
    .A1(net74),
    .S(_0997_),
    .X(_0029_));
 sky130_fd_sc_hd__nor2_1 _2101_ (.A(net130),
    .B(net96),
    .Y(_1004_));
 sky130_fd_sc_hd__and3_4 _2102_ (.A(\MAR[2] ),
    .B(net141),
    .C(_1004_),
    .X(_1005_));
 sky130_fd_sc_hd__o2111a_4 _2103_ (.A1(_0989_),
    .A2(net101),
    .B1(_0557_),
    .C1(net116),
    .D1(net119),
    .X(_1006_));
 sky130_fd_sc_hd__inv_2 _2104_ (.A(_1006_),
    .Y(_1007_));
 sky130_fd_sc_hd__nand2_4 _2105_ (.A(_1005_),
    .B(_1006_),
    .Y(_1008_));
 sky130_fd_sc_hd__mux2_1 _2106_ (.A0(net93),
    .A1(net579),
    .S(_1008_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _2107_ (.A0(net88),
    .A1(net537),
    .S(_1008_),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _2108_ (.A0(net83),
    .A1(net903),
    .S(_1008_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _2109_ (.A0(net80),
    .A1(net367),
    .S(_1008_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _2110_ (.A0(net75),
    .A1(net941),
    .S(_1008_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _2111_ (.A0(net71),
    .A1(net787),
    .S(_1008_),
    .X(_0035_));
 sky130_fd_sc_hd__o2111a_4 _2112_ (.A1(_0989_),
    .A2(net101),
    .B1(net113),
    .C1(net137),
    .D1(net129),
    .X(_1009_));
 sky130_fd_sc_hd__nand2_4 _2113_ (.A(_0995_),
    .B(_1009_),
    .Y(_1010_));
 sky130_fd_sc_hd__mux2_1 _2114_ (.A0(net94),
    .A1(net851),
    .S(_1010_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _2115_ (.A0(net90),
    .A1(net543),
    .S(_1010_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _2116_ (.A0(net87),
    .A1(net863),
    .S(_1010_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _2117_ (.A0(net82),
    .A1(net883),
    .S(_1010_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _2118_ (.A0(net78),
    .A1(net557),
    .S(_1010_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _2119_ (.A0(net74),
    .A1(net645),
    .S(_1010_),
    .X(_0041_));
 sky130_fd_sc_hd__and3_1 _2120_ (.A(\last_addr[2] ),
    .B(\last_addr[1] ),
    .C(\last_addr[0] ),
    .X(_1011_));
 sky130_fd_sc_hd__and2_1 _2121_ (.A(\last_addr[3] ),
    .B(_1011_),
    .X(_1012_));
 sky130_fd_sc_hd__and3_1 _2122_ (.A(\last_addr[5] ),
    .B(\last_addr[4] ),
    .C(_1012_),
    .X(_1013_));
 sky130_fd_sc_hd__and2_1 _2123_ (.A(\last_addr[6] ),
    .B(_1013_),
    .X(_1014_));
 sky130_fd_sc_hd__and3_1 _2124_ (.A(net1063),
    .B(\last_addr[7] ),
    .C(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__and2_1 _2125_ (.A(net1044),
    .B(_1015_),
    .X(_1016_));
 sky130_fd_sc_hd__nor2_1 _2126_ (.A(\last_addr[10] ),
    .B(_1016_),
    .Y(_1017_));
 sky130_fd_sc_hd__nand2_1 _2127_ (.A(\last_addr[10] ),
    .B(_1016_),
    .Y(_1018_));
 sky130_fd_sc_hd__nor2_1 _2128_ (.A(\last_addr[11] ),
    .B(\ROM_addr_buff[11] ),
    .Y(_1019_));
 sky130_fd_sc_hd__and2_1 _2129_ (.A(\last_addr[11] ),
    .B(\ROM_addr_buff[11] ),
    .X(_1020_));
 sky130_fd_sc_hd__o221a_1 _2130_ (.A1(\ROM_addr_buff[10] ),
    .A2(_1017_),
    .B1(_1019_),
    .B2(_1020_),
    .C1(_1018_),
    .X(_1021_));
 sky130_fd_sc_hd__a21bo_1 _2131_ (.A1(net1016),
    .A2(_1017_),
    .B1_N(_1021_),
    .X(_1022_));
 sky130_fd_sc_hd__or4b_1 _2132_ (.A(\last_addr[11] ),
    .B(\ROM_addr_buff[10] ),
    .C(_1018_),
    .D_N(\ROM_addr_buff[11] ),
    .X(_1023_));
 sky130_fd_sc_hd__nor2_1 _2133_ (.A(net1044),
    .B(_1015_),
    .Y(_1024_));
 sky130_fd_sc_hd__o21ai_1 _2134_ (.A1(_1016_),
    .A2(_1024_),
    .B1(\ROM_addr_buff[9] ),
    .Y(_1025_));
 sky130_fd_sc_hd__or3_1 _2135_ (.A(\ROM_addr_buff[9] ),
    .B(_1016_),
    .C(_1024_),
    .X(_1026_));
 sky130_fd_sc_hd__a21oi_1 _2136_ (.A1(\last_addr[7] ),
    .A2(_1014_),
    .B1(\last_addr[8] ),
    .Y(_1027_));
 sky130_fd_sc_hd__or2_1 _2137_ (.A(_1015_),
    .B(_1027_),
    .X(_1028_));
 sky130_fd_sc_hd__xnor2_1 _2138_ (.A(\ROM_addr_buff[8] ),
    .B(_1028_),
    .Y(_1029_));
 sky130_fd_sc_hd__xnor2_1 _2139_ (.A(\last_addr[7] ),
    .B(_1014_),
    .Y(_1030_));
 sky130_fd_sc_hd__a21oi_1 _2140_ (.A1(\last_addr[4] ),
    .A2(_1012_),
    .B1(\last_addr[5] ),
    .Y(_1031_));
 sky130_fd_sc_hd__or2_1 _2141_ (.A(_1013_),
    .B(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__xnor2_1 _2142_ (.A(\ROM_addr_buff[5] ),
    .B(_1032_),
    .Y(_1033_));
 sky130_fd_sc_hd__xnor2_1 _2143_ (.A(\last_addr[4] ),
    .B(_1012_),
    .Y(_1034_));
 sky130_fd_sc_hd__xnor2_1 _2144_ (.A(\ROM_addr_buff[4] ),
    .B(_1034_),
    .Y(_1035_));
 sky130_fd_sc_hd__nor2_1 _2145_ (.A(\last_addr[3] ),
    .B(_1011_),
    .Y(_1036_));
 sky130_fd_sc_hd__or2_1 _2146_ (.A(_1012_),
    .B(_1036_),
    .X(_1037_));
 sky130_fd_sc_hd__xnor2_1 _2147_ (.A(\ROM_addr_buff[3] ),
    .B(_1037_),
    .Y(_1038_));
 sky130_fd_sc_hd__a21oi_1 _2148_ (.A1(\last_addr[1] ),
    .A2(\last_addr[0] ),
    .B1(\last_addr[2] ),
    .Y(_1039_));
 sky130_fd_sc_hd__nor3_1 _2149_ (.A(\ROM_addr_buff[2] ),
    .B(_1011_),
    .C(_1039_),
    .Y(_1040_));
 sky130_fd_sc_hd__o21a_1 _2150_ (.A1(_1011_),
    .A2(_1039_),
    .B1(\ROM_addr_buff[2] ),
    .X(_1041_));
 sky130_fd_sc_hd__xnor2_1 _2151_ (.A(\last_addr[1] ),
    .B(\ROM_addr_buff[1] ),
    .Y(_1042_));
 sky130_fd_sc_hd__mux2_1 _2152_ (.A0(\last_addr[0] ),
    .A1(\ROM_addr_buff[0] ),
    .S(_1042_),
    .X(_1043_));
 sky130_fd_sc_hd__nor3_2 _2153_ (.A(net1188),
    .B(_0553_),
    .C(_0572_),
    .Y(_1044_));
 sky130_fd_sc_hd__nor2_1 _2154_ (.A(\last_addr[6] ),
    .B(_1013_),
    .Y(_1045_));
 sky130_fd_sc_hd__or2_1 _2155_ (.A(_1014_),
    .B(_1045_),
    .X(_1046_));
 sky130_fd_sc_hd__xnor2_1 _2156_ (.A(\ROM_addr_buff[6] ),
    .B(_1046_),
    .Y(_1047_));
 sky130_fd_sc_hd__a21oi_1 _2157_ (.A1(\mem_cycle[1] ),
    .A2(_0746_),
    .B1(net1182),
    .Y(_1048_));
 sky130_fd_sc_hd__nand2_2 _2158_ (.A(_0570_),
    .B(_0574_),
    .Y(_1049_));
 sky130_fd_sc_hd__and4b_1 _2159_ (.A_N(_0613_),
    .B(_0585_),
    .C(net145),
    .D(_0588_),
    .X(_1050_));
 sky130_fd_sc_hd__o31a_1 _2160_ (.A1(net1170),
    .A2(_0574_),
    .A3(_1050_),
    .B1(_0969_),
    .X(_1051_));
 sky130_fd_sc_hd__xnor2_1 _2161_ (.A(net1074),
    .B(_1030_),
    .Y(_1052_));
 sky130_fd_sc_hd__a2111o_1 _2162_ (.A1(\last_addr[0] ),
    .A2(\ROM_addr_buff[0] ),
    .B1(_1038_),
    .C1(_1040_),
    .D1(_1041_),
    .X(_1053_));
 sky130_fd_sc_hd__or4b_1 _2163_ (.A(_1033_),
    .B(_1035_),
    .C(_1053_),
    .D_N(_1043_),
    .X(_1054_));
 sky130_fd_sc_hd__or4_1 _2164_ (.A(_1029_),
    .B(_1047_),
    .C(_1052_),
    .D(_1054_),
    .X(_1055_));
 sky130_fd_sc_hd__a21bo_1 _2165_ (.A1(_1022_),
    .A2(_1023_),
    .B1_N(_1044_),
    .X(_1056_));
 sky130_fd_sc_hd__and4bb_2 _2166_ (.A_N(_1055_),
    .B_N(_1056_),
    .C(_1025_),
    .D(_1026_),
    .X(_1057_));
 sky130_fd_sc_hd__or3_1 _2167_ (.A(net106),
    .B(_1048_),
    .C(_1049_),
    .X(_1058_));
 sky130_fd_sc_hd__o221a_1 _2168_ (.A1(net1182),
    .A2(_1051_),
    .B1(_1057_),
    .B2(_1058_),
    .C1(net154),
    .X(_0042_));
 sky130_fd_sc_hd__nor2_1 _2169_ (.A(_0553_),
    .B(_0970_),
    .Y(_1059_));
 sky130_fd_sc_hd__o21ai_1 _2170_ (.A1(net1182),
    .A2(_0746_),
    .B1(net1188),
    .Y(_1060_));
 sky130_fd_sc_hd__o221a_1 _2171_ (.A1(net1188),
    .A2(_1059_),
    .B1(net1189),
    .B2(_0970_),
    .C1(net154),
    .X(_0043_));
 sky130_fd_sc_hd__o21a_1 _2172_ (.A1(_0633_),
    .A2(_0970_),
    .B1(_0554_),
    .X(_1061_));
 sky130_fd_sc_hd__a31oi_2 _2173_ (.A1(net1188),
    .A2(_0553_),
    .A3(_0746_),
    .B1(_1044_),
    .Y(_1062_));
 sky130_fd_sc_hd__o21ai_1 _2174_ (.A1(_0554_),
    .A2(_0633_),
    .B1(_1062_),
    .Y(_1063_));
 sky130_fd_sc_hd__a211oi_1 _2175_ (.A1(_0969_),
    .A2(_1063_),
    .B1(net1206),
    .C1(net147),
    .Y(_0044_));
 sky130_fd_sc_hd__and4_1 _2176_ (.A(\mem_cycle[1] ),
    .B(\mem_cycle[0] ),
    .C(net1178),
    .D(\mem_cycle[2] ),
    .X(_1064_));
 sky130_fd_sc_hd__inv_2 _2177_ (.A(_1064_),
    .Y(_1065_));
 sky130_fd_sc_hd__a31o_1 _2178_ (.A1(\mem_cycle[1] ),
    .A2(\mem_cycle[0] ),
    .A3(\mem_cycle[2] ),
    .B1(net1178),
    .X(_1066_));
 sky130_fd_sc_hd__a31o_1 _2179_ (.A1(_1062_),
    .A2(_1065_),
    .A3(_1066_),
    .B1(_0970_),
    .X(_1067_));
 sky130_fd_sc_hd__o221a_1 _2180_ (.A1(net1178),
    .A2(_0969_),
    .B1(_1057_),
    .B2(_1067_),
    .C1(net154),
    .X(_0045_));
 sky130_fd_sc_hd__nand2_1 _2181_ (.A(net1168),
    .B(_1064_),
    .Y(_1068_));
 sky130_fd_sc_hd__or2_1 _2182_ (.A(net1168),
    .B(_1064_),
    .X(_1069_));
 sky130_fd_sc_hd__a31o_1 _2183_ (.A1(_1062_),
    .A2(_1068_),
    .A3(_1069_),
    .B1(_0970_),
    .X(_1070_));
 sky130_fd_sc_hd__o221a_1 _2184_ (.A1(net1168),
    .A2(_0969_),
    .B1(_1057_),
    .B2(_1070_),
    .C1(net154),
    .X(_0046_));
 sky130_fd_sc_hd__or4_4 _2185_ (.A(_0559_),
    .B(net141),
    .C(net131),
    .D(net96),
    .X(_1071_));
 sky130_fd_sc_hd__nor2_2 _2186_ (.A(_0996_),
    .B(_1071_),
    .Y(_1072_));
 sky130_fd_sc_hd__mux2_1 _2187_ (.A0(net323),
    .A1(net94),
    .S(_1072_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _2188_ (.A0(net201),
    .A1(net90),
    .S(_1072_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _2189_ (.A0(net353),
    .A1(net86),
    .S(_1072_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _2190_ (.A0(net419),
    .A1(net82),
    .S(_1072_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _2191_ (.A0(net385),
    .A1(net78),
    .S(_1072_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _2192_ (.A0(net181),
    .A1(net74),
    .S(_1072_),
    .X(_0052_));
 sky130_fd_sc_hd__nor2_1 _2193_ (.A(net116),
    .B(net96),
    .Y(_1073_));
 sky130_fd_sc_hd__and3b_4 _2194_ (.A_N(net120),
    .B(_1073_),
    .C(net117),
    .X(_1074_));
 sky130_fd_sc_hd__or4_4 _2195_ (.A(_0557_),
    .B(net116),
    .C(net120),
    .D(net96),
    .X(_1075_));
 sky130_fd_sc_hd__nand2_4 _2196_ (.A(_1009_),
    .B(_1074_),
    .Y(_1076_));
 sky130_fd_sc_hd__mux2_1 _2197_ (.A0(_0998_),
    .A1(net779),
    .S(_1076_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _2198_ (.A0(net89),
    .A1(net917),
    .S(_1076_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _2199_ (.A0(net84),
    .A1(net639),
    .S(_1076_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _2200_ (.A0(net79),
    .A1(net717),
    .S(_1076_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _2201_ (.A0(net76),
    .A1(net713),
    .S(_1076_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _2202_ (.A0(net71),
    .A1(net673),
    .S(_1076_),
    .X(_0058_));
 sky130_fd_sc_hd__nand2_4 _2203_ (.A(_0995_),
    .B(_1005_),
    .Y(_1077_));
 sky130_fd_sc_hd__mux2_1 _2204_ (.A0(net94),
    .A1(net965),
    .S(_1077_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _2205_ (.A0(net90),
    .A1(net875),
    .S(_1077_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _2206_ (.A0(net86),
    .A1(net943),
    .S(_1077_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _2207_ (.A0(net82),
    .A1(net927),
    .S(_1077_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _2208_ (.A0(net78),
    .A1(net635),
    .S(_1077_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _2209_ (.A0(net74),
    .A1(net953),
    .S(_1077_),
    .X(_0064_));
 sky130_fd_sc_hd__and3_4 _2210_ (.A(net117),
    .B(net120),
    .C(_1073_),
    .X(_1078_));
 sky130_fd_sc_hd__inv_2 _2211_ (.A(_1078_),
    .Y(_1079_));
 sky130_fd_sc_hd__nand2_4 _2212_ (.A(_1005_),
    .B(_1078_),
    .Y(_1080_));
 sky130_fd_sc_hd__mux2_1 _2213_ (.A0(net92),
    .A1(net637),
    .S(_1080_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _2214_ (.A0(net89),
    .A1(net731),
    .S(_1080_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _2215_ (.A0(net83),
    .A1(net435),
    .S(_1080_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _2216_ (.A0(net79),
    .A1(net835),
    .S(_1080_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _2217_ (.A0(net76),
    .A1(net733),
    .S(_1080_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _2218_ (.A0(net71),
    .A1(net745),
    .S(_1080_),
    .X(_0070_));
 sky130_fd_sc_hd__and4bb_4 _2219_ (.A_N(net135),
    .B_N(net96),
    .C(net127),
    .D(\MAR[2] ),
    .X(_1081_));
 sky130_fd_sc_hd__nand2_2 _2220_ (.A(_0995_),
    .B(_1081_),
    .Y(_1082_));
 sky130_fd_sc_hd__mux2_1 _2221_ (.A0(net94),
    .A1(net373),
    .S(_1082_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _2222_ (.A0(net90),
    .A1(net457),
    .S(_1082_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _2223_ (.A0(net86),
    .A1(net339),
    .S(_1082_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _2224_ (.A0(net82),
    .A1(net581),
    .S(_1082_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _2225_ (.A0(net78),
    .A1(net355),
    .S(_1082_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _2226_ (.A0(net74),
    .A1(net497),
    .S(_1082_),
    .X(_0076_));
 sky130_fd_sc_hd__nor4_2 _2227_ (.A(net117),
    .B(_0558_),
    .C(net119),
    .D(net96),
    .Y(_1083_));
 sky130_fd_sc_hd__or4_4 _2228_ (.A(net117),
    .B(_0558_),
    .C(net119),
    .D(net96),
    .X(_1084_));
 sky130_fd_sc_hd__a31o_4 _2229_ (.A1(net124),
    .A2(net139),
    .A3(net129),
    .B1(net96),
    .X(_1085_));
 sky130_fd_sc_hd__nand2_4 _2230_ (.A(net1265),
    .B(_1085_),
    .Y(_1086_));
 sky130_fd_sc_hd__mux2_1 _2231_ (.A0(net93),
    .A1(net695),
    .S(_1086_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _2232_ (.A0(net88),
    .A1(net555),
    .S(_1086_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _2233_ (.A0(net85),
    .A1(net677),
    .S(_1086_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _2234_ (.A0(net80),
    .A1(net691),
    .S(_1086_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _2235_ (.A0(net75),
    .A1(net517),
    .S(_1086_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _2236_ (.A0(net72),
    .A1(net867),
    .S(_1086_),
    .X(_0082_));
 sky130_fd_sc_hd__nand2_2 _2237_ (.A(_0995_),
    .B(_1085_),
    .Y(_1087_));
 sky130_fd_sc_hd__mux2_1 _2238_ (.A0(net94),
    .A1(net769),
    .S(_1087_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _2239_ (.A0(net90),
    .A1(net729),
    .S(_1087_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _2240_ (.A0(net86),
    .A1(net721),
    .S(_1087_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _2241_ (.A0(net82),
    .A1(net949),
    .S(_1087_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _2242_ (.A0(net78),
    .A1(net877),
    .S(_1087_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _2243_ (.A0(net74),
    .A1(net737),
    .S(_1087_),
    .X(_0088_));
 sky130_fd_sc_hd__and3_2 _2244_ (.A(net113),
    .B(net141),
    .C(_1004_),
    .X(_1088_));
 sky130_fd_sc_hd__or4b_4 _2245_ (.A(net124),
    .B(net130),
    .C(_0993_),
    .D_N(net140),
    .X(_1089_));
 sky130_fd_sc_hd__nor2_4 _2246_ (.A(_0996_),
    .B(_1089_),
    .Y(_1090_));
 sky130_fd_sc_hd__mux2_1 _2247_ (.A0(net441),
    .A1(net94),
    .S(_1090_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _2248_ (.A0(net253),
    .A1(net90),
    .S(_1090_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _2249_ (.A0(net223),
    .A1(net87),
    .S(_1090_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _2250_ (.A0(net199),
    .A1(net82),
    .S(_1090_),
    .X(_0092_));
 sky130_fd_sc_hd__mux2_1 _2251_ (.A0(net179),
    .A1(net78),
    .S(_1090_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _2252_ (.A0(net243),
    .A1(net74),
    .S(_1090_),
    .X(_0094_));
 sky130_fd_sc_hd__nor2_4 _2253_ (.A(_1071_),
    .B(_1075_),
    .Y(_1091_));
 sky130_fd_sc_hd__mux2_1 _2254_ (.A0(net363),
    .A1(_0998_),
    .S(_1091_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _2255_ (.A0(net307),
    .A1(net89),
    .S(_1091_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _2256_ (.A0(net591),
    .A1(net83),
    .S(_1091_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _2257_ (.A0(net313),
    .A1(net79),
    .S(_1091_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _2258_ (.A0(net325),
    .A1(net76),
    .S(_1091_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _2259_ (.A0(net845),
    .A1(net71),
    .S(_1091_),
    .X(_0100_));
 sky130_fd_sc_hd__nand2_4 _2260_ (.A(_1006_),
    .B(_1009_),
    .Y(_1092_));
 sky130_fd_sc_hd__mux2_1 _2261_ (.A0(net93),
    .A1(net933),
    .S(_1092_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _2262_ (.A0(net88),
    .A1(net857),
    .S(_1092_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _2263_ (.A0(net85),
    .A1(net509),
    .S(_1092_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _2264_ (.A0(net80),
    .A1(net823),
    .S(_1092_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _2265_ (.A0(net75),
    .A1(net657),
    .S(_1092_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _2266_ (.A0(net72),
    .A1(net583),
    .S(_1092_),
    .X(_0106_));
 sky130_fd_sc_hd__a21oi_2 _2267_ (.A1(net156),
    .A2(_0993_),
    .B1(net105),
    .Y(_1093_));
 sky130_fd_sc_hd__or2_1 _2268_ (.A(net1227),
    .B(_1093_),
    .X(_1094_));
 sky130_fd_sc_hd__o311a_1 _2269_ (.A1(net105),
    .A2(_0993_),
    .A3(net94),
    .B1(_1094_),
    .C1(net156),
    .X(_0107_));
 sky130_fd_sc_hd__or2_1 _2270_ (.A(net1215),
    .B(_1093_),
    .X(_1095_));
 sky130_fd_sc_hd__o311a_1 _2271_ (.A1(net105),
    .A2(_0993_),
    .A3(net90),
    .B1(_1095_),
    .C1(net156),
    .X(_0108_));
 sky130_fd_sc_hd__or2_1 _2272_ (.A(net1212),
    .B(_1093_),
    .X(_1096_));
 sky130_fd_sc_hd__o311a_1 _2273_ (.A1(net105),
    .A2(_0993_),
    .A3(net87),
    .B1(_1096_),
    .C1(net156),
    .X(_0109_));
 sky130_fd_sc_hd__or2_1 _2274_ (.A(net1221),
    .B(_1093_),
    .X(_1097_));
 sky130_fd_sc_hd__o311a_1 _2275_ (.A1(_0643_),
    .A2(_0993_),
    .A3(net82),
    .B1(_1097_),
    .C1(net156),
    .X(_0110_));
 sky130_fd_sc_hd__or2_1 _2276_ (.A(net1201),
    .B(_1093_),
    .X(_1098_));
 sky130_fd_sc_hd__o311a_1 _2277_ (.A1(_0643_),
    .A2(_0993_),
    .A3(net78),
    .B1(_1098_),
    .C1(net156),
    .X(_0111_));
 sky130_fd_sc_hd__or2_1 _2278_ (.A(net1213),
    .B(_1093_),
    .X(_1099_));
 sky130_fd_sc_hd__o311a_1 _2279_ (.A1(_0643_),
    .A2(net96),
    .A3(net74),
    .B1(_1099_),
    .C1(net156),
    .X(_0112_));
 sky130_fd_sc_hd__a31o_4 _2280_ (.A1(net118),
    .A2(net116),
    .A3(net121),
    .B1(net96),
    .X(_1100_));
 sky130_fd_sc_hd__inv_2 _2281_ (.A(_1100_),
    .Y(_1101_));
 sky130_fd_sc_hd__nand2_4 _2282_ (.A(_1088_),
    .B(_1100_),
    .Y(_1102_));
 sky130_fd_sc_hd__mux2_1 _2283_ (.A0(net94),
    .A1(net615),
    .S(_1102_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _2284_ (.A0(net90),
    .A1(net529),
    .S(_1102_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _2285_ (.A0(net87),
    .A1(net681),
    .S(_1102_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _2286_ (.A0(net82),
    .A1(net837),
    .S(_1102_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _2287_ (.A0(net77),
    .A1(net755),
    .S(_1102_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _2288_ (.A0(net74),
    .A1(net811),
    .S(_1102_),
    .X(_0118_));
 sky130_fd_sc_hd__or4_4 _2289_ (.A(net124),
    .B(net136),
    .C(net128),
    .D(net96),
    .X(_1103_));
 sky130_fd_sc_hd__nor2_2 _2290_ (.A(_0996_),
    .B(_1103_),
    .Y(_1104_));
 sky130_fd_sc_hd__mux2_1 _2291_ (.A0(net309),
    .A1(net94),
    .S(_1104_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _2292_ (.A0(net233),
    .A1(net90),
    .S(_1104_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _2293_ (.A0(net229),
    .A1(net87),
    .S(_1104_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _2294_ (.A0(net251),
    .A1(net82),
    .S(_1104_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _2295_ (.A0(net267),
    .A1(net78),
    .S(_1104_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _2296_ (.A0(net219),
    .A1(net74),
    .S(_1104_),
    .X(_0124_));
 sky130_fd_sc_hd__o21a_1 _2297_ (.A1(_0571_),
    .A2(_0574_),
    .B1(net108),
    .X(_1105_));
 sky130_fd_sc_hd__inv_2 _2298_ (.A(_1105_),
    .Y(_1106_));
 sky130_fd_sc_hd__or4_1 _2299_ (.A(_0552_),
    .B(\mem_cycle[3] ),
    .C(\mem_cycle[2] ),
    .D(_0573_),
    .X(_1107_));
 sky130_fd_sc_hd__inv_2 _2300_ (.A(_1107_),
    .Y(_1108_));
 sky130_fd_sc_hd__and3_1 _2301_ (.A(_0552_),
    .B(\mem_cycle[1] ),
    .C(_0553_),
    .X(_1109_));
 sky130_fd_sc_hd__or3b_1 _2302_ (.A(_0573_),
    .B(\mem_cycle[4] ),
    .C_N(\mem_cycle[3] ),
    .X(_1110_));
 sky130_fd_sc_hd__or3b_2 _2303_ (.A(_1108_),
    .B(_1109_),
    .C_N(_1110_),
    .X(_1111_));
 sky130_fd_sc_hd__or4_1 _2304_ (.A(\startup_cycle[6] ),
    .B(\startup_cycle[5] ),
    .C(_0543_),
    .D(_0568_),
    .X(_1112_));
 sky130_fd_sc_hd__or3_1 _2305_ (.A(net1090),
    .B(net1208),
    .C(_0568_),
    .X(_1113_));
 sky130_fd_sc_hd__nand2_1 _2306_ (.A(_0542_),
    .B(net1208),
    .Y(_1114_));
 sky130_fd_sc_hd__or3_1 _2307_ (.A(_0544_),
    .B(net1123),
    .C(_0567_),
    .X(_1115_));
 sky130_fd_sc_hd__nor3_1 _2308_ (.A(net1088),
    .B(_1114_),
    .C(_1115_),
    .Y(_1116_));
 sky130_fd_sc_hd__nand2_2 _2309_ (.A(net1234),
    .B(net1123),
    .Y(_1117_));
 sky130_fd_sc_hd__or4_2 _2310_ (.A(net1088),
    .B(_0567_),
    .C(_1114_),
    .D(_1117_),
    .X(_1118_));
 sky130_fd_sc_hd__nand3b_2 _2311_ (.A_N(_1116_),
    .B(_1118_),
    .C(_1113_),
    .Y(_1119_));
 sky130_fd_sc_hd__o211ai_4 _2312_ (.A1(_1049_),
    .A2(_1111_),
    .B1(_1119_),
    .C1(_1105_),
    .Y(_1120_));
 sky130_fd_sc_hd__and3_1 _2313_ (.A(\mem_cycle[3] ),
    .B(_0554_),
    .C(_1109_),
    .X(_1121_));
 sky130_fd_sc_hd__o211a_1 _2314_ (.A1(net1036),
    .A2(net1205),
    .B1(_1109_),
    .C1(net1178),
    .X(_1122_));
 sky130_fd_sc_hd__nor2_1 _2315_ (.A(_0554_),
    .B(_1110_),
    .Y(_1123_));
 sky130_fd_sc_hd__nor2_1 _2316_ (.A(net1205),
    .B(_1110_),
    .Y(_1124_));
 sky130_fd_sc_hd__a221o_1 _2317_ (.A1(net1114),
    .A2(_1123_),
    .B1(_1124_),
    .B2(net1193),
    .C1(_1122_),
    .X(_1125_));
 sky130_fd_sc_hd__nand2b_1 _2318_ (.A_N(net1218),
    .B(_1120_),
    .Y(_1126_));
 sky130_fd_sc_hd__a211o_1 _2319_ (.A1(_0570_),
    .A2(_1125_),
    .B1(_1120_),
    .C1(_1116_),
    .X(_1127_));
 sky130_fd_sc_hd__and3_1 _2320_ (.A(net154),
    .B(net1219),
    .C(_1127_),
    .X(_0125_));
 sky130_fd_sc_hd__a22o_1 _2321_ (.A1(\ROM_addr_buff[6] ),
    .A2(_1121_),
    .B1(_1124_),
    .B2(net1016),
    .X(_1128_));
 sky130_fd_sc_hd__a211o_1 _2322_ (.A1(\ROM_addr_buff[2] ),
    .A2(_1123_),
    .B1(_1128_),
    .C1(_1108_),
    .X(_1129_));
 sky130_fd_sc_hd__nand2_1 _2323_ (.A(_0570_),
    .B(_1129_),
    .Y(_1130_));
 sky130_fd_sc_hd__a21oi_1 _2324_ (.A1(_1118_),
    .A2(_1130_),
    .B1(_1120_),
    .Y(_1131_));
 sky130_fd_sc_hd__a211o_1 _2325_ (.A1(net1018),
    .A2(_1120_),
    .B1(_1131_),
    .C1(net147),
    .X(_0126_));
 sky130_fd_sc_hd__o211a_1 _2326_ (.A1(\ROM_addr_buff[7] ),
    .A2(\mem_cycle[2] ),
    .B1(_1109_),
    .C1(\mem_cycle[3] ),
    .X(_1132_));
 sky130_fd_sc_hd__a22o_1 _2327_ (.A1(\ROM_addr_buff[3] ),
    .A2(_1123_),
    .B1(_1124_),
    .B2(\ROM_addr_buff[11] ),
    .X(_1133_));
 sky130_fd_sc_hd__o21a_1 _2328_ (.A1(_1132_),
    .A2(_1133_),
    .B1(_0570_),
    .X(_1134_));
 sky130_fd_sc_hd__o21ba_1 _2329_ (.A1(_1116_),
    .A2(_1134_),
    .B1_N(_1120_),
    .X(_1135_));
 sky130_fd_sc_hd__a211o_1 _2330_ (.A1(net1020),
    .A2(_1120_),
    .B1(_1135_),
    .C1(net147),
    .X(_0127_));
 sky130_fd_sc_hd__nand2_4 _2331_ (.A(_1006_),
    .B(_1081_),
    .Y(_1136_));
 sky130_fd_sc_hd__mux2_1 _2332_ (.A0(net93),
    .A1(net801),
    .S(_1136_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _2333_ (.A0(net88),
    .A1(net593),
    .S(_1136_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _2334_ (.A0(net83),
    .A1(net923),
    .S(_1136_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _2335_ (.A0(net80),
    .A1(net483),
    .S(_1136_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _2336_ (.A0(net75),
    .A1(net589),
    .S(_1136_),
    .X(_0132_));
 sky130_fd_sc_hd__mux2_1 _2337_ (.A0(net72),
    .A1(net921),
    .S(_1136_),
    .X(_0133_));
 sky130_fd_sc_hd__nand2_2 _2338_ (.A(_1009_),
    .B(_1100_),
    .Y(_1137_));
 sky130_fd_sc_hd__a31o_1 _2339_ (.A1(net94),
    .A2(_1009_),
    .A3(_1100_),
    .B1(net147),
    .X(_1138_));
 sky130_fd_sc_hd__a21o_1 _2340_ (.A1(net961),
    .A2(_1137_),
    .B1(_1138_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _2341_ (.A0(net90),
    .A1(net1069),
    .S(_1137_),
    .X(_1139_));
 sky130_fd_sc_hd__or2_1 _2342_ (.A(net147),
    .B(net1070),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _2343_ (.A0(net87),
    .A1(net1058),
    .S(_1137_),
    .X(_1140_));
 sky130_fd_sc_hd__or2_1 _2344_ (.A(net147),
    .B(_1140_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _2345_ (.A0(net82),
    .A1(net1061),
    .S(_1137_),
    .X(_1141_));
 sky130_fd_sc_hd__or2_1 _2346_ (.A(net147),
    .B(net1062),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _2347_ (.A0(net78),
    .A1(net1073),
    .S(_1137_),
    .X(_1142_));
 sky130_fd_sc_hd__or2_1 _2348_ (.A(net147),
    .B(_1142_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _2349_ (.A0(net74),
    .A1(net1078),
    .S(_1137_),
    .X(_1143_));
 sky130_fd_sc_hd__or2_1 _2350_ (.A(net147),
    .B(net1079),
    .X(_0139_));
 sky130_fd_sc_hd__nor2_2 _2351_ (.A(_0994_),
    .B(_1101_),
    .Y(_1144_));
 sky130_fd_sc_hd__or2_1 _2352_ (.A(_0994_),
    .B(_1101_),
    .X(_1145_));
 sky130_fd_sc_hd__or2_1 _2353_ (.A(net95),
    .B(_1145_),
    .X(_1146_));
 sky130_fd_sc_hd__o211a_1 _2354_ (.A1(net1163),
    .A2(_1144_),
    .B1(_1146_),
    .C1(net156),
    .X(_0140_));
 sky130_fd_sc_hd__or2_1 _2355_ (.A(net90),
    .B(_1145_),
    .X(_1147_));
 sky130_fd_sc_hd__o211a_1 _2356_ (.A1(net1172),
    .A2(_1144_),
    .B1(_1147_),
    .C1(net156),
    .X(_0141_));
 sky130_fd_sc_hd__or2_1 _2357_ (.A(net86),
    .B(_1145_),
    .X(_1148_));
 sky130_fd_sc_hd__o211a_1 _2358_ (.A1(net1159),
    .A2(_1144_),
    .B1(_1148_),
    .C1(net156),
    .X(_0142_));
 sky130_fd_sc_hd__or2_1 _2359_ (.A(_1001_),
    .B(_1145_),
    .X(_1149_));
 sky130_fd_sc_hd__o211a_1 _2360_ (.A1(net1134),
    .A2(_1144_),
    .B1(_1149_),
    .C1(net157),
    .X(_0143_));
 sky130_fd_sc_hd__or2_1 _2361_ (.A(net77),
    .B(_1145_),
    .X(_1150_));
 sky130_fd_sc_hd__o211a_1 _2362_ (.A1(net1140),
    .A2(_1144_),
    .B1(_1150_),
    .C1(net157),
    .X(_0144_));
 sky130_fd_sc_hd__or2_1 _2363_ (.A(net73),
    .B(_1145_),
    .X(_1151_));
 sky130_fd_sc_hd__o211a_1 _2364_ (.A1(net1173),
    .A2(_1144_),
    .B1(_1151_),
    .C1(net157),
    .X(_0145_));
 sky130_fd_sc_hd__nand2_4 _2365_ (.A(_1006_),
    .B(_1085_),
    .Y(_1152_));
 sky130_fd_sc_hd__mux2_1 _2366_ (.A0(net93),
    .A1(net843),
    .S(_1152_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _2367_ (.A0(net88),
    .A1(net501),
    .S(_1152_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _2368_ (.A0(net83),
    .A1(net955),
    .S(_1152_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _2369_ (.A0(net80),
    .A1(net469),
    .S(_1152_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _2370_ (.A0(net75),
    .A1(net671),
    .S(_1152_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _2371_ (.A0(net72),
    .A1(net853),
    .S(_1152_),
    .X(_0151_));
 sky130_fd_sc_hd__nor2_2 _2372_ (.A(_1101_),
    .B(_1103_),
    .Y(_1153_));
 sky130_fd_sc_hd__mux2_1 _2373_ (.A0(net375),
    .A1(net94),
    .S(_1153_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _2374_ (.A0(net215),
    .A1(net90),
    .S(_1153_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _2375_ (.A0(net311),
    .A1(net87),
    .S(_1153_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _2376_ (.A0(net293),
    .A1(net82),
    .S(_1153_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _2377_ (.A0(net265),
    .A1(net78),
    .S(_1153_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _2378_ (.A0(net235),
    .A1(net74),
    .S(_1153_),
    .X(_0157_));
 sky130_fd_sc_hd__nand2_4 _2379_ (.A(_1005_),
    .B(_1074_),
    .Y(_1154_));
 sky130_fd_sc_hd__mux2_1 _2380_ (.A0(_0998_),
    .A1(net925),
    .S(_1154_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _2381_ (.A0(net89),
    .A1(net641),
    .S(_1154_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _2382_ (.A0(net83),
    .A1(net913),
    .S(_1154_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _2383_ (.A0(net79),
    .A1(net813),
    .S(_1154_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _2384_ (.A0(net76),
    .A1(net687),
    .S(_1154_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _2385_ (.A0(net71),
    .A1(net679),
    .S(_1154_),
    .X(_0163_));
 sky130_fd_sc_hd__or2_4 _2386_ (.A(_0994_),
    .B(_1007_),
    .X(_1155_));
 sky130_fd_sc_hd__mux2_1 _2387_ (.A0(net93),
    .A1(net929),
    .S(_1155_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_1 _2388_ (.A0(net88),
    .A1(net931),
    .S(_1155_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _2389_ (.A0(net85),
    .A1(net541),
    .S(_1155_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _2390_ (.A0(net80),
    .A1(net967),
    .S(_1155_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _2391_ (.A0(net75),
    .A1(net741),
    .S(_1155_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _2392_ (.A0(net72),
    .A1(net471),
    .S(_1155_),
    .X(_0169_));
 sky130_fd_sc_hd__nand2_4 _2393_ (.A(_1074_),
    .B(_1081_),
    .Y(_1156_));
 sky130_fd_sc_hd__mux2_1 _2394_ (.A0(net92),
    .A1(net951),
    .S(_1156_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _2395_ (.A0(net89),
    .A1(net817),
    .S(_1156_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _2396_ (.A0(net84),
    .A1(net653),
    .S(_1156_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_1 _2397_ (.A0(net79),
    .A1(net723),
    .S(_1156_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _2398_ (.A0(net76),
    .A1(net647),
    .S(_1156_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _2399_ (.A0(net71),
    .A1(net655),
    .S(_1156_),
    .X(_0175_));
 sky130_fd_sc_hd__or2_4 _2400_ (.A(_1007_),
    .B(_1089_),
    .X(_1157_));
 sky130_fd_sc_hd__mux2_1 _2401_ (.A0(net93),
    .A1(net715),
    .S(_1157_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _2402_ (.A0(net88),
    .A1(net577),
    .S(_1157_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _2403_ (.A0(net85),
    .A1(net831),
    .S(_1157_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _2404_ (.A0(net80),
    .A1(net873),
    .S(_1157_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _2405_ (.A0(net75),
    .A1(net551),
    .S(_1157_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _2406_ (.A0(net72),
    .A1(net899),
    .S(_1157_),
    .X(_0181_));
 sky130_fd_sc_hd__nand2_4 _2407_ (.A(_1074_),
    .B(_1085_),
    .Y(_1158_));
 sky130_fd_sc_hd__mux2_1 _2408_ (.A0(net92),
    .A1(net305),
    .S(_1158_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _2409_ (.A0(net89),
    .A1(net803),
    .S(_1158_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _2410_ (.A0(net84),
    .A1(net763),
    .S(_1158_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _2411_ (.A0(net79),
    .A1(net887),
    .S(_1158_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _2412_ (.A0(net76),
    .A1(net533),
    .S(_1158_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _2413_ (.A0(net71),
    .A1(net833),
    .S(_1158_),
    .X(_0187_));
 sky130_fd_sc_hd__nor2_4 _2414_ (.A(_1007_),
    .B(_1103_),
    .Y(_1159_));
 sky130_fd_sc_hd__mux2_1 _2415_ (.A0(net347),
    .A1(net93),
    .S(_1159_),
    .X(_0188_));
 sky130_fd_sc_hd__mux2_1 _2416_ (.A0(net281),
    .A1(net88),
    .S(_1159_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _2417_ (.A0(net827),
    .A1(net85),
    .S(_1159_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _2418_ (.A0(net911),
    .A1(net80),
    .S(_1159_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _2419_ (.A0(net295),
    .A1(net75),
    .S(_1159_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _2420_ (.A0(net395),
    .A1(net72),
    .S(_1159_),
    .X(_0193_));
 sky130_fd_sc_hd__nor2_2 _2421_ (.A(_1079_),
    .B(_1103_),
    .Y(_1160_));
 sky130_fd_sc_hd__mux2_1 _2422_ (.A0(net321),
    .A1(net92),
    .S(_1160_),
    .X(_0194_));
 sky130_fd_sc_hd__mux2_1 _2423_ (.A0(net495),
    .A1(net89),
    .S(_1160_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _2424_ (.A0(net261),
    .A1(net83),
    .S(_1160_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2_1 _2425_ (.A0(net455),
    .A1(net79),
    .S(_1160_),
    .X(_0197_));
 sky130_fd_sc_hd__mux2_1 _2426_ (.A0(net487),
    .A1(net76),
    .S(_1160_),
    .X(_0198_));
 sky130_fd_sc_hd__mux2_1 _2427_ (.A0(net335),
    .A1(net71),
    .S(_1160_),
    .X(_0199_));
 sky130_fd_sc_hd__or4_4 _2428_ (.A(net118),
    .B(net61),
    .C(net122),
    .D(net96),
    .X(_1161_));
 sky130_fd_sc_hd__inv_2 _2429_ (.A(_1161_),
    .Y(_1162_));
 sky130_fd_sc_hd__and2_2 _2430_ (.A(_1009_),
    .B(_1162_),
    .X(_1163_));
 sky130_fd_sc_hd__mux2_1 _2431_ (.A0(net919),
    .A1(net95),
    .S(_1163_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2_1 _2432_ (.A0(net525),
    .A1(net91),
    .S(_1163_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _2433_ (.A0(net939),
    .A1(net86),
    .S(_1163_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _2434_ (.A0(net807),
    .A1(net81),
    .S(_1163_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _2435_ (.A0(net523),
    .A1(net77),
    .S(_1163_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _2436_ (.A0(net751),
    .A1(net73),
    .S(_1163_),
    .X(_0205_));
 sky130_fd_sc_hd__o311a_4 _2437_ (.A1(net147),
    .A2(_0989_),
    .A3(net101),
    .B1(_1085_),
    .C1(_1100_),
    .X(_1164_));
 sky130_fd_sc_hd__mux2_1 _2438_ (.A0(net1119),
    .A1(net94),
    .S(_1164_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _2439_ (.A0(net1146),
    .A1(net90),
    .S(_1164_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _2440_ (.A0(net1158),
    .A1(net87),
    .S(_1164_),
    .X(_0208_));
 sky130_fd_sc_hd__mux2_1 _2441_ (.A0(net1059),
    .A1(net82),
    .S(_1164_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_1 _2442_ (.A0(net1149),
    .A1(net78),
    .S(_1164_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_1 _2443_ (.A0(net1133),
    .A1(net74),
    .S(_1164_),
    .X(_0211_));
 sky130_fd_sc_hd__nand2_4 _2444_ (.A(_1081_),
    .B(net1265),
    .Y(_1165_));
 sky130_fd_sc_hd__mux2_1 _2445_ (.A0(net93),
    .A1(net753),
    .S(_1165_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_1 _2446_ (.A0(net88),
    .A1(net959),
    .S(_1165_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_1 _2447_ (.A0(net85),
    .A1(net895),
    .S(_1165_),
    .X(_0214_));
 sky130_fd_sc_hd__mux2_1 _2448_ (.A0(net80),
    .A1(net815),
    .S(_1165_),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _2449_ (.A0(net75),
    .A1(net727),
    .S(_1165_),
    .X(_0216_));
 sky130_fd_sc_hd__mux2_1 _2450_ (.A0(net72),
    .A1(net897),
    .S(_1165_),
    .X(_0217_));
 sky130_fd_sc_hd__and2_2 _2451_ (.A(_1081_),
    .B(_1162_),
    .X(_1166_));
 sky130_fd_sc_hd__mux2_1 _2452_ (.A0(net187),
    .A1(net94),
    .S(_1166_),
    .X(_0218_));
 sky130_fd_sc_hd__mux2_1 _2453_ (.A0(net211),
    .A1(net91),
    .S(_1166_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _2454_ (.A0(net183),
    .A1(net87),
    .S(_1166_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _2455_ (.A0(net493),
    .A1(net81),
    .S(_1166_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_1 _2456_ (.A0(net213),
    .A1(net77),
    .S(_1166_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_1 _2457_ (.A0(net283),
    .A1(net73),
    .S(_1166_),
    .X(_0223_));
 sky130_fd_sc_hd__nand2_4 _2458_ (.A(_1005_),
    .B(net1265),
    .Y(_1167_));
 sky130_fd_sc_hd__mux2_1 _2459_ (.A0(net93),
    .A1(net459),
    .S(_1167_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_1 _2460_ (.A0(net88),
    .A1(net511),
    .S(_1167_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _2461_ (.A0(net85),
    .A1(net871),
    .S(_1167_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_1 _2462_ (.A0(net80),
    .A1(net915),
    .S(_1167_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_1 _2463_ (.A0(net75),
    .A1(net977),
    .S(_1167_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_1 _2464_ (.A0(net72),
    .A1(net793),
    .S(_1167_),
    .X(_0229_));
 sky130_fd_sc_hd__nand2_4 _2465_ (.A(_1085_),
    .B(_1162_),
    .Y(_1168_));
 sky130_fd_sc_hd__mux2_1 _2466_ (.A0(net94),
    .A1(net445),
    .S(_1168_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_1 _2467_ (.A0(net91),
    .A1(net411),
    .S(_1168_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_1 _2468_ (.A0(net87),
    .A1(net409),
    .S(_1168_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_1 _2469_ (.A0(net81),
    .A1(net765),
    .S(_1168_),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _2470_ (.A0(net78),
    .A1(net709),
    .S(_1168_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_1 _2471_ (.A0(net73),
    .A1(net429),
    .S(_1168_),
    .X(_0235_));
 sky130_fd_sc_hd__nor2_2 _2472_ (.A(_1071_),
    .B(_1084_),
    .Y(_1169_));
 sky130_fd_sc_hd__mux2_1 _2473_ (.A0(net485),
    .A1(net93),
    .S(_1169_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_1 _2474_ (.A0(net383),
    .A1(net88),
    .S(_1169_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_1 _2475_ (.A0(net349),
    .A1(net85),
    .S(_1169_),
    .X(_0238_));
 sky130_fd_sc_hd__mux2_1 _2476_ (.A0(net317),
    .A1(net80),
    .S(_1169_),
    .X(_0239_));
 sky130_fd_sc_hd__mux2_1 _2477_ (.A0(net649),
    .A1(net75),
    .S(_1169_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _2478_ (.A0(net531),
    .A1(net72),
    .S(_1169_),
    .X(_0241_));
 sky130_fd_sc_hd__and3_4 _2479_ (.A(_0557_),
    .B(net120),
    .C(_1073_),
    .X(_1170_));
 sky130_fd_sc_hd__or4b_4 _2480_ (.A(net118),
    .B(net61),
    .C(net96),
    .D_N(net122),
    .X(_1171_));
 sky130_fd_sc_hd__nor2_2 _2481_ (.A(_1103_),
    .B(_1171_),
    .Y(_1172_));
 sky130_fd_sc_hd__mux2_1 _2482_ (.A0(net559),
    .A1(net95),
    .S(_1172_),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _2483_ (.A0(net231),
    .A1(net90),
    .S(_1172_),
    .X(_0243_));
 sky130_fd_sc_hd__mux2_1 _2484_ (.A0(net247),
    .A1(net86),
    .S(_1172_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _2485_ (.A0(net431),
    .A1(net81),
    .S(_1172_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _2486_ (.A0(net239),
    .A1(net77),
    .S(_1172_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _2487_ (.A0(net207),
    .A1(net73),
    .S(_1172_),
    .X(_0247_));
 sky130_fd_sc_hd__nand2_4 _2488_ (.A(_1005_),
    .B(_1100_),
    .Y(_1173_));
 sky130_fd_sc_hd__mux2_1 _2489_ (.A0(net94),
    .A1(net403),
    .S(_1173_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _2490_ (.A0(net90),
    .A1(net627),
    .S(_1173_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _2491_ (.A0(net87),
    .A1(net859),
    .S(_1173_),
    .X(_0250_));
 sky130_fd_sc_hd__mux2_1 _2492_ (.A0(net82),
    .A1(net619),
    .S(_1173_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _2493_ (.A0(net78),
    .A1(net507),
    .S(_1173_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _2494_ (.A0(net74),
    .A1(net865),
    .S(_1173_),
    .X(_0253_));
 sky130_fd_sc_hd__and3_1 _2495_ (.A(net151),
    .B(\ROM_dest[1] ),
    .C(_0574_),
    .X(_1174_));
 sky130_fd_sc_hd__or4b_1 _2496_ (.A(\ROM_dest[2] ),
    .B(net106),
    .C(_0635_),
    .D_N(_1174_),
    .X(_1175_));
 sky130_fd_sc_hd__or2_1 _2497_ (.A(_0634_),
    .B(_1175_),
    .X(_1176_));
 sky130_fd_sc_hd__mux2_1 _2498_ (.A0(net13),
    .A1(net1001),
    .S(_1176_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _2499_ (.A0(net14),
    .A1(net1011),
    .S(_1176_),
    .X(_0255_));
 sky130_fd_sc_hd__nand2_4 _2500_ (.A(_1009_),
    .B(_1083_),
    .Y(_1177_));
 sky130_fd_sc_hd__mux2_1 _2501_ (.A0(net92),
    .A1(net775),
    .S(_1177_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _2502_ (.A0(net88),
    .A1(net781),
    .S(_1177_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _2503_ (.A0(net84),
    .A1(net659),
    .S(_1177_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _2504_ (.A0(net80),
    .A1(net453),
    .S(_1177_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _2505_ (.A0(net75),
    .A1(net665),
    .S(_1177_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _2506_ (.A0(net72),
    .A1(net841),
    .S(_1177_),
    .X(_0261_));
 sky130_fd_sc_hd__nor2_2 _2507_ (.A(_1103_),
    .B(_1161_),
    .Y(_1178_));
 sky130_fd_sc_hd__mux2_1 _2508_ (.A0(net371),
    .A1(net95),
    .S(_1178_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _2509_ (.A0(net693),
    .A1(net91),
    .S(_1178_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _2510_ (.A0(net465),
    .A1(net86),
    .S(_1178_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _2511_ (.A0(net299),
    .A1(net81),
    .S(_1178_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _2512_ (.A0(net189),
    .A1(net77),
    .S(_1178_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _2513_ (.A0(net461),
    .A1(net73),
    .S(_1178_),
    .X(_0267_));
 sky130_fd_sc_hd__nor2_2 _2514_ (.A(_0994_),
    .B(_1084_),
    .Y(_1179_));
 sky130_fd_sc_hd__mux2_1 _2515_ (.A0(net433),
    .A1(net92),
    .S(_1179_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _2516_ (.A0(net327),
    .A1(net88),
    .S(_1179_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _2517_ (.A0(net389),
    .A1(net84),
    .S(_1179_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _2518_ (.A0(net663),
    .A1(net80),
    .S(_1179_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _2519_ (.A0(net279),
    .A1(net75),
    .S(_1179_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2_1 _2520_ (.A0(net707),
    .A1(net72),
    .S(_1179_),
    .X(_0273_));
 sky130_fd_sc_hd__nor2_2 _2521_ (.A(_0994_),
    .B(_1171_),
    .Y(_1180_));
 sky130_fd_sc_hd__mux2_1 _2522_ (.A0(net703),
    .A1(net95),
    .S(_1180_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _2523_ (.A0(net315),
    .A1(net91),
    .S(_1180_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _2524_ (.A0(net359),
    .A1(net86),
    .S(_1180_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _2525_ (.A0(net255),
    .A1(net81),
    .S(_1180_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _2526_ (.A0(net473),
    .A1(net77),
    .S(_1180_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _2527_ (.A0(net503),
    .A1(net73),
    .S(_1180_),
    .X(_0279_));
 sky130_fd_sc_hd__and2_2 _2528_ (.A(_1005_),
    .B(_1162_),
    .X(_1181_));
 sky130_fd_sc_hd__mux2_1 _2529_ (.A0(net195),
    .A1(net95),
    .S(_1181_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_1 _2530_ (.A0(net275),
    .A1(net91),
    .S(_1181_),
    .X(_0281_));
 sky130_fd_sc_hd__mux2_1 _2531_ (.A0(net423),
    .A1(net86),
    .S(_1181_),
    .X(_0282_));
 sky130_fd_sc_hd__mux2_1 _2532_ (.A0(net699),
    .A1(net81),
    .S(_1181_),
    .X(_0283_));
 sky130_fd_sc_hd__mux2_1 _2533_ (.A0(net451),
    .A1(net78),
    .S(_1181_),
    .X(_0284_));
 sky130_fd_sc_hd__mux2_1 _2534_ (.A0(net467),
    .A1(net73),
    .S(_1181_),
    .X(_0285_));
 sky130_fd_sc_hd__nor2_4 _2535_ (.A(_1084_),
    .B(_1089_),
    .Y(_1182_));
 sky130_fd_sc_hd__mux2_1 _2536_ (.A0(net337),
    .A1(net92),
    .S(_1182_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _2537_ (.A0(net245),
    .A1(net88),
    .S(_1182_),
    .X(_0287_));
 sky130_fd_sc_hd__mux2_1 _2538_ (.A0(net391),
    .A1(net84),
    .S(_1182_),
    .X(_0288_));
 sky130_fd_sc_hd__mux2_1 _2539_ (.A0(net443),
    .A1(net79),
    .S(_1182_),
    .X(_0289_));
 sky130_fd_sc_hd__mux2_1 _2540_ (.A0(net273),
    .A1(net75),
    .S(_1182_),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _2541_ (.A0(net193),
    .A1(net71),
    .S(_1182_),
    .X(_0291_));
 sky130_fd_sc_hd__nand2_4 _2542_ (.A(_1009_),
    .B(_1170_),
    .Y(_1183_));
 sky130_fd_sc_hd__mux2_1 _2543_ (.A0(net95),
    .A1(net819),
    .S(_1183_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _2544_ (.A0(net91),
    .A1(net905),
    .S(_1183_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _2545_ (.A0(net86),
    .A1(net829),
    .S(_1183_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _2546_ (.A0(net81),
    .A1(net617),
    .S(_1183_),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _2547_ (.A0(net77),
    .A1(net907),
    .S(_1183_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _2548_ (.A0(net73),
    .A1(net847),
    .S(_1183_),
    .X(_0297_));
 sky130_fd_sc_hd__nor2_2 _2549_ (.A(_1084_),
    .B(_1103_),
    .Y(_1184_));
 sky130_fd_sc_hd__mux2_1 _2550_ (.A0(net197),
    .A1(net92),
    .S(_1184_),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _2551_ (.A0(net379),
    .A1(net88),
    .S(_1184_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _2552_ (.A0(net297),
    .A1(net84),
    .S(_1184_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _2553_ (.A0(net191),
    .A1(net80),
    .S(_1184_),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _2554_ (.A0(net397),
    .A1(net76),
    .S(_1184_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _2555_ (.A0(net499),
    .A1(net72),
    .S(_1184_),
    .X(_0303_));
 sky130_fd_sc_hd__nor2_2 _2556_ (.A(_1071_),
    .B(_1171_),
    .Y(_1185_));
 sky130_fd_sc_hd__mux2_1 _2557_ (.A0(net361),
    .A1(net95),
    .S(_1185_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _2558_ (.A0(net319),
    .A1(net91),
    .S(_1185_),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _2559_ (.A0(net413),
    .A1(net86),
    .S(_1185_),
    .X(_0306_));
 sky130_fd_sc_hd__mux2_1 _2560_ (.A0(net287),
    .A1(net81),
    .S(_1185_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _2561_ (.A0(net421),
    .A1(net77),
    .S(_1185_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _2562_ (.A0(net603),
    .A1(net73),
    .S(_1185_),
    .X(_0309_));
 sky130_fd_sc_hd__nand2_4 _2563_ (.A(_1078_),
    .B(_1085_),
    .Y(_1186_));
 sky130_fd_sc_hd__mux2_1 _2564_ (.A0(net92),
    .A1(net891),
    .S(_1186_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _2565_ (.A0(net89),
    .A1(net821),
    .S(_1186_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _2566_ (.A0(net83),
    .A1(net805),
    .S(_1186_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _2567_ (.A0(net79),
    .A1(net605),
    .S(_1186_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _2568_ (.A0(net76),
    .A1(net631),
    .S(_1186_),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _2569_ (.A0(net71),
    .A1(net879),
    .S(_1186_),
    .X(_0315_));
 sky130_fd_sc_hd__nand2_4 _2570_ (.A(_1005_),
    .B(_1170_),
    .Y(_1187_));
 sky130_fd_sc_hd__mux2_1 _2571_ (.A0(net95),
    .A1(net623),
    .S(_1187_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _2572_ (.A0(net91),
    .A1(net357),
    .S(_1187_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_1 _2573_ (.A0(net86),
    .A1(net725),
    .S(_1187_),
    .X(_0318_));
 sky130_fd_sc_hd__mux2_1 _2574_ (.A0(net81),
    .A1(net401),
    .S(_1187_),
    .X(_0319_));
 sky130_fd_sc_hd__mux2_1 _2575_ (.A0(net77),
    .A1(net399),
    .S(_1187_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _2576_ (.A0(net73),
    .A1(net607),
    .S(_1187_),
    .X(_0321_));
 sky130_fd_sc_hd__nand2_4 _2577_ (.A(_1078_),
    .B(_1081_),
    .Y(_1188_));
 sky130_fd_sc_hd__mux2_1 _2578_ (.A0(net92),
    .A1(net901),
    .S(_1188_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_1 _2579_ (.A0(net89),
    .A1(net893),
    .S(_1188_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_1 _2580_ (.A0(net83),
    .A1(net539),
    .S(_1188_),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_1 _2581_ (.A0(net79),
    .A1(net685),
    .S(_1188_),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _2582_ (.A0(net76),
    .A1(net519),
    .S(_1188_),
    .X(_0326_));
 sky130_fd_sc_hd__mux2_1 _2583_ (.A0(net71),
    .A1(net621),
    .S(_1188_),
    .X(_0327_));
 sky130_fd_sc_hd__nand2_2 _2584_ (.A(_1081_),
    .B(_1170_),
    .Y(_1189_));
 sky130_fd_sc_hd__mux2_1 _2585_ (.A0(net92),
    .A1(net405),
    .S(_1189_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _2586_ (.A0(net89),
    .A1(net549),
    .S(_1189_),
    .X(_0329_));
 sky130_fd_sc_hd__mux2_1 _2587_ (.A0(net83),
    .A1(net947),
    .S(_1189_),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _2588_ (.A0(net81),
    .A1(net975),
    .S(_1189_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _2589_ (.A0(net77),
    .A1(net969),
    .S(_1189_),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _2590_ (.A0(net73),
    .A1(net935),
    .S(_1189_),
    .X(_0333_));
 sky130_fd_sc_hd__nor2_4 _2591_ (.A(_0994_),
    .B(_1161_),
    .Y(_1190_));
 sky130_fd_sc_hd__mux2_1 _2592_ (.A0(net271),
    .A1(net95),
    .S(_1190_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2_1 _2593_ (.A0(net289),
    .A1(net91),
    .S(_1190_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _2594_ (.A0(net369),
    .A1(net87),
    .S(_1190_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _2595_ (.A0(net221),
    .A1(net81),
    .S(_1190_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_1 _2596_ (.A0(net351),
    .A1(net77),
    .S(_1190_),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_1 _2597_ (.A0(net449),
    .A1(_1003_),
    .S(_1190_),
    .X(_0339_));
 sky130_fd_sc_hd__nand2_4 _2598_ (.A(_1085_),
    .B(_1170_),
    .Y(_1191_));
 sky130_fd_sc_hd__mux2_1 _2599_ (.A0(net92),
    .A1(net437),
    .S(_1191_),
    .X(_0340_));
 sky130_fd_sc_hd__mux2_1 _2600_ (.A0(net91),
    .A1(net573),
    .S(_1191_),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_1 _2601_ (.A0(net83),
    .A1(net789),
    .S(_1191_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _2602_ (.A0(net81),
    .A1(net711),
    .S(_1191_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_1 _2603_ (.A0(net77),
    .A1(net735),
    .S(_1191_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _2604_ (.A0(net73),
    .A1(net791),
    .S(_1191_),
    .X(_0345_));
 sky130_fd_sc_hd__or2_4 _2605_ (.A(_1071_),
    .B(_1079_),
    .X(_1192_));
 sky130_fd_sc_hd__mux2_1 _2606_ (.A0(net92),
    .A1(net849),
    .S(_1192_),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _2607_ (.A0(net89),
    .A1(net643),
    .S(_1192_),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _2608_ (.A0(net83),
    .A1(net683),
    .S(_1192_),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _2609_ (.A0(net79),
    .A1(net661),
    .S(_1192_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _2610_ (.A0(net76),
    .A1(net861),
    .S(_1192_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _2611_ (.A0(net71),
    .A1(net609),
    .S(_1192_),
    .X(_0351_));
 sky130_fd_sc_hd__nor2_2 _2612_ (.A(_1075_),
    .B(_1103_),
    .Y(_1193_));
 sky130_fd_sc_hd__mux2_1 _2613_ (.A0(net225),
    .A1(net93),
    .S(_1193_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _2614_ (.A0(net333),
    .A1(net89),
    .S(_1193_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _2615_ (.A0(net285),
    .A1(net84),
    .S(_1193_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _2616_ (.A0(net669),
    .A1(_1001_),
    .S(_1193_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _2617_ (.A0(net185),
    .A1(net76),
    .S(_1193_),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _2618_ (.A0(net249),
    .A1(_1003_),
    .S(_1193_),
    .X(_0357_));
 sky130_fd_sc_hd__nand2_4 _2619_ (.A(_1009_),
    .B(_1078_),
    .Y(_1194_));
 sky130_fd_sc_hd__mux2_1 _2620_ (.A0(net92),
    .A1(net957),
    .S(_1194_),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _2621_ (.A0(net89),
    .A1(net881),
    .S(_1194_),
    .X(_0359_));
 sky130_fd_sc_hd__mux2_1 _2622_ (.A0(net83),
    .A1(net909),
    .S(_1194_),
    .X(_0360_));
 sky130_fd_sc_hd__mux2_1 _2623_ (.A0(net79),
    .A1(net889),
    .S(_1194_),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_1 _2624_ (.A0(_1002_),
    .A1(net759),
    .S(_1194_),
    .X(_0362_));
 sky130_fd_sc_hd__mux2_1 _2625_ (.A0(net71),
    .A1(net739),
    .S(_1194_),
    .X(_0363_));
 sky130_fd_sc_hd__nor2_2 _2626_ (.A(_1075_),
    .B(_1089_),
    .Y(_1195_));
 sky130_fd_sc_hd__mux2_1 _2627_ (.A0(net241),
    .A1(_0998_),
    .S(_1195_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _2628_ (.A0(net757),
    .A1(net89),
    .S(_1195_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_1 _2629_ (.A0(net439),
    .A1(net84),
    .S(_1195_),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_1 _2630_ (.A0(net205),
    .A1(net79),
    .S(_1195_),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_1 _2631_ (.A0(net387),
    .A1(net76),
    .S(_1195_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _2632_ (.A0(net545),
    .A1(net72),
    .S(_1195_),
    .X(_0369_));
 sky130_fd_sc_hd__or2_4 _2633_ (.A(_0994_),
    .B(_1079_),
    .X(_1196_));
 sky130_fd_sc_hd__mux2_1 _2634_ (.A0(net92),
    .A1(net809),
    .S(_1196_),
    .X(_0370_));
 sky130_fd_sc_hd__mux2_1 _2635_ (.A0(net89),
    .A1(net973),
    .S(_1196_),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _2636_ (.A0(net83),
    .A1(net425),
    .S(_1196_),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_1 _2637_ (.A0(net79),
    .A1(net839),
    .S(_1196_),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_1 _2638_ (.A0(_1002_),
    .A1(net777),
    .S(_1196_),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_1 _2639_ (.A0(net71),
    .A1(net689),
    .S(_1196_),
    .X(_0375_));
 sky130_fd_sc_hd__nor2_2 _2640_ (.A(_0994_),
    .B(_1075_),
    .Y(_1197_));
 sky130_fd_sc_hd__mux2_1 _2641_ (.A0(net227),
    .A1(net93),
    .S(_1197_),
    .X(_0376_));
 sky130_fd_sc_hd__mux2_1 _2642_ (.A0(net797),
    .A1(_0999_),
    .S(_1197_),
    .X(_0377_));
 sky130_fd_sc_hd__mux2_1 _2643_ (.A0(net597),
    .A1(net84),
    .S(_1197_),
    .X(_0378_));
 sky130_fd_sc_hd__mux2_1 _2644_ (.A0(net783),
    .A1(net79),
    .S(_1197_),
    .X(_0379_));
 sky130_fd_sc_hd__mux2_1 _2645_ (.A0(net329),
    .A1(net76),
    .S(_1197_),
    .X(_0380_));
 sky130_fd_sc_hd__mux2_1 _2646_ (.A0(net477),
    .A1(net71),
    .S(_1197_),
    .X(_0381_));
 sky130_fd_sc_hd__nand2_4 _2647_ (.A(_1081_),
    .B(_1100_),
    .Y(_1198_));
 sky130_fd_sc_hd__mux2_1 _2648_ (.A0(net94),
    .A1(net629),
    .S(_1198_),
    .X(_0382_));
 sky130_fd_sc_hd__mux2_1 _2649_ (.A0(net90),
    .A1(net515),
    .S(_1198_),
    .X(_0383_));
 sky130_fd_sc_hd__mux2_1 _2650_ (.A0(net87),
    .A1(net535),
    .S(_1198_),
    .X(_0384_));
 sky130_fd_sc_hd__mux2_1 _2651_ (.A0(net82),
    .A1(net633),
    .S(_1198_),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _2652_ (.A0(net78),
    .A1(net561),
    .S(_1198_),
    .X(_0386_));
 sky130_fd_sc_hd__mux2_1 _2653_ (.A0(net74),
    .A1(net575),
    .S(_1198_),
    .X(_0387_));
 sky130_fd_sc_hd__nand2_4 _2654_ (.A(_1078_),
    .B(_1088_),
    .Y(_1199_));
 sky130_fd_sc_hd__mux2_1 _2655_ (.A0(net92),
    .A1(net611),
    .S(_1199_),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _2656_ (.A0(net89),
    .A1(net547),
    .S(_1199_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _2657_ (.A0(net83),
    .A1(net291),
    .S(_1199_),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _2658_ (.A0(net79),
    .A1(net481),
    .S(_1199_),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_1 _2659_ (.A0(net76),
    .A1(net571),
    .S(_1199_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _2660_ (.A0(net71),
    .A1(net479),
    .S(_1199_),
    .X(_0393_));
 sky130_fd_sc_hd__nor2_2 _2661_ (.A(_1089_),
    .B(_1161_),
    .Y(_1200_));
 sky130_fd_sc_hd__mux2_1 _2662_ (.A0(net415),
    .A1(net95),
    .S(_1200_),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_1 _2663_ (.A0(net331),
    .A1(net91),
    .S(_1200_),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _2664_ (.A0(net381),
    .A1(net86),
    .S(_1200_),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_1 _2665_ (.A0(net565),
    .A1(net81),
    .S(_1200_),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _2666_ (.A0(net341),
    .A1(net77),
    .S(_1200_),
    .X(_0398_));
 sky130_fd_sc_hd__mux2_1 _2667_ (.A0(net393),
    .A1(net73),
    .S(_1200_),
    .X(_0399_));
 sky130_fd_sc_hd__and2_4 _2668_ (.A(_0578_),
    .B(_0591_),
    .X(_1201_));
 sky130_fd_sc_hd__and3_2 _2669_ (.A(_0550_),
    .B(_0578_),
    .C(_0591_),
    .X(_1202_));
 sky130_fd_sc_hd__or3_1 _2670_ (.A(\insin[0] ),
    .B(\insin[1] ),
    .C(\insin[2] ),
    .X(_1203_));
 sky130_fd_sc_hd__and2_1 _2671_ (.A(\A[5] ),
    .B(_0742_),
    .X(_1204_));
 sky130_fd_sc_hd__nor2_1 _2672_ (.A(\A[5] ),
    .B(_0742_),
    .Y(_1205_));
 sky130_fd_sc_hd__or2_1 _2673_ (.A(_1204_),
    .B(_1205_),
    .X(_1206_));
 sky130_fd_sc_hd__and2b_1 _2674_ (.A_N(_0692_),
    .B(\A[4] ),
    .X(_1207_));
 sky130_fd_sc_hd__and2_1 _2675_ (.A(\A[4] ),
    .B(_0692_),
    .X(_1208_));
 sky130_fd_sc_hd__or2_1 _2676_ (.A(\A[4] ),
    .B(_0692_),
    .X(_1209_));
 sky130_fd_sc_hd__nand2b_2 _2677_ (.A_N(_1208_),
    .B(_1209_),
    .Y(_1210_));
 sky130_fd_sc_hd__and2b_1 _2678_ (.A_N(_0947_),
    .B(\A[3] ),
    .X(_1211_));
 sky130_fd_sc_hd__and2_1 _2679_ (.A(\A[2] ),
    .B(_0897_),
    .X(_1212_));
 sky130_fd_sc_hd__or2_1 _2680_ (.A(\A[2] ),
    .B(_0897_),
    .X(_1213_));
 sky130_fd_sc_hd__xnor2_4 _2681_ (.A(\A[2] ),
    .B(_0897_),
    .Y(_1214_));
 sky130_fd_sc_hd__nand3_2 _2682_ (.A(\A[1] ),
    .B(_0845_),
    .C(_0846_),
    .Y(_1215_));
 sky130_fd_sc_hd__a21o_1 _2683_ (.A1(_0845_),
    .A2(_0846_),
    .B1(\A[1] ),
    .X(_1216_));
 sky130_fd_sc_hd__nand2_1 _2684_ (.A(_1215_),
    .B(_1216_),
    .Y(_1217_));
 sky130_fd_sc_hd__a21bo_1 _2685_ (.A1(_0794_),
    .A2(_0795_),
    .B1_N(\A[0] ),
    .X(_1218_));
 sky130_fd_sc_hd__a21oi_2 _2686_ (.A1(_1215_),
    .A2(_1216_),
    .B1(_1218_),
    .Y(_1219_));
 sky130_fd_sc_hd__and2_1 _2687_ (.A(\A[1] ),
    .B(_0847_),
    .X(_1220_));
 sky130_fd_sc_hd__o21ai_2 _2688_ (.A1(_1219_),
    .A2(_1220_),
    .B1(_1214_),
    .Y(_1221_));
 sky130_fd_sc_hd__nand2_1 _2689_ (.A(\A[2] ),
    .B(_0898_),
    .Y(_1222_));
 sky130_fd_sc_hd__and2_1 _2690_ (.A(\A[3] ),
    .B(_0947_),
    .X(_1223_));
 sky130_fd_sc_hd__or2_1 _2691_ (.A(\A[3] ),
    .B(_0947_),
    .X(_1224_));
 sky130_fd_sc_hd__xnor2_4 _2692_ (.A(\A[3] ),
    .B(_0947_),
    .Y(_1225_));
 sky130_fd_sc_hd__inv_2 _2693_ (.A(_1225_),
    .Y(_1226_));
 sky130_fd_sc_hd__a31oi_2 _2694_ (.A1(\A[2] ),
    .A2(_0898_),
    .A3(_1225_),
    .B1(_1211_),
    .Y(_1227_));
 sky130_fd_sc_hd__o211ai_2 _2695_ (.A1(_1219_),
    .A2(_1220_),
    .B1(_1225_),
    .C1(_1214_),
    .Y(_1228_));
 sky130_fd_sc_hd__nand2_1 _2696_ (.A(_1227_),
    .B(_1228_),
    .Y(_1229_));
 sky130_fd_sc_hd__a21boi_1 _2697_ (.A1(_1227_),
    .A2(_1228_),
    .B1_N(_1210_),
    .Y(_1230_));
 sky130_fd_sc_hd__or3_1 _2698_ (.A(_1206_),
    .B(_1207_),
    .C(_1230_),
    .X(_1231_));
 sky130_fd_sc_hd__o21ai_2 _2699_ (.A1(_1207_),
    .A2(_1230_),
    .B1(_1206_),
    .Y(_1232_));
 sky130_fd_sc_hd__xor2_2 _2700_ (.A(_1210_),
    .B(_1229_),
    .X(_1233_));
 sky130_fd_sc_hd__xnor2_2 _2701_ (.A(\A[0] ),
    .B(_0796_),
    .Y(_1234_));
 sky130_fd_sc_hd__and2_1 _2702_ (.A(_1217_),
    .B(_1234_),
    .X(_1235_));
 sky130_fd_sc_hd__or3_1 _2703_ (.A(_1214_),
    .B(_1219_),
    .C(_1220_),
    .X(_1236_));
 sky130_fd_sc_hd__and3_1 _2704_ (.A(_1221_),
    .B(_1235_),
    .C(_1236_),
    .X(_1237_));
 sky130_fd_sc_hd__nand3_1 _2705_ (.A(_1221_),
    .B(_1222_),
    .C(_1226_),
    .Y(_1238_));
 sky130_fd_sc_hd__a21o_1 _2706_ (.A1(_1221_),
    .A2(_1222_),
    .B1(_1226_),
    .X(_1239_));
 sky130_fd_sc_hd__and3_1 _2707_ (.A(_1237_),
    .B(_1238_),
    .C(_1239_),
    .X(_1240_));
 sky130_fd_sc_hd__nand2_1 _2708_ (.A(_1233_),
    .B(_1240_),
    .Y(_1241_));
 sky130_fd_sc_hd__and4_1 _2709_ (.A(_1231_),
    .B(_1232_),
    .C(_1233_),
    .D(_1240_),
    .X(_1242_));
 sky130_fd_sc_hd__nor2_1 _2710_ (.A(_1203_),
    .B(_1242_),
    .Y(_1243_));
 sky130_fd_sc_hd__o21ai_1 _2711_ (.A1(_0547_),
    .A2(_0742_),
    .B1(_1232_),
    .Y(_1244_));
 sky130_fd_sc_hd__or3_1 _2712_ (.A(_0548_),
    .B(\insin[1] ),
    .C(\insin[2] ),
    .X(_1245_));
 sky130_fd_sc_hd__or3b_1 _2713_ (.A(_1242_),
    .B(_1245_),
    .C_N(_1244_),
    .X(_1246_));
 sky130_fd_sc_hd__xnor2_1 _2714_ (.A(_0953_),
    .B(_1234_),
    .Y(_1247_));
 sky130_fd_sc_hd__nor2_1 _2715_ (.A(net51),
    .B(_1247_),
    .Y(_1248_));
 sky130_fd_sc_hd__nand2_2 _2716_ (.A(net51),
    .B(_1247_),
    .Y(_1249_));
 sky130_fd_sc_hd__nand2_2 _2717_ (.A(net1223),
    .B(net1160),
    .Y(_1250_));
 sky130_fd_sc_hd__or3b_1 _2718_ (.A(_1248_),
    .B(_1250_),
    .C_N(_1249_),
    .X(_1251_));
 sky130_fd_sc_hd__nor2_2 _2719_ (.A(\insin[2] ),
    .B(_0595_),
    .Y(_1252_));
 sky130_fd_sc_hd__and3_1 _2720_ (.A(\A[0] ),
    .B(_0794_),
    .C(_0795_),
    .X(_1253_));
 sky130_fd_sc_hd__nand2_1 _2721_ (.A(_1252_),
    .B(_1253_),
    .Y(_1254_));
 sky130_fd_sc_hd__or3_2 _2722_ (.A(\insin[0] ),
    .B(\insin[1] ),
    .C(_0549_),
    .X(_1255_));
 sky130_fd_sc_hd__inv_2 _2723_ (.A(_1255_),
    .Y(_1256_));
 sky130_fd_sc_hd__o211a_1 _2724_ (.A1(\insin[0] ),
    .A2(_1234_),
    .B1(_1254_),
    .C1(_1203_),
    .X(_1257_));
 sky130_fd_sc_hd__a31o_1 _2725_ (.A1(_1246_),
    .A2(_1251_),
    .A3(_1257_),
    .B1(_1243_),
    .X(_1258_));
 sky130_fd_sc_hd__nand2_1 _2726_ (.A(_1202_),
    .B(_1258_),
    .Y(_1259_));
 sky130_fd_sc_hd__o21a_2 _2727_ (.A1(\insin[4] ),
    .A2(_0579_),
    .B1(_0609_),
    .X(_1260_));
 sky130_fd_sc_hd__mux2_1 _2728_ (.A0(_0796_),
    .A1(net1086),
    .S(_1260_),
    .X(_1261_));
 sky130_fd_sc_hd__o211a_1 _2729_ (.A1(_1202_),
    .A2(_1261_),
    .B1(_1259_),
    .C1(net114),
    .X(_1262_));
 sky130_fd_sc_hd__a21oi_4 _2730_ (.A1(_0639_),
    .A2(net103),
    .B1(net102),
    .Y(_1263_));
 sky130_fd_sc_hd__a21o_2 _2731_ (.A1(_0639_),
    .A2(net103),
    .B1(net102),
    .X(_1264_));
 sky130_fd_sc_hd__a21o_1 _2732_ (.A1(net144),
    .A2(net585),
    .B1(_1264_),
    .X(_1265_));
 sky130_fd_sc_hd__o221a_1 _2733_ (.A1(net1086),
    .A2(_1263_),
    .B1(_1265_),
    .B2(_1262_),
    .C1(net150),
    .X(_0400_));
 sky130_fd_sc_hd__and3_1 _2734_ (.A(_1215_),
    .B(_1216_),
    .C(_1218_),
    .X(_1266_));
 sky130_fd_sc_hd__or2_1 _2735_ (.A(_1219_),
    .B(_1266_),
    .X(_1267_));
 sky130_fd_sc_hd__xor2_1 _2736_ (.A(_1217_),
    .B(_1253_),
    .X(_1268_));
 sky130_fd_sc_hd__mux2_1 _2737_ (.A0(_1267_),
    .A1(_1268_),
    .S(_0954_),
    .X(_1269_));
 sky130_fd_sc_hd__nor2_1 _2738_ (.A(_1249_),
    .B(_1269_),
    .Y(_1270_));
 sky130_fd_sc_hd__a21o_1 _2739_ (.A1(_1249_),
    .A2(_1269_),
    .B1(_1250_),
    .X(_1271_));
 sky130_fd_sc_hd__and2b_1 _2740_ (.A_N(_1234_),
    .B(_1267_),
    .X(_1272_));
 sky130_fd_sc_hd__or2_2 _2741_ (.A(_0549_),
    .B(_0592_),
    .X(_1273_));
 sky130_fd_sc_hd__or3_1 _2742_ (.A(\insin[2] ),
    .B(_0595_),
    .C(_1215_),
    .X(_1274_));
 sky130_fd_sc_hd__o211a_1 _2743_ (.A1(_0990_),
    .A2(_1217_),
    .B1(_1274_),
    .C1(_1201_),
    .X(_1275_));
 sky130_fd_sc_hd__o32a_1 _2744_ (.A1(_1235_),
    .A2(_1272_),
    .A3(_1273_),
    .B1(_1255_),
    .B2(_1268_),
    .X(_1276_));
 sky130_fd_sc_hd__o211a_1 _2745_ (.A1(_1270_),
    .A2(_1271_),
    .B1(_1275_),
    .C1(_1276_),
    .X(_1277_));
 sky130_fd_sc_hd__inv_2 _2746_ (.A(_1277_),
    .Y(_1278_));
 sky130_fd_sc_hd__mux2_1 _2747_ (.A0(_0848_),
    .A1(net1096),
    .S(_1260_),
    .X(_1279_));
 sky130_fd_sc_hd__o221a_1 _2748_ (.A1(\insin[4] ),
    .A2(_1278_),
    .B1(_1279_),
    .B2(_1202_),
    .C1(net114),
    .X(_1280_));
 sky130_fd_sc_hd__a21o_1 _2749_ (.A1(net144),
    .A2(net761),
    .B1(_1264_),
    .X(_1281_));
 sky130_fd_sc_hd__o221a_1 _2750_ (.A1(net1096),
    .A2(_1263_),
    .B1(_1280_),
    .B2(_1281_),
    .C1(net150),
    .X(_0401_));
 sky130_fd_sc_hd__mux2_1 _2751_ (.A0(_0897_),
    .A1(net1101),
    .S(_1260_),
    .X(_1282_));
 sky130_fd_sc_hd__inv_2 _2752_ (.A(_1282_),
    .Y(_1283_));
 sky130_fd_sc_hd__a21bo_1 _2753_ (.A1(_1216_),
    .A2(_1253_),
    .B1_N(_1215_),
    .X(_1284_));
 sky130_fd_sc_hd__xor2_1 _2754_ (.A(_1214_),
    .B(_1284_),
    .X(_1285_));
 sky130_fd_sc_hd__nand3_1 _2755_ (.A(_0953_),
    .B(_1221_),
    .C(_1236_),
    .Y(_1286_));
 sky130_fd_sc_hd__or2_1 _2756_ (.A(_0953_),
    .B(_1285_),
    .X(_1287_));
 sky130_fd_sc_hd__o211a_1 _2757_ (.A1(_1249_),
    .A2(_1269_),
    .B1(_1286_),
    .C1(_1287_),
    .X(_1288_));
 sky130_fd_sc_hd__a211oi_2 _2758_ (.A1(_1286_),
    .A2(_1287_),
    .B1(_1249_),
    .C1(_1269_),
    .Y(_1289_));
 sky130_fd_sc_hd__nand2_1 _2759_ (.A(_1212_),
    .B(_1252_),
    .Y(_1290_));
 sky130_fd_sc_hd__o221a_1 _2760_ (.A1(_0990_),
    .A2(_1214_),
    .B1(_1255_),
    .B2(_1285_),
    .C1(_1290_),
    .X(_1291_));
 sky130_fd_sc_hd__a21oi_1 _2761_ (.A1(_1221_),
    .A2(_1236_),
    .B1(_1235_),
    .Y(_1292_));
 sky130_fd_sc_hd__or3_1 _2762_ (.A(_1237_),
    .B(_1273_),
    .C(_1292_),
    .X(_1293_));
 sky130_fd_sc_hd__o311a_1 _2763_ (.A1(_1250_),
    .A2(_1288_),
    .A3(_1289_),
    .B1(_1291_),
    .C1(_1293_),
    .X(_1294_));
 sky130_fd_sc_hd__mux2_1 _2764_ (.A0(_1283_),
    .A1(_1294_),
    .S(_1202_),
    .X(_1295_));
 sky130_fd_sc_hd__nor2_1 _2765_ (.A(net144),
    .B(_1295_),
    .Y(_1296_));
 sky130_fd_sc_hd__a21o_1 _2766_ (.A1(net144),
    .A2(net885),
    .B1(_1264_),
    .X(_1297_));
 sky130_fd_sc_hd__o221a_1 _2767_ (.A1(net1101),
    .A2(_1263_),
    .B1(_1296_),
    .B2(_1297_),
    .C1(net150),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _2768_ (.A0(_0947_),
    .A1(net1071),
    .S(_1260_),
    .X(_1298_));
 sky130_fd_sc_hd__inv_2 _2769_ (.A(_1298_),
    .Y(_1299_));
 sky130_fd_sc_hd__a21o_1 _2770_ (.A1(_1213_),
    .A2(_1284_),
    .B1(_1212_),
    .X(_1300_));
 sky130_fd_sc_hd__xnor2_1 _2771_ (.A(_1225_),
    .B(_1300_),
    .Y(_1301_));
 sky130_fd_sc_hd__a21o_1 _2772_ (.A1(_1238_),
    .A2(_1239_),
    .B1(_0954_),
    .X(_1302_));
 sky130_fd_sc_hd__or2_1 _2773_ (.A(_0953_),
    .B(_1301_),
    .X(_1303_));
 sky130_fd_sc_hd__a21oi_1 _2774_ (.A1(_1302_),
    .A2(_1303_),
    .B1(_1289_),
    .Y(_1304_));
 sky130_fd_sc_hd__and3_1 _2775_ (.A(_1289_),
    .B(_1302_),
    .C(_1303_),
    .X(_1305_));
 sky130_fd_sc_hd__a2bb2o_1 _2776_ (.A1_N(_0990_),
    .A2_N(_1225_),
    .B1(_1252_),
    .B2(_1223_),
    .X(_1306_));
 sky130_fd_sc_hd__a21oi_1 _2777_ (.A1(_1256_),
    .A2(_1301_),
    .B1(_1306_),
    .Y(_1307_));
 sky130_fd_sc_hd__a21oi_1 _2778_ (.A1(_1238_),
    .A2(_1239_),
    .B1(_1237_),
    .Y(_1308_));
 sky130_fd_sc_hd__or3_1 _2779_ (.A(_1240_),
    .B(_1273_),
    .C(_1308_),
    .X(_1309_));
 sky130_fd_sc_hd__o311a_1 _2780_ (.A1(_1250_),
    .A2(_1304_),
    .A3(_1305_),
    .B1(_1307_),
    .C1(_1309_),
    .X(_1310_));
 sky130_fd_sc_hd__mux2_1 _2781_ (.A0(_1299_),
    .A1(_1310_),
    .S(_1202_),
    .X(_1311_));
 sky130_fd_sc_hd__nor2_1 _2782_ (.A(net144),
    .B(_1311_),
    .Y(_1312_));
 sky130_fd_sc_hd__a21o_1 _2783_ (.A1(net144),
    .A2(net747),
    .B1(_1264_),
    .X(_1313_));
 sky130_fd_sc_hd__o221a_1 _2784_ (.A1(net1071),
    .A2(_1263_),
    .B1(_1312_),
    .B2(_1313_),
    .C1(net150),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _2785_ (.A0(_0692_),
    .A1(net1082),
    .S(_1260_),
    .X(_1314_));
 sky130_fd_sc_hd__inv_2 _2786_ (.A(_1314_),
    .Y(_1315_));
 sky130_fd_sc_hd__o21a_1 _2787_ (.A1(_1223_),
    .A2(_1300_),
    .B1(_1224_),
    .X(_1316_));
 sky130_fd_sc_hd__xnor2_1 _2788_ (.A(_1210_),
    .B(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__mux2_1 _2789_ (.A0(_1233_),
    .A1(_1317_),
    .S(_0954_),
    .X(_1318_));
 sky130_fd_sc_hd__or2_1 _2790_ (.A(_1305_),
    .B(_1318_),
    .X(_1319_));
 sky130_fd_sc_hd__a21oi_1 _2791_ (.A1(_1305_),
    .A2(_1318_),
    .B1(_1250_),
    .Y(_1320_));
 sky130_fd_sc_hd__a2bb2o_1 _2792_ (.A1_N(_0990_),
    .A2_N(_1210_),
    .B1(_1252_),
    .B2(_1208_),
    .X(_1321_));
 sky130_fd_sc_hd__o21ba_1 _2793_ (.A1(_1233_),
    .A2(_1240_),
    .B1_N(_1273_),
    .X(_1322_));
 sky130_fd_sc_hd__a221o_1 _2794_ (.A1(_1256_),
    .A2(_1317_),
    .B1(_1322_),
    .B2(_1241_),
    .C1(_1321_),
    .X(_1323_));
 sky130_fd_sc_hd__a21oi_2 _2795_ (.A1(_1319_),
    .A2(_1320_),
    .B1(_1323_),
    .Y(_1324_));
 sky130_fd_sc_hd__mux2_1 _2796_ (.A0(_1315_),
    .A1(_1324_),
    .S(_1202_),
    .X(_1325_));
 sky130_fd_sc_hd__nor2_1 _2797_ (.A(net144),
    .B(_1325_),
    .Y(_1326_));
 sky130_fd_sc_hd__a21o_1 _2798_ (.A1(net144),
    .A2(net743),
    .B1(_1264_),
    .X(_1327_));
 sky130_fd_sc_hd__o221a_1 _2799_ (.A1(net1082),
    .A2(_1263_),
    .B1(_1326_),
    .B2(_1327_),
    .C1(net150),
    .X(_0404_));
 sky130_fd_sc_hd__a21o_1 _2800_ (.A1(_1231_),
    .A2(_1232_),
    .B1(_0954_),
    .X(_1328_));
 sky130_fd_sc_hd__o21a_1 _2801_ (.A1(_1208_),
    .A2(_1316_),
    .B1(_1209_),
    .X(_1329_));
 sky130_fd_sc_hd__xnor2_1 _2802_ (.A(_1206_),
    .B(_1329_),
    .Y(_1330_));
 sky130_fd_sc_hd__and3_1 _2803_ (.A(_0953_),
    .B(_1231_),
    .C(_1232_),
    .X(_1331_));
 sky130_fd_sc_hd__a221oi_1 _2804_ (.A1(_1305_),
    .A2(_1318_),
    .B1(_1330_),
    .B2(_0954_),
    .C1(_1331_),
    .Y(_1332_));
 sky130_fd_sc_hd__o2111a_1 _2805_ (.A1(_0953_),
    .A2(_1330_),
    .B1(_1328_),
    .C1(_1318_),
    .D1(_1305_),
    .X(_1333_));
 sky130_fd_sc_hd__a2bb2o_1 _2806_ (.A1_N(_0990_),
    .A2_N(_1206_),
    .B1(_1252_),
    .B2(_1204_),
    .X(_1334_));
 sky130_fd_sc_hd__a21oi_1 _2807_ (.A1(_1256_),
    .A2(_1330_),
    .B1(_1334_),
    .Y(_1335_));
 sky130_fd_sc_hd__a22o_1 _2808_ (.A1(_1231_),
    .A2(_1232_),
    .B1(_1233_),
    .B2(_1240_),
    .X(_1336_));
 sky130_fd_sc_hd__or3b_1 _2809_ (.A(_1242_),
    .B(_1273_),
    .C_N(_1336_),
    .X(_1337_));
 sky130_fd_sc_hd__o311a_1 _2810_ (.A1(_1250_),
    .A2(_1332_),
    .A3(_1333_),
    .B1(_1335_),
    .C1(_1337_),
    .X(_1338_));
 sky130_fd_sc_hd__nand2_1 _2811_ (.A(_1202_),
    .B(_1338_),
    .Y(_1339_));
 sky130_fd_sc_hd__mux2_1 _2812_ (.A0(_0742_),
    .A1(net1112),
    .S(_1260_),
    .X(_1340_));
 sky130_fd_sc_hd__o211a_1 _2813_ (.A1(_1202_),
    .A2(_1340_),
    .B1(_1339_),
    .C1(net114),
    .X(_1341_));
 sky130_fd_sc_hd__a21o_1 _2814_ (.A1(net144),
    .A2(net937),
    .B1(_1264_),
    .X(_1342_));
 sky130_fd_sc_hd__o221a_1 _2815_ (.A1(net1112),
    .A2(_1263_),
    .B1(_1341_),
    .B2(_1342_),
    .C1(net150),
    .X(_0405_));
 sky130_fd_sc_hd__nand2_1 _2816_ (.A(_1201_),
    .B(_1258_),
    .Y(_1343_));
 sky130_fd_sc_hd__o211a_1 _2817_ (.A1(net1086),
    .A2(_1201_),
    .B1(_1343_),
    .C1(net114),
    .X(_1344_));
 sky130_fd_sc_hd__a211o_1 _2818_ (.A1(net1038),
    .A2(_0988_),
    .B1(_1201_),
    .C1(_0639_),
    .X(_1345_));
 sky130_fd_sc_hd__and2_1 _2819_ (.A(net145),
    .B(_0601_),
    .X(_1346_));
 sky130_fd_sc_hd__o21a_1 _2820_ (.A1(_0638_),
    .A2(_1346_),
    .B1(_0622_),
    .X(_1347_));
 sky130_fd_sc_hd__o21ai_1 _2821_ (.A1(_0582_),
    .A2(_0586_),
    .B1(net145),
    .Y(_1348_));
 sky130_fd_sc_hd__and3_1 _2822_ (.A(_0604_),
    .B(_1347_),
    .C(_1348_),
    .X(_1349_));
 sky130_fd_sc_hd__inv_2 _2823_ (.A(_1349_),
    .Y(_1350_));
 sky130_fd_sc_hd__and2_2 _2824_ (.A(_1345_),
    .B(_1349_),
    .X(_1351_));
 sky130_fd_sc_hd__nand2_2 _2825_ (.A(_1345_),
    .B(_1349_),
    .Y(_1352_));
 sky130_fd_sc_hd__a221o_1 _2826_ (.A1(net1096),
    .A2(_0627_),
    .B1(net104),
    .B2(net799),
    .C1(_1352_),
    .X(_1353_));
 sky130_fd_sc_hd__o221a_1 _2827_ (.A1(net1156),
    .A2(_1351_),
    .B1(_1353_),
    .B2(_1344_),
    .C1(net150),
    .X(_0406_));
 sky130_fd_sc_hd__o211a_1 _2828_ (.A1(net1096),
    .A2(_1201_),
    .B1(_1278_),
    .C1(net114),
    .X(_1354_));
 sky130_fd_sc_hd__a221o_1 _2829_ (.A1(net1101),
    .A2(_0627_),
    .B1(net104),
    .B2(net825),
    .C1(_1352_),
    .X(_1355_));
 sky130_fd_sc_hd__o221a_1 _2830_ (.A1(net1121),
    .A2(_1351_),
    .B1(_1354_),
    .B2(_1355_),
    .C1(net150),
    .X(_0407_));
 sky130_fd_sc_hd__nand2_1 _2831_ (.A(_1201_),
    .B(_1294_),
    .Y(_1356_));
 sky130_fd_sc_hd__o211a_1 _2832_ (.A1(\A[2] ),
    .A2(_1201_),
    .B1(_1356_),
    .C1(net114),
    .X(_1357_));
 sky130_fd_sc_hd__a221o_1 _2833_ (.A1(\A[3] ),
    .A2(_0627_),
    .B1(net104),
    .B2(net505),
    .C1(_1352_),
    .X(_1358_));
 sky130_fd_sc_hd__o221a_1 _2834_ (.A1(net1028),
    .A2(_1351_),
    .B1(_1357_),
    .B2(_1358_),
    .C1(net150),
    .X(_0408_));
 sky130_fd_sc_hd__nand2_1 _2835_ (.A(_1201_),
    .B(_1310_),
    .Y(_1359_));
 sky130_fd_sc_hd__o211a_1 _2836_ (.A1(net1071),
    .A2(_1201_),
    .B1(_1359_),
    .C1(net114),
    .X(_1360_));
 sky130_fd_sc_hd__a221o_1 _2837_ (.A1(net1082),
    .A2(_0627_),
    .B1(net104),
    .B2(net785),
    .C1(_1352_),
    .X(_1361_));
 sky130_fd_sc_hd__o221a_1 _2838_ (.A1(net1128),
    .A2(_1351_),
    .B1(_1360_),
    .B2(_1361_),
    .C1(net150),
    .X(_0409_));
 sky130_fd_sc_hd__nand2_1 _2839_ (.A(_1201_),
    .B(_1324_),
    .Y(_1362_));
 sky130_fd_sc_hd__o211a_1 _2840_ (.A1(\A[4] ),
    .A2(_1201_),
    .B1(_1362_),
    .C1(net114),
    .X(_1363_));
 sky130_fd_sc_hd__a221o_1 _2841_ (.A1(\A[5] ),
    .A2(_0627_),
    .B1(net104),
    .B2(net513),
    .C1(_1352_),
    .X(_1364_));
 sky130_fd_sc_hd__o221a_1 _2842_ (.A1(net1030),
    .A2(_1351_),
    .B1(_1363_),
    .B2(_1364_),
    .C1(net150),
    .X(_0410_));
 sky130_fd_sc_hd__nand2_1 _2843_ (.A(_1201_),
    .B(_1338_),
    .Y(_1365_));
 sky130_fd_sc_hd__o211a_1 _2844_ (.A1(\A[5] ),
    .A2(_1201_),
    .B1(_1365_),
    .C1(net114),
    .X(_1366_));
 sky130_fd_sc_hd__a31o_1 _2845_ (.A1(net1174),
    .A2(_0581_),
    .A3(_0987_),
    .B1(_0599_),
    .X(_1367_));
 sky130_fd_sc_hd__or2_1 _2846_ (.A(net257),
    .B(_0600_),
    .X(_1368_));
 sky130_fd_sc_hd__a31o_1 _2847_ (.A1(net144),
    .A2(_1367_),
    .A3(_1368_),
    .B1(_1352_),
    .X(_1369_));
 sky130_fd_sc_hd__o221a_1 _2848_ (.A1(net1103),
    .A2(_1351_),
    .B1(_1366_),
    .B2(_1369_),
    .C1(net150),
    .X(_0411_));
 sky130_fd_sc_hd__a21oi_1 _2849_ (.A1(_0953_),
    .A2(_1244_),
    .B1(_1333_),
    .Y(_1370_));
 sky130_fd_sc_hd__o21bai_1 _2850_ (.A1(_1242_),
    .A2(_1244_),
    .B1_N(_1273_),
    .Y(_1371_));
 sky130_fd_sc_hd__nor2_1 _2851_ (.A(_1204_),
    .B(_1329_),
    .Y(_1372_));
 sky130_fd_sc_hd__o41a_1 _2852_ (.A1(net1226),
    .A2(_0549_),
    .A3(_1205_),
    .A4(_1372_),
    .B1(_1371_),
    .X(_1373_));
 sky130_fd_sc_hd__o21ai_1 _2853_ (.A1(_1250_),
    .A2(_1370_),
    .B1(_1373_),
    .Y(_1374_));
 sky130_fd_sc_hd__or4bb_1 _2854_ (.A(net1150),
    .B(net102),
    .C_N(_1345_),
    .D_N(_1347_),
    .X(_1375_));
 sky130_fd_sc_hd__o211a_1 _2855_ (.A1(net1086),
    .A2(_0582_),
    .B1(_0587_),
    .C1(_0627_),
    .X(_1376_));
 sky130_fd_sc_hd__a211o_1 _2856_ (.A1(net971),
    .A2(net104),
    .B1(_1375_),
    .C1(_1376_),
    .X(_1377_));
 sky130_fd_sc_hd__a31o_1 _2857_ (.A1(net114),
    .A2(_1201_),
    .A3(_1374_),
    .B1(_1377_),
    .X(_1378_));
 sky130_fd_sc_hd__nand2b_1 _2858_ (.A_N(net1174),
    .B(_1375_),
    .Y(_1379_));
 sky130_fd_sc_hd__and3_1 _2859_ (.A(net150),
    .B(_1378_),
    .C(_1379_),
    .X(_0412_));
 sky130_fd_sc_hd__or3_1 _2860_ (.A(\A[3] ),
    .B(\A[2] ),
    .C(\A[1] ),
    .X(_1380_));
 sky130_fd_sc_hd__or3_1 _2861_ (.A(\A[5] ),
    .B(net1082),
    .C(_1380_),
    .X(_1381_));
 sky130_fd_sc_hd__o221a_1 _2862_ (.A1(_0562_),
    .A2(_0600_),
    .B1(_1367_),
    .B2(_1381_),
    .C1(net144),
    .X(_1382_));
 sky130_fd_sc_hd__and3_1 _2863_ (.A(_1277_),
    .B(_1294_),
    .C(_1310_),
    .X(_1383_));
 sky130_fd_sc_hd__o21a_1 _2864_ (.A1(\A[0] ),
    .A2(_1381_),
    .B1(_0988_),
    .X(_1384_));
 sky130_fd_sc_hd__o21ai_1 _2865_ (.A1(net40),
    .A2(_0988_),
    .B1(net1038),
    .Y(_1385_));
 sky130_fd_sc_hd__o21ai_1 _2866_ (.A1(\insin[4] ),
    .A2(_0579_),
    .B1(net40),
    .Y(_1386_));
 sky130_fd_sc_hd__or3_1 _2867_ (.A(_0848_),
    .B(_0897_),
    .C(_0947_),
    .X(_1387_));
 sky130_fd_sc_hd__or4_1 _2868_ (.A(\insin[4] ),
    .B(_0579_),
    .C(_0692_),
    .D(_0742_),
    .X(_1388_));
 sky130_fd_sc_hd__o31a_1 _2869_ (.A1(_0796_),
    .A2(_1387_),
    .A3(_1388_),
    .B1(_1386_),
    .X(_1389_));
 sky130_fd_sc_hd__o22a_1 _2870_ (.A1(_1384_),
    .A2(_1385_),
    .B1(_1389_),
    .B2(net1038),
    .X(_1390_));
 sky130_fd_sc_hd__nor2_1 _2871_ (.A(_1201_),
    .B(_1390_),
    .Y(_1391_));
 sky130_fd_sc_hd__a41o_1 _2872_ (.A1(_1258_),
    .A2(_1324_),
    .A3(_1338_),
    .A4(_1383_),
    .B1(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__o21ba_1 _2873_ (.A1(net144),
    .A2(_1392_),
    .B1_N(_1382_),
    .X(_1393_));
 sky130_fd_sc_hd__or2_1 _2874_ (.A(net1228),
    .B(_1349_),
    .X(_1394_));
 sky130_fd_sc_hd__o211a_1 _2875_ (.A1(_1350_),
    .A2(_1393_),
    .B1(net1229),
    .C1(net150),
    .X(_0413_));
 sky130_fd_sc_hd__or3_1 _2876_ (.A(net146),
    .B(net114),
    .C(_0601_),
    .X(_1395_));
 sky130_fd_sc_hd__o311a_2 _2877_ (.A1(net146),
    .A2(net114),
    .A3(_0585_),
    .B1(_1395_),
    .C1(_0575_),
    .X(_1396_));
 sky130_fd_sc_hd__or3_2 _2878_ (.A(_0586_),
    .B(_0614_),
    .C(_0620_),
    .X(_1397_));
 sky130_fd_sc_hd__nor2_1 _2879_ (.A(net40),
    .B(\insin[4] ),
    .Y(_1398_));
 sky130_fd_sc_hd__a211o_1 _2880_ (.A1(net1174),
    .A2(\insin[4] ),
    .B1(_0592_),
    .C1(_1398_),
    .X(_1399_));
 sky130_fd_sc_hd__o311a_1 _2881_ (.A1(net40),
    .A2(_0548_),
    .A3(\insin[1] ),
    .B1(_0593_),
    .C1(_0638_),
    .X(_1400_));
 sky130_fd_sc_hd__a21oi_1 _2882_ (.A1(net1175),
    .A2(_1400_),
    .B1(net146),
    .Y(_1401_));
 sky130_fd_sc_hd__a21boi_4 _2883_ (.A1(_1397_),
    .A2(net1176),
    .B1_N(_1396_),
    .Y(_1402_));
 sky130_fd_sc_hd__a22oi_1 _2884_ (.A1(net427),
    .A2(net104),
    .B1(_0796_),
    .B2(net115),
    .Y(_1403_));
 sky130_fd_sc_hd__or3b_4 _2885_ (.A(net1116),
    .B(_0545_),
    .C_N(net979),
    .X(_1404_));
 sky130_fd_sc_hd__inv_2 _2886_ (.A(_1404_),
    .Y(_1405_));
 sky130_fd_sc_hd__o21a_2 _2887_ (.A1(net146),
    .A2(_0627_),
    .B1(_1404_),
    .X(_1406_));
 sky130_fd_sc_hd__o21ai_4 _2888_ (.A1(net146),
    .A2(_0627_),
    .B1(_1404_),
    .Y(_1407_));
 sky130_fd_sc_hd__o221ai_2 _2889_ (.A1(net146),
    .A2(_1403_),
    .B1(_1407_),
    .B2(net1053),
    .C1(_1402_),
    .Y(_1408_));
 sky130_fd_sc_hd__o211a_1 _2890_ (.A1(net1053),
    .A2(_1402_),
    .B1(_1408_),
    .C1(net152),
    .X(_0414_));
 sky130_fd_sc_hd__o2bb2a_1 _2891_ (.A1_N(net217),
    .A2_N(net104),
    .B1(_0847_),
    .B2(net145),
    .X(_1409_));
 sky130_fd_sc_hd__xnor2_1 _2892_ (.A(net1130),
    .B(net1053),
    .Y(_1410_));
 sky130_fd_sc_hd__o221ai_1 _2893_ (.A1(net146),
    .A2(_1409_),
    .B1(_1410_),
    .B2(_1407_),
    .C1(net70),
    .Y(_1411_));
 sky130_fd_sc_hd__o211a_1 _2894_ (.A1(net1130),
    .A2(net70),
    .B1(net1167),
    .C1(net150),
    .X(_0415_));
 sky130_fd_sc_hd__o22a_1 _2895_ (.A1(net773),
    .A2(_0694_),
    .B1(_0897_),
    .B2(net145),
    .X(_1412_));
 sky130_fd_sc_hd__a21oi_1 _2896_ (.A1(\PC[1] ),
    .A2(\PC[0] ),
    .B1(net1026),
    .Y(_1413_));
 sky130_fd_sc_hd__and3_1 _2897_ (.A(net1026),
    .B(\PC[1] ),
    .C(\PC[0] ),
    .X(_1414_));
 sky130_fd_sc_hd__o21ai_1 _2898_ (.A1(_1413_),
    .A2(_1414_),
    .B1(_1406_),
    .Y(_1415_));
 sky130_fd_sc_hd__o21ai_1 _2899_ (.A1(net146),
    .A2(_1412_),
    .B1(_1415_),
    .Y(_1416_));
 sky130_fd_sc_hd__nand2_1 _2900_ (.A(net70),
    .B(_1416_),
    .Y(_1417_));
 sky130_fd_sc_hd__o211a_1 _2901_ (.A1(net1026),
    .A2(net70),
    .B1(_1417_),
    .C1(net152),
    .X(_0416_));
 sky130_fd_sc_hd__a22oi_1 _2902_ (.A1(net749),
    .A2(net104),
    .B1(_0947_),
    .B2(net115),
    .Y(_1418_));
 sky130_fd_sc_hd__and2_1 _2903_ (.A(net1022),
    .B(_1414_),
    .X(_1419_));
 sky130_fd_sc_hd__or2_1 _2904_ (.A(net1022),
    .B(_1414_),
    .X(_1420_));
 sky130_fd_sc_hd__or3b_1 _2905_ (.A(_1407_),
    .B(_1419_),
    .C_N(_1420_),
    .X(_1421_));
 sky130_fd_sc_hd__o211ai_1 _2906_ (.A1(net146),
    .A2(_1418_),
    .B1(_1421_),
    .C1(_1402_),
    .Y(_1422_));
 sky130_fd_sc_hd__o211a_1 _2907_ (.A1(net1022),
    .A2(net70),
    .B1(_1422_),
    .C1(net153),
    .X(_0417_));
 sky130_fd_sc_hd__a22oi_1 _2908_ (.A1(net115),
    .A2(_0692_),
    .B1(net104),
    .B2(net567),
    .Y(_1423_));
 sky130_fd_sc_hd__xnor2_1 _2909_ (.A(net1137),
    .B(_1419_),
    .Y(_1424_));
 sky130_fd_sc_hd__o221ai_1 _2910_ (.A1(net146),
    .A2(_1423_),
    .B1(_1424_),
    .B2(_1407_),
    .C1(_1402_),
    .Y(_1425_));
 sky130_fd_sc_hd__o211a_1 _2911_ (.A1(net1137),
    .A2(_1402_),
    .B1(_1425_),
    .C1(net153),
    .X(_0418_));
 sky130_fd_sc_hd__a22o_1 _2912_ (.A1(net675),
    .A2(net104),
    .B1(_0742_),
    .B2(net115),
    .X(_1426_));
 sky130_fd_sc_hd__a21oi_1 _2913_ (.A1(\PC[4] ),
    .A2(_1419_),
    .B1(net1032),
    .Y(_1427_));
 sky130_fd_sc_hd__and3_1 _2914_ (.A(net1032),
    .B(net1137),
    .C(_1419_),
    .X(_1428_));
 sky130_fd_sc_hd__o31a_1 _2915_ (.A1(_1407_),
    .A2(_1427_),
    .A3(_1428_),
    .B1(net70),
    .X(_1429_));
 sky130_fd_sc_hd__a21bo_1 _2916_ (.A1(_0545_),
    .A2(_1426_),
    .B1_N(_1429_),
    .X(_1430_));
 sky130_fd_sc_hd__o211a_1 _2917_ (.A1(net1032),
    .A2(net70),
    .B1(_1430_),
    .C1(net153),
    .X(_0419_));
 sky130_fd_sc_hd__a22oi_1 _2918_ (.A1(net115),
    .A2(\P[0] ),
    .B1(net377),
    .B2(net104),
    .Y(_1431_));
 sky130_fd_sc_hd__and2_1 _2919_ (.A(net1084),
    .B(_1428_),
    .X(_1432_));
 sky130_fd_sc_hd__o21ai_1 _2920_ (.A1(net1084),
    .A2(_1428_),
    .B1(_1406_),
    .Y(_1433_));
 sky130_fd_sc_hd__o221ai_1 _2921_ (.A1(net146),
    .A2(_1431_),
    .B1(_1432_),
    .B2(_1433_),
    .C1(net70),
    .Y(_1434_));
 sky130_fd_sc_hd__o211a_1 _2922_ (.A1(net1084),
    .A2(_1402_),
    .B1(_1434_),
    .C1(net152),
    .X(_0420_));
 sky130_fd_sc_hd__a22oi_1 _2923_ (.A1(net115),
    .A2(\P[1] ),
    .B1(net475),
    .B2(net104),
    .Y(_1435_));
 sky130_fd_sc_hd__and3_1 _2924_ (.A(net1153),
    .B(net1084),
    .C(_1428_),
    .X(_1436_));
 sky130_fd_sc_hd__o21ai_1 _2925_ (.A1(net1153),
    .A2(_1432_),
    .B1(_1406_),
    .Y(_1437_));
 sky130_fd_sc_hd__o221ai_1 _2926_ (.A1(net1170),
    .A2(_1435_),
    .B1(_1436_),
    .B2(_1437_),
    .C1(net70),
    .Y(_1438_));
 sky130_fd_sc_hd__o211a_1 _2927_ (.A1(net1153),
    .A2(net70),
    .B1(net1171),
    .C1(net152),
    .X(_0421_));
 sky130_fd_sc_hd__a22o_1 _2928_ (.A1(net115),
    .A2(\P[2] ),
    .B1(net491),
    .B2(net104),
    .X(_1439_));
 sky130_fd_sc_hd__and2_1 _2929_ (.A(net1245),
    .B(_1436_),
    .X(_1440_));
 sky130_fd_sc_hd__a32o_1 _2930_ (.A1(_0546_),
    .A2(_1406_),
    .A3(_1436_),
    .B1(_1439_),
    .B2(_0545_),
    .X(_1441_));
 sky130_fd_sc_hd__o21ai_1 _2931_ (.A1(_1407_),
    .A2(_1440_),
    .B1(net70),
    .Y(_1442_));
 sky130_fd_sc_hd__a22o_1 _2932_ (.A1(net70),
    .A2(_1441_),
    .B1(_1442_),
    .B2(net1245),
    .X(_1443_));
 sky130_fd_sc_hd__and2_1 _2933_ (.A(net152),
    .B(net1246),
    .X(_0422_));
 sky130_fd_sc_hd__a22o_1 _2934_ (.A1(net115),
    .A2(net1243),
    .B1(net587),
    .B2(net104),
    .X(_1444_));
 sky130_fd_sc_hd__nand2_1 _2935_ (.A(_1406_),
    .B(_1440_),
    .Y(_1445_));
 sky130_fd_sc_hd__o2bb2a_1 _2936_ (.A1_N(_0545_),
    .A2_N(_1444_),
    .B1(_1445_),
    .B2(net1236),
    .X(_1446_));
 sky130_fd_sc_hd__inv_2 _2937_ (.A(_1446_),
    .Y(_1447_));
 sky130_fd_sc_hd__a22o_1 _2938_ (.A1(net1236),
    .A2(_1442_),
    .B1(_1447_),
    .B2(net70),
    .X(_1448_));
 sky130_fd_sc_hd__and2_1 _2939_ (.A(net152),
    .B(net1244),
    .X(_0423_));
 sky130_fd_sc_hd__a22o_1 _2940_ (.A1(net115),
    .A2(net1241),
    .B1(net625),
    .B2(net104),
    .X(_1449_));
 sky130_fd_sc_hd__and3_1 _2941_ (.A(net1236),
    .B(net1263),
    .C(_1436_),
    .X(_1450_));
 sky130_fd_sc_hd__a21oi_1 _2942_ (.A1(net1066),
    .A2(_1450_),
    .B1(_1407_),
    .Y(_1451_));
 sky130_fd_sc_hd__a22o_1 _2943_ (.A1(_0545_),
    .A2(_1449_),
    .B1(net1237),
    .B2(_1451_),
    .X(_1452_));
 sky130_fd_sc_hd__nand2b_1 _2944_ (.A_N(_1451_),
    .B(net70),
    .Y(_1453_));
 sky130_fd_sc_hd__a22o_1 _2945_ (.A1(net70),
    .A2(_1452_),
    .B1(_1453_),
    .B2(net1066),
    .X(_1454_));
 sky130_fd_sc_hd__and2_1 _2946_ (.A(net152),
    .B(_1454_),
    .X(_0424_));
 sky130_fd_sc_hd__a22o_1 _2947_ (.A1(net115),
    .A2(net1186),
    .B1(net527),
    .B2(_0693_),
    .X(_1455_));
 sky130_fd_sc_hd__nor2_1 _2948_ (.A(net1198),
    .B(_1407_),
    .Y(_1456_));
 sky130_fd_sc_hd__a32o_1 _2949_ (.A1(net1066),
    .A2(net1237),
    .A3(_1456_),
    .B1(_1455_),
    .B2(_0545_),
    .X(_1457_));
 sky130_fd_sc_hd__a22o_1 _2950_ (.A1(net1198),
    .A2(_1453_),
    .B1(_1457_),
    .B2(net70),
    .X(_1458_));
 sky130_fd_sc_hd__and2_1 _2951_ (.A(net152),
    .B(_1458_),
    .X(_0425_));
 sky130_fd_sc_hd__o21ai_1 _2952_ (.A1(_0576_),
    .A2(_1395_),
    .B1(net1038),
    .Y(_1459_));
 sky130_fd_sc_hd__o31a_1 _2953_ (.A1(net1038),
    .A2(_0576_),
    .A3(_1395_),
    .B1(net149),
    .X(_1460_));
 sky130_fd_sc_hd__nand2_1 _2954_ (.A(net1039),
    .B(_1460_),
    .Y(_0426_));
 sky130_fd_sc_hd__or2_2 _2955_ (.A(_0747_),
    .B(_1175_),
    .X(_1461_));
 sky130_fd_sc_hd__mux2_1 _2956_ (.A0(net13),
    .A1(net601),
    .S(_1461_),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_1 _2957_ (.A0(net14),
    .A1(net795),
    .S(_1461_),
    .X(_0428_));
 sky130_fd_sc_hd__mux2_1 _2958_ (.A0(net15),
    .A1(net993),
    .S(_1461_),
    .X(_0429_));
 sky130_fd_sc_hd__mux2_1 _2959_ (.A0(net16),
    .A1(net1005),
    .S(_1461_),
    .X(_0430_));
 sky130_fd_sc_hd__nand2_1 _2960_ (.A(_0575_),
    .B(_1405_),
    .Y(_1462_));
 sky130_fd_sc_hd__nor2_1 _2961_ (.A(net148),
    .B(_1462_),
    .Y(_1463_));
 sky130_fd_sc_hd__mux2_1 _2962_ (.A0(net427),
    .A1(net1253),
    .S(net98),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _2963_ (.A0(net217),
    .A1(net1261),
    .S(net97),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_1 _2964_ (.A0(net773),
    .A1(net1252),
    .S(net98),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_1 _2965_ (.A0(net749),
    .A1(net1258),
    .S(net97),
    .X(_0434_));
 sky130_fd_sc_hd__mux2_1 _2966_ (.A0(net567),
    .A1(net1262),
    .S(net98),
    .X(_0435_));
 sky130_fd_sc_hd__mux2_1 _2967_ (.A0(net675),
    .A1(net1257),
    .S(net97),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _2968_ (.A0(net377),
    .A1(net1260),
    .S(net97),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _2969_ (.A0(net475),
    .A1(net30),
    .S(net97),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _2970_ (.A0(net491),
    .A1(net31),
    .S(net97),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_1 _2971_ (.A0(net587),
    .A1(net32),
    .S(net97),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _2972_ (.A0(net625),
    .A1(net33),
    .S(net97),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _2973_ (.A0(net527),
    .A1(net34),
    .S(net97),
    .X(_0442_));
 sky130_fd_sc_hd__mux2_1 _2974_ (.A0(net971),
    .A1(net51),
    .S(net99),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_1 _2975_ (.A0(net997),
    .A1(net40),
    .S(net99),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_1 _2976_ (.A0(net585),
    .A1(\A[0] ),
    .S(net99),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _2977_ (.A0(net761),
    .A1(\A[1] ),
    .S(net99),
    .X(_0446_));
 sky130_fd_sc_hd__mux2_1 _2978_ (.A0(net885),
    .A1(\A[2] ),
    .S(net99),
    .X(_0447_));
 sky130_fd_sc_hd__mux2_1 _2979_ (.A0(net747),
    .A1(net1264),
    .S(net99),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _2980_ (.A0(net743),
    .A1(\A[4] ),
    .S(net99),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _2981_ (.A0(net937),
    .A1(\A[5] ),
    .S(net99),
    .X(_0450_));
 sky130_fd_sc_hd__mux2_1 _2982_ (.A0(net799),
    .A1(net1251),
    .S(net99),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _2983_ (.A0(net825),
    .A1(net1250),
    .S(net99),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _2984_ (.A0(net505),
    .A1(net1259),
    .S(net99),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _2985_ (.A0(net785),
    .A1(net1254),
    .S(net99),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_1 _2986_ (.A0(net513),
    .A1(net1256),
    .S(net99),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _2987_ (.A0(net257),
    .A1(net1255),
    .S(net99),
    .X(_0456_));
 sky130_fd_sc_hd__mux2_1 _2988_ (.A0(net697),
    .A1(net134),
    .S(net98),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _2989_ (.A0(net667),
    .A1(net126),
    .S(net98),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _2990_ (.A0(net767),
    .A1(net123),
    .S(net98),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _2991_ (.A0(net613),
    .A1(net119),
    .S(net98),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _2992_ (.A0(net595),
    .A1(net118),
    .S(net98),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _2993_ (.A0(net651),
    .A1(net116),
    .S(net97),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _2994_ (.A0(net417),
    .A1(net1247),
    .S(net97),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _2995_ (.A0(net983),
    .A1(\P[1] ),
    .S(net97),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _2996_ (.A0(net563),
    .A1(net1248),
    .S(net97),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _2997_ (.A0(net463),
    .A1(net1243),
    .S(net97),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _2998_ (.A0(net945),
    .A1(net1241),
    .S(net97),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _2999_ (.A0(net553),
    .A1(net1186),
    .S(net97),
    .X(_0468_));
 sky130_fd_sc_hd__and2b_1 _3000_ (.A_N(last_inter),
    .B(net12),
    .X(_1464_));
 sky130_fd_sc_hd__o211a_1 _3001_ (.A1(net979),
    .A2(_1464_),
    .B1(_1462_),
    .C1(net153),
    .X(_0469_));
 sky130_fd_sc_hd__o21ai_1 _3002_ (.A1(net102),
    .A2(_0694_),
    .B1(net1116),
    .Y(_1465_));
 sky130_fd_sc_hd__a21oi_1 _3003_ (.A1(_1462_),
    .A2(net1117),
    .B1(net148),
    .Y(_0470_));
 sky130_fd_sc_hd__nand2_1 _3004_ (.A(spi_clkdiv),
    .B(net106),
    .Y(_1466_));
 sky130_fd_sc_hd__nand2_2 _3005_ (.A(net1007),
    .B(net1164),
    .Y(_1467_));
 sky130_fd_sc_hd__nor2_1 _3006_ (.A(_1117_),
    .B(_1467_),
    .Y(_1468_));
 sky130_fd_sc_hd__or2_1 _3007_ (.A(_1117_),
    .B(_1467_),
    .X(_1469_));
 sky130_fd_sc_hd__nand2_1 _3008_ (.A(_0544_),
    .B(net1123),
    .Y(_1470_));
 sky130_fd_sc_hd__o21a_1 _3009_ (.A1(_0567_),
    .A2(_1470_),
    .B1(_1469_),
    .X(_1471_));
 sky130_fd_sc_hd__nor2_1 _3010_ (.A(_0569_),
    .B(_1471_),
    .Y(_1472_));
 sky130_fd_sc_hd__nand2b_2 _3011_ (.A_N(\startup_cycle[0] ),
    .B(net1007),
    .Y(_1473_));
 sky130_fd_sc_hd__or3_1 _3012_ (.A(_0544_),
    .B(\startup_cycle[2] ),
    .C(_1473_),
    .X(_1474_));
 sky130_fd_sc_hd__a21oi_1 _3013_ (.A1(_1471_),
    .A2(_1474_),
    .B1(_0569_),
    .Y(_1475_));
 sky130_fd_sc_hd__or3_1 _3014_ (.A(_0544_),
    .B(\startup_cycle[2] ),
    .C(_1467_),
    .X(_1476_));
 sky130_fd_sc_hd__o21a_1 _3015_ (.A1(_0567_),
    .A2(_1117_),
    .B1(_1476_),
    .X(_1477_));
 sky130_fd_sc_hd__o21ba_1 _3016_ (.A1(_0569_),
    .A2(_1477_),
    .B1_N(_1475_),
    .X(_1478_));
 sky130_fd_sc_hd__o31a_1 _3017_ (.A1(_0569_),
    .A2(_1467_),
    .A3(_1470_),
    .B1(_1478_),
    .X(_1479_));
 sky130_fd_sc_hd__or3b_1 _3018_ (.A(_0569_),
    .B(net1007),
    .C_N(\startup_cycle[0] ),
    .X(_1480_));
 sky130_fd_sc_hd__o21ai_1 _3019_ (.A1(_0566_),
    .A2(_1480_),
    .B1(_1479_),
    .Y(_1481_));
 sky130_fd_sc_hd__nor2_1 _3020_ (.A(net106),
    .B(_0570_),
    .Y(_1482_));
 sky130_fd_sc_hd__or2_2 _3021_ (.A(net1009),
    .B(net108),
    .X(_1483_));
 sky130_fd_sc_hd__o21a_1 _3022_ (.A1(net106),
    .A2(_1481_),
    .B1(_1483_),
    .X(_1484_));
 sky130_fd_sc_hd__or2_1 _3023_ (.A(net1238),
    .B(_1484_),
    .X(_1485_));
 sky130_fd_sc_hd__nand2_1 _3024_ (.A(net1238),
    .B(_1483_),
    .Y(_1486_));
 sky130_fd_sc_hd__and3_1 _3025_ (.A(net155),
    .B(_1485_),
    .C(_1486_),
    .X(_0471_));
 sky130_fd_sc_hd__or4b_1 _3026_ (.A(net1231),
    .B(_0563_),
    .C(_1486_),
    .D_N(net1224),
    .X(_1487_));
 sky130_fd_sc_hd__xnor2_1 _3027_ (.A(net1231),
    .B(_1486_),
    .Y(_1488_));
 sky130_fd_sc_hd__and3_1 _3028_ (.A(net155),
    .B(_1487_),
    .C(net1232),
    .X(_0472_));
 sky130_fd_sc_hd__a31o_1 _3029_ (.A1(\ROM_spi_cycle[1] ),
    .A2(\ROM_spi_cycle[0] ),
    .A3(_1483_),
    .B1(net1098),
    .X(_1489_));
 sky130_fd_sc_hd__and4_1 _3030_ (.A(net1098),
    .B(\ROM_spi_cycle[1] ),
    .C(\ROM_spi_cycle[0] ),
    .D(_1483_),
    .X(_1490_));
 sky130_fd_sc_hd__and3b_1 _3031_ (.A_N(_1490_),
    .B(net155),
    .C(net1099),
    .X(_0473_));
 sky130_fd_sc_hd__or2_1 _3032_ (.A(net1107),
    .B(_1490_),
    .X(_1491_));
 sky130_fd_sc_hd__nand2_1 _3033_ (.A(net1107),
    .B(_1490_),
    .Y(_1492_));
 sky130_fd_sc_hd__and3_1 _3034_ (.A(net155),
    .B(_1491_),
    .C(net1108),
    .X(_0474_));
 sky130_fd_sc_hd__xnor2_1 _3035_ (.A(net1224),
    .B(net1108),
    .Y(_1493_));
 sky130_fd_sc_hd__and3_1 _3036_ (.A(net155),
    .B(_1487_),
    .C(_1493_),
    .X(_0475_));
 sky130_fd_sc_hd__or4_1 _3037_ (.A(_0542_),
    .B(_0543_),
    .C(_0566_),
    .D(_1473_),
    .X(_1494_));
 sky130_fd_sc_hd__nor2_1 _3038_ (.A(\startup_cycle[5] ),
    .B(_1494_),
    .Y(_1495_));
 sky130_fd_sc_hd__o21a_1 _3039_ (.A1(net1164),
    .A2(_1495_),
    .B1(_1482_),
    .X(_1496_));
 sky130_fd_sc_hd__nor2_1 _3040_ (.A(net1164),
    .B(_1482_),
    .Y(_1497_));
 sky130_fd_sc_hd__o21ai_1 _3041_ (.A1(_1496_),
    .A2(_1497_),
    .B1(net154),
    .Y(_0476_));
 sky130_fd_sc_hd__o21ai_1 _3042_ (.A1(net1007),
    .A2(_1496_),
    .B1(net154),
    .Y(_1498_));
 sky130_fd_sc_hd__a21oi_1 _3043_ (.A1(net1007),
    .A2(_1496_),
    .B1(_1498_),
    .Y(_0477_));
 sky130_fd_sc_hd__o21ai_1 _3044_ (.A1(net106),
    .A2(_1467_),
    .B1(net1123),
    .Y(_1499_));
 sky130_fd_sc_hd__or4_1 _3045_ (.A(net1123),
    .B(net106),
    .C(_0570_),
    .D(_1467_),
    .X(_1500_));
 sky130_fd_sc_hd__a21oi_1 _3046_ (.A1(net1124),
    .A2(_1500_),
    .B1(net147),
    .Y(_0478_));
 sky130_fd_sc_hd__a31o_1 _3047_ (.A1(net1007),
    .A2(net1164),
    .A3(net108),
    .B1(_1470_),
    .X(_1501_));
 sky130_fd_sc_hd__and3_1 _3048_ (.A(net108),
    .B(_0571_),
    .C(_1468_),
    .X(_1502_));
 sky130_fd_sc_hd__o2111a_1 _3049_ (.A1(net107),
    .A2(_1469_),
    .B1(_1501_),
    .C1(_0566_),
    .D1(net154),
    .X(_0479_));
 sky130_fd_sc_hd__a221o_1 _3050_ (.A1(_1482_),
    .A2(_1495_),
    .B1(_1502_),
    .B2(net1088),
    .C1(net147),
    .X(_1503_));
 sky130_fd_sc_hd__o21ba_1 _3051_ (.A1(net1088),
    .A2(_1502_),
    .B1_N(_1503_),
    .X(_0480_));
 sky130_fd_sc_hd__a21o_1 _3052_ (.A1(net1088),
    .A2(_1502_),
    .B1(net1208),
    .X(_1504_));
 sky130_fd_sc_hd__and3_1 _3053_ (.A(net1208),
    .B(net1088),
    .C(_1468_),
    .X(_1505_));
 sky130_fd_sc_hd__nand2_1 _3054_ (.A(_1482_),
    .B(_1505_),
    .Y(_1506_));
 sky130_fd_sc_hd__and3_1 _3055_ (.A(net154),
    .B(net1209),
    .C(_1506_),
    .X(_0481_));
 sky130_fd_sc_hd__o311a_1 _3056_ (.A1(_0570_),
    .A2(_1495_),
    .A3(_1505_),
    .B1(net108),
    .C1(net1090),
    .X(_1507_));
 sky130_fd_sc_hd__a211oi_1 _3057_ (.A1(_0542_),
    .A2(_1506_),
    .B1(_1507_),
    .C1(net147),
    .Y(_0482_));
 sky130_fd_sc_hd__and2_1 _3058_ (.A(net156),
    .B(net12),
    .X(_0483_));
 sky130_fd_sc_hd__or4b_2 _3059_ (.A(net1182),
    .B(net1178),
    .C(\mem_cycle[2] ),
    .D_N(net1188),
    .X(_1508_));
 sky130_fd_sc_hd__nor2_1 _3060_ (.A(\mem_cycle[4] ),
    .B(_1508_),
    .Y(_1509_));
 sky130_fd_sc_hd__o21ba_1 _3061_ (.A1(_1044_),
    .A2(_1509_),
    .B1_N(_1057_),
    .X(_1510_));
 sky130_fd_sc_hd__o21a_1 _3062_ (.A1(_1049_),
    .A2(_1510_),
    .B1(_1105_),
    .X(_1511_));
 sky130_fd_sc_hd__or3b_1 _3063_ (.A(_1470_),
    .B(net1007),
    .C_N(\startup_cycle[0] ),
    .X(_1512_));
 sky130_fd_sc_hd__o21a_1 _3064_ (.A1(_0566_),
    .A2(_1473_),
    .B1(_1115_),
    .X(_1513_));
 sky130_fd_sc_hd__or3_1 _3065_ (.A(_0542_),
    .B(\startup_cycle[5] ),
    .C(\startup_cycle[4] ),
    .X(_1514_));
 sky130_fd_sc_hd__o21a_1 _3066_ (.A1(_1473_),
    .A2(_1514_),
    .B1(_1480_),
    .X(_1515_));
 sky130_fd_sc_hd__a31o_1 _3067_ (.A1(_0568_),
    .A2(_1512_),
    .A3(_1513_),
    .B1(_0569_),
    .X(_1516_));
 sky130_fd_sc_hd__o21ai_1 _3068_ (.A1(_1117_),
    .A2(_1515_),
    .B1(_1516_),
    .Y(_1517_));
 sky130_fd_sc_hd__o21ai_1 _3069_ (.A1(_1481_),
    .A2(_1517_),
    .B1(_1511_),
    .Y(_1518_));
 sky130_fd_sc_hd__o31a_1 _3070_ (.A1(\mem_cycle[4] ),
    .A2(_0571_),
    .A3(_1508_),
    .B1(_1517_),
    .X(_1519_));
 sky130_fd_sc_hd__a221o_1 _3071_ (.A1(net1024),
    .A2(_1518_),
    .B1(_1519_),
    .B2(_1511_),
    .C1(net147),
    .X(_0484_));
 sky130_fd_sc_hd__o21ai_1 _3072_ (.A1(net1182),
    .A2(_0572_),
    .B1(_1068_),
    .Y(_1520_));
 sky130_fd_sc_hd__o21ai_1 _3073_ (.A1(_1057_),
    .A2(_1520_),
    .B1(_0969_),
    .Y(_1521_));
 sky130_fd_sc_hd__or4b_1 _3074_ (.A(\startup_cycle[6] ),
    .B(\startup_cycle[5] ),
    .C(_0543_),
    .D_N(_0566_),
    .X(_1522_));
 sky130_fd_sc_hd__and3_1 _3075_ (.A(_1114_),
    .B(_1514_),
    .C(_1522_),
    .X(_1523_));
 sky130_fd_sc_hd__o21ai_1 _3076_ (.A1(_0567_),
    .A2(_1523_),
    .B1(_0571_),
    .Y(_1524_));
 sky130_fd_sc_hd__or3b_1 _3077_ (.A(\startup_cycle[5] ),
    .B(\startup_cycle[4] ),
    .C_N(_1117_),
    .X(_1525_));
 sky130_fd_sc_hd__a21oi_1 _3078_ (.A1(net1090),
    .A2(_1525_),
    .B1(_1473_),
    .Y(_1526_));
 sky130_fd_sc_hd__a211o_1 _3079_ (.A1(_0569_),
    .A2(_1526_),
    .B1(_1524_),
    .C1(net107),
    .X(_1527_));
 sky130_fd_sc_hd__and3_1 _3080_ (.A(_1483_),
    .B(_1521_),
    .C(_1527_),
    .X(_1528_));
 sky130_fd_sc_hd__nor2_2 _3081_ (.A(\mem_cycle[1] ),
    .B(_0572_),
    .Y(_1529_));
 sky130_fd_sc_hd__a2111o_1 _3082_ (.A1(net1195),
    .A2(_0746_),
    .B1(_1529_),
    .C1(_0553_),
    .D1(_0571_),
    .X(_1530_));
 sky130_fd_sc_hd__a21o_1 _3083_ (.A1(_1524_),
    .A2(_1530_),
    .B1(net107),
    .X(_1531_));
 sky130_fd_sc_hd__o21ai_1 _3084_ (.A1(\ROM_spi_cycle[0] ),
    .A2(net108),
    .B1(_1531_),
    .Y(_1532_));
 sky130_fd_sc_hd__mux2_1 _3085_ (.A0(net1203),
    .A1(_1532_),
    .S(_1528_),
    .X(_1533_));
 sky130_fd_sc_hd__and2_1 _3086_ (.A(net155),
    .B(net1204),
    .X(_0485_));
 sky130_fd_sc_hd__o221a_1 _3087_ (.A1(\ROM_spi_cycle[0] ),
    .A2(net108),
    .B1(_0970_),
    .B2(_1111_),
    .C1(_1483_),
    .X(_1534_));
 sky130_fd_sc_hd__o31a_1 _3088_ (.A1(net107),
    .A2(_0570_),
    .A3(_1119_),
    .B1(_1534_),
    .X(_1535_));
 sky130_fd_sc_hd__or3b_1 _3089_ (.A(_1109_),
    .B(_1123_),
    .C_N(\ROM_addr_buff[8] ),
    .X(_1536_));
 sky130_fd_sc_hd__a22oi_1 _3090_ (.A1(net1105),
    .A2(_1121_),
    .B1(_1123_),
    .B2(net1076),
    .Y(_1537_));
 sky130_fd_sc_hd__a31o_1 _3091_ (.A1(_1107_),
    .A2(_1536_),
    .A3(_1537_),
    .B1(_0571_),
    .X(_1538_));
 sky130_fd_sc_hd__nor2_1 _3092_ (.A(net991),
    .B(net108),
    .Y(_1539_));
 sky130_fd_sc_hd__a31o_1 _3093_ (.A1(net109),
    .A2(_1118_),
    .A3(_1538_),
    .B1(_1539_),
    .X(_1540_));
 sky130_fd_sc_hd__mux2_1 _3094_ (.A0(_0541_),
    .A1(_1540_),
    .S(_1535_),
    .X(_1541_));
 sky130_fd_sc_hd__nor2_1 _3095_ (.A(net147),
    .B(net1148),
    .Y(_0486_));
 sky130_fd_sc_hd__and3_1 _3096_ (.A(_0570_),
    .B(_0574_),
    .C(_1508_),
    .X(_1542_));
 sky130_fd_sc_hd__or3_1 _3097_ (.A(_0543_),
    .B(_0568_),
    .C(_1114_),
    .X(_1543_));
 sky130_fd_sc_hd__a211o_1 _3098_ (.A1(_1113_),
    .A2(_1543_),
    .B1(_1542_),
    .C1(_1106_),
    .X(_1544_));
 sky130_fd_sc_hd__o31a_1 _3099_ (.A1(_0552_),
    .A2(_0571_),
    .A3(_1508_),
    .B1(_1543_),
    .X(_1545_));
 sky130_fd_sc_hd__mux2_1 _3100_ (.A0(_1545_),
    .A1(_0540_),
    .S(_1544_),
    .X(_1546_));
 sky130_fd_sc_hd__nand2_1 _3101_ (.A(net152),
    .B(net1192),
    .Y(_0487_));
 sky130_fd_sc_hd__o21ai_1 _3102_ (.A1(net106),
    .A2(_1112_),
    .B1(net985),
    .Y(_1547_));
 sky130_fd_sc_hd__nand2_1 _3103_ (.A(net152),
    .B(net986),
    .Y(_0488_));
 sky130_fd_sc_hd__o21a_2 _3104_ (.A1(\ROM_spi_cycle[0] ),
    .A2(_1466_),
    .B1(_1484_),
    .X(_1548_));
 sky130_fd_sc_hd__o21ai_4 _3105_ (.A1(\ROM_spi_cycle[0] ),
    .A2(_1466_),
    .B1(_1484_),
    .Y(_1549_));
 sky130_fd_sc_hd__o211a_1 _3106_ (.A1(_1475_),
    .A2(_1479_),
    .B1(_1548_),
    .C1(net108),
    .X(_1550_));
 sky130_fd_sc_hd__a21oi_1 _3107_ (.A1(net963),
    .A2(_1549_),
    .B1(_1550_),
    .Y(_1551_));
 sky130_fd_sc_hd__nor2_1 _3108_ (.A(net147),
    .B(net964),
    .Y(_0489_));
 sky130_fd_sc_hd__mux2_1 _3109_ (.A0(net963),
    .A1(_1473_),
    .S(net108),
    .X(_1552_));
 sky130_fd_sc_hd__or2_1 _3110_ (.A(_1549_),
    .B(_1552_),
    .X(_1553_));
 sky130_fd_sc_hd__o211a_1 _3111_ (.A1(net981),
    .A2(_1548_),
    .B1(_1553_),
    .C1(net154),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _3112_ (.A0(net981),
    .A1(_1478_),
    .S(net108),
    .X(_1554_));
 sky130_fd_sc_hd__or2_1 _3113_ (.A(_1549_),
    .B(_1554_),
    .X(_1555_));
 sky130_fd_sc_hd__o211a_1 _3114_ (.A1(net1003),
    .A2(_1548_),
    .B1(_1555_),
    .C1(net154),
    .X(_0491_));
 sky130_fd_sc_hd__o21a_1 _3115_ (.A1(_1472_),
    .A2(_1479_),
    .B1(net108),
    .X(_1556_));
 sky130_fd_sc_hd__a211o_1 _3116_ (.A1(\ROM_spi_dat_out[2] ),
    .A2(net107),
    .B1(_1549_),
    .C1(_1556_),
    .X(_1557_));
 sky130_fd_sc_hd__o211a_1 _3117_ (.A1(net995),
    .A2(_1548_),
    .B1(_1557_),
    .C1(net154),
    .X(_0492_));
 sky130_fd_sc_hd__or2_1 _3118_ (.A(net107),
    .B(_1479_),
    .X(_1558_));
 sky130_fd_sc_hd__o21ai_1 _3119_ (.A1(net995),
    .A2(net108),
    .B1(_1558_),
    .Y(_1559_));
 sky130_fd_sc_hd__nand2_1 _3120_ (.A(_1548_),
    .B(_1559_),
    .Y(_1560_));
 sky130_fd_sc_hd__o211a_1 _3121_ (.A1(net999),
    .A2(_1548_),
    .B1(_1560_),
    .C1(net154),
    .X(_0493_));
 sky130_fd_sc_hd__a211o_1 _3122_ (.A1(\ROM_spi_dat_out[4] ),
    .A2(net107),
    .B1(_1549_),
    .C1(_1556_),
    .X(_1561_));
 sky130_fd_sc_hd__o211a_1 _3123_ (.A1(net987),
    .A2(_1548_),
    .B1(_1561_),
    .C1(net154),
    .X(_0494_));
 sky130_fd_sc_hd__nor2_1 _3124_ (.A(_0569_),
    .B(_1469_),
    .Y(_1562_));
 sky130_fd_sc_hd__o22a_1 _3125_ (.A1(net987),
    .A2(net108),
    .B1(_1558_),
    .B2(_1562_),
    .X(_1563_));
 sky130_fd_sc_hd__or2_1 _3126_ (.A(_1549_),
    .B(_1563_),
    .X(_1564_));
 sky130_fd_sc_hd__o211a_1 _3127_ (.A1(net989),
    .A2(_1548_),
    .B1(_1564_),
    .C1(net154),
    .X(_0495_));
 sky130_fd_sc_hd__a211o_1 _3128_ (.A1(net989),
    .A2(net107),
    .B1(_1549_),
    .C1(_1556_),
    .X(_1565_));
 sky130_fd_sc_hd__o211a_1 _3129_ (.A1(net991),
    .A2(_1548_),
    .B1(_1565_),
    .C1(net154),
    .X(_0496_));
 sky130_fd_sc_hd__nor2_2 _3130_ (.A(_0599_),
    .B(_1397_),
    .Y(_1566_));
 sky130_fd_sc_hd__o21a_4 _3131_ (.A1(net1170),
    .A2(_1566_),
    .B1(_1396_),
    .X(_1567_));
 sky130_fd_sc_hd__o21ai_4 _3132_ (.A1(net1170),
    .A2(_1566_),
    .B1(_1396_),
    .Y(_1568_));
 sky130_fd_sc_hd__a21o_1 _3133_ (.A1(net1053),
    .A2(_1404_),
    .B1(_1568_),
    .X(_1569_));
 sky130_fd_sc_hd__o211a_1 _3134_ (.A1(net1076),
    .A2(_1567_),
    .B1(_1569_),
    .C1(net153),
    .X(_0497_));
 sky130_fd_sc_hd__a21o_1 _3135_ (.A1(net1130),
    .A2(_1404_),
    .B1(_1568_),
    .X(_1570_));
 sky130_fd_sc_hd__o211a_1 _3136_ (.A1(net1114),
    .A2(_1567_),
    .B1(net1131),
    .C1(net153),
    .X(_0498_));
 sky130_fd_sc_hd__or3_1 _3137_ (.A(net1026),
    .B(_1405_),
    .C(_1568_),
    .X(_1571_));
 sky130_fd_sc_hd__o211a_1 _3138_ (.A1(net1135),
    .A2(_1567_),
    .B1(_1571_),
    .C1(net153),
    .X(_0499_));
 sky130_fd_sc_hd__a21o_1 _3139_ (.A1(net1022),
    .A2(_1404_),
    .B1(_1568_),
    .X(_1572_));
 sky130_fd_sc_hd__o211a_1 _3140_ (.A1(net1144),
    .A2(_1567_),
    .B1(_1572_),
    .C1(net153),
    .X(_0500_));
 sky130_fd_sc_hd__a21o_1 _3141_ (.A1(net1137),
    .A2(_1404_),
    .B1(_1568_),
    .X(_1573_));
 sky130_fd_sc_hd__o211a_1 _3142_ (.A1(net1105),
    .A2(_1567_),
    .B1(net1138),
    .C1(net153),
    .X(_0501_));
 sky130_fd_sc_hd__a21o_1 _3143_ (.A1(net1032),
    .A2(_1404_),
    .B1(_1568_),
    .X(_1574_));
 sky130_fd_sc_hd__o211a_1 _3144_ (.A1(net1036),
    .A2(_1567_),
    .B1(_1574_),
    .C1(net153),
    .X(_0502_));
 sky130_fd_sc_hd__a21o_1 _3145_ (.A1(net1084),
    .A2(_1404_),
    .B1(_1568_),
    .X(_1575_));
 sky130_fd_sc_hd__o211a_1 _3146_ (.A1(net1092),
    .A2(_1567_),
    .B1(_1575_),
    .C1(net153),
    .X(_0503_));
 sky130_fd_sc_hd__a21o_1 _3147_ (.A1(net1153),
    .A2(_1404_),
    .B1(_1568_),
    .X(_1576_));
 sky130_fd_sc_hd__o211a_1 _3148_ (.A1(net1074),
    .A2(_1567_),
    .B1(net1154),
    .C1(net152),
    .X(_0504_));
 sky130_fd_sc_hd__a21o_1 _3149_ (.A1(net31),
    .A2(_1404_),
    .B1(_1568_),
    .X(_1577_));
 sky130_fd_sc_hd__o211a_1 _3150_ (.A1(net1180),
    .A2(_1567_),
    .B1(_1577_),
    .C1(net152),
    .X(_0505_));
 sky130_fd_sc_hd__a21o_1 _3151_ (.A1(net32),
    .A2(_1404_),
    .B1(_1568_),
    .X(_1578_));
 sky130_fd_sc_hd__o211a_1 _3152_ (.A1(net1193),
    .A2(_1567_),
    .B1(_1578_),
    .C1(net152),
    .X(_0506_));
 sky130_fd_sc_hd__a21o_1 _3153_ (.A1(net1066),
    .A2(_1404_),
    .B1(_1568_),
    .X(_1579_));
 sky130_fd_sc_hd__o211a_1 _3154_ (.A1(net1016),
    .A2(_1567_),
    .B1(net1067),
    .C1(net152),
    .X(_0507_));
 sky130_fd_sc_hd__a21o_1 _3155_ (.A1(net1198),
    .A2(_1404_),
    .B1(_1568_),
    .X(_1580_));
 sky130_fd_sc_hd__o211a_1 _3156_ (.A1(net1126),
    .A2(_1567_),
    .B1(_1580_),
    .C1(net152),
    .X(_0508_));
 sky130_fd_sc_hd__and3_4 _3157_ (.A(\mem_cycle[0] ),
    .B(_0969_),
    .C(_1529_),
    .X(_1581_));
 sky130_fd_sc_hd__nand2_4 _3158_ (.A(_1059_),
    .B(_1529_),
    .Y(_1582_));
 sky130_fd_sc_hd__or2_1 _3159_ (.A(net1141),
    .B(_1581_),
    .X(_1583_));
 sky130_fd_sc_hd__o211a_1 _3160_ (.A1(net1076),
    .A2(_1582_),
    .B1(net1142),
    .C1(net155),
    .X(_0509_));
 sky130_fd_sc_hd__or2_1 _3161_ (.A(\last_addr[1] ),
    .B(_1581_),
    .X(_1584_));
 sky130_fd_sc_hd__o211a_1 _3162_ (.A1(net1114),
    .A2(_1582_),
    .B1(_1584_),
    .C1(net153),
    .X(_0510_));
 sky130_fd_sc_hd__or2_1 _3163_ (.A(net1055),
    .B(_1581_),
    .X(_1585_));
 sky130_fd_sc_hd__o211a_1 _3164_ (.A1(\ROM_addr_buff[2] ),
    .A2(_1582_),
    .B1(net1056),
    .C1(net153),
    .X(_0511_));
 sky130_fd_sc_hd__or2_1 _3165_ (.A(net1041),
    .B(_1581_),
    .X(_1586_));
 sky130_fd_sc_hd__o211a_1 _3166_ (.A1(\ROM_addr_buff[3] ),
    .A2(_1582_),
    .B1(net1042),
    .C1(net153),
    .X(_0512_));
 sky130_fd_sc_hd__or2_1 _3167_ (.A(\last_addr[4] ),
    .B(_1581_),
    .X(_1587_));
 sky130_fd_sc_hd__o211a_1 _3168_ (.A1(net1105),
    .A2(_1582_),
    .B1(_1587_),
    .C1(net157),
    .X(_0513_));
 sky130_fd_sc_hd__or2_1 _3169_ (.A(net1047),
    .B(_1581_),
    .X(_1588_));
 sky130_fd_sc_hd__o211a_1 _3170_ (.A1(net1036),
    .A2(_1582_),
    .B1(net1048),
    .C1(net157),
    .X(_0514_));
 sky130_fd_sc_hd__or2_1 _3171_ (.A(net1050),
    .B(_1581_),
    .X(_1589_));
 sky130_fd_sc_hd__o211a_1 _3172_ (.A1(\ROM_addr_buff[6] ),
    .A2(_1582_),
    .B1(net1051),
    .C1(net157),
    .X(_0515_));
 sky130_fd_sc_hd__or2_1 _3173_ (.A(\last_addr[7] ),
    .B(_1581_),
    .X(_1590_));
 sky130_fd_sc_hd__o211a_1 _3174_ (.A1(net1074),
    .A2(_1582_),
    .B1(_1590_),
    .C1(net156),
    .X(_0516_));
 sky130_fd_sc_hd__or2_1 _3175_ (.A(net1063),
    .B(_1581_),
    .X(_1591_));
 sky130_fd_sc_hd__o211a_1 _3176_ (.A1(\ROM_addr_buff[8] ),
    .A2(_1582_),
    .B1(net1064),
    .C1(net156),
    .X(_0517_));
 sky130_fd_sc_hd__or2_1 _3177_ (.A(net1044),
    .B(_1581_),
    .X(_1592_));
 sky130_fd_sc_hd__o211a_1 _3178_ (.A1(\ROM_addr_buff[9] ),
    .A2(_1582_),
    .B1(net1045),
    .C1(net156),
    .X(_0518_));
 sky130_fd_sc_hd__or2_1 _3179_ (.A(\last_addr[10] ),
    .B(_1581_),
    .X(_1593_));
 sky130_fd_sc_hd__o211a_1 _3180_ (.A1(net1016),
    .A2(_1582_),
    .B1(_1593_),
    .C1(net156),
    .X(_0519_));
 sky130_fd_sc_hd__or2_1 _3181_ (.A(\last_addr[11] ),
    .B(_1581_),
    .X(_1594_));
 sky130_fd_sc_hd__o211a_1 _3182_ (.A1(net1126),
    .A2(_1582_),
    .B1(_1594_),
    .C1(net155),
    .X(_0520_));
 sky130_fd_sc_hd__nand2_1 _3183_ (.A(net1009),
    .B(net108),
    .Y(_1595_));
 sky130_fd_sc_hd__a21oi_1 _3184_ (.A1(_1483_),
    .A2(net1010),
    .B1(net148),
    .Y(_0521_));
 sky130_fd_sc_hd__nor2_4 _3185_ (.A(_1071_),
    .B(_1161_),
    .Y(_1596_));
 sky130_fd_sc_hd__mux2_1 _3186_ (.A0(net209),
    .A1(net95),
    .S(_1596_),
    .X(_0522_));
 sky130_fd_sc_hd__mux2_1 _3187_ (.A0(net301),
    .A1(net91),
    .S(_1596_),
    .X(_0523_));
 sky130_fd_sc_hd__mux2_1 _3188_ (.A0(net345),
    .A1(net86),
    .S(_1596_),
    .X(_0524_));
 sky130_fd_sc_hd__mux2_1 _3189_ (.A0(net277),
    .A1(net81),
    .S(_1596_),
    .X(_0525_));
 sky130_fd_sc_hd__mux2_1 _3190_ (.A0(net259),
    .A1(net77),
    .S(_1596_),
    .X(_0526_));
 sky130_fd_sc_hd__mux2_1 _3191_ (.A0(net237),
    .A1(net73),
    .S(_1596_),
    .X(_0527_));
 sky130_fd_sc_hd__or2_4 _3192_ (.A(_1007_),
    .B(_1071_),
    .X(_1597_));
 sky130_fd_sc_hd__mux2_1 _3193_ (.A0(net93),
    .A1(net719),
    .S(_1597_),
    .X(_0528_));
 sky130_fd_sc_hd__mux2_1 _3194_ (.A0(net88),
    .A1(net407),
    .S(_1597_),
    .X(_0529_));
 sky130_fd_sc_hd__mux2_1 _3195_ (.A0(net83),
    .A1(net705),
    .S(_1597_),
    .X(_0530_));
 sky130_fd_sc_hd__mux2_1 _3196_ (.A0(net80),
    .A1(net365),
    .S(_1597_),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_1 _3197_ (.A0(net75),
    .A1(net869),
    .S(_1597_),
    .X(_0532_));
 sky130_fd_sc_hd__mux2_1 _3198_ (.A0(net72),
    .A1(net701),
    .S(_1597_),
    .X(_0533_));
 sky130_fd_sc_hd__nor2_4 _3199_ (.A(_1089_),
    .B(_1171_),
    .Y(_1598_));
 sky130_fd_sc_hd__mux2_1 _3200_ (.A0(net447),
    .A1(net95),
    .S(_1598_),
    .X(_0534_));
 sky130_fd_sc_hd__mux2_1 _3201_ (.A0(net303),
    .A1(net91),
    .S(_1598_),
    .X(_0535_));
 sky130_fd_sc_hd__mux2_1 _3202_ (.A0(net855),
    .A1(net86),
    .S(_1598_),
    .X(_0536_));
 sky130_fd_sc_hd__mux2_1 _3203_ (.A0(net599),
    .A1(net81),
    .S(_1598_),
    .X(_0537_));
 sky130_fd_sc_hd__mux2_1 _3204_ (.A0(net771),
    .A1(net77),
    .S(_1598_),
    .X(_0538_));
 sky130_fd_sc_hd__mux2_1 _3205_ (.A0(net521),
    .A1(net73),
    .S(_1598_),
    .X(_0539_));
 sky130_fd_sc_hd__dfxtp_1 _3206_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(net570),
    .Q(\RAM[50][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3207_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net344),
    .Q(\RAM[50][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3208_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(net270),
    .Q(\RAM[50][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3209_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net264),
    .Q(\RAM[50][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3210_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(net490),
    .Q(\RAM[50][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3211_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net204),
    .Q(\RAM[50][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3212_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net580),
    .Q(\RAM[45][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3213_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net538),
    .Q(\RAM[45][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3214_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net904),
    .Q(\RAM[45][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3215_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net368),
    .Q(\RAM[45][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3216_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net942),
    .Q(\RAM[45][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3217_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net788),
    .Q(\RAM[45][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3218_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(net852),
    .Q(\RAM[51][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3219_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net544),
    .Q(\RAM[51][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3220_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(net864),
    .Q(\RAM[51][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3221_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net884),
    .Q(\RAM[51][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3222_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(net558),
    .Q(\RAM[51][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3223_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net646),
    .Q(\RAM[51][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3224_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net1183),
    .Q(\mem_cycle[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3225_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net1190),
    .Q(\mem_cycle[1] ));
 sky130_fd_sc_hd__dfxtp_2 _3226_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(net1207),
    .Q(\mem_cycle[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3227_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net1179),
    .Q(\mem_cycle[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3228_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net1169),
    .Q(\mem_cycle[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3229_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net324),
    .Q(\RAM[52][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3230_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net202),
    .Q(\RAM[52][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3231_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net354),
    .Q(\RAM[52][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3232_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net420),
    .Q(\RAM[52][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3233_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net386),
    .Q(\RAM[52][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3234_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net182),
    .Q(\RAM[52][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3235_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net780),
    .Q(\RAM[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3236_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net918),
    .Q(\RAM[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3237_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net640),
    .Q(\RAM[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3238_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net718),
    .Q(\RAM[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3239_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net714),
    .Q(\RAM[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3240_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net674),
    .Q(\RAM[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3241_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(net1035),
    .Q(\ROM_dest[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3242_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(net1015),
    .Q(\ROM_dest[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3243_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(net1095),
    .Q(\ROM_dest[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3244_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net966),
    .Q(\RAM[53][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3245_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net876),
    .Q(\RAM[53][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3246_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net944),
    .Q(\RAM[53][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3247_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net928),
    .Q(\RAM[53][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3248_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net636),
    .Q(\RAM[53][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3249_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net954),
    .Q(\RAM[53][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3250_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net638),
    .Q(\RAM[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3251_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net732),
    .Q(\RAM[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3252_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net436),
    .Q(\RAM[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3253_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net836),
    .Q(\RAM[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3254_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net734),
    .Q(\RAM[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3255_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net746),
    .Q(\RAM[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3256_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net374),
    .Q(\RAM[54][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3257_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net458),
    .Q(\RAM[54][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3258_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net340),
    .Q(\RAM[54][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3259_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net582),
    .Q(\RAM[54][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3260_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net356),
    .Q(\RAM[54][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3261_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net498),
    .Q(\RAM[54][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3262_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net696),
    .Q(\RAM[39][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3263_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net556),
    .Q(\RAM[39][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3264_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net678),
    .Q(\RAM[39][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3265_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net692),
    .Q(\RAM[39][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3266_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net518),
    .Q(\RAM[39][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3267_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net868),
    .Q(\RAM[39][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3268_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net770),
    .Q(\RAM[55][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3269_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net730),
    .Q(\RAM[55][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3270_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net722),
    .Q(\RAM[55][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3271_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net950),
    .Q(\RAM[55][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3272_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net878),
    .Q(\RAM[55][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3273_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net738),
    .Q(\RAM[55][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3274_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(net442),
    .Q(\RAM[49][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3275_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net254),
    .Q(\RAM[49][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3276_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(net224),
    .Q(\RAM[49][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3277_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(net200),
    .Q(\RAM[49][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3278_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net180),
    .Q(\RAM[49][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3279_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(net244),
    .Q(\RAM[49][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3280_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net364),
    .Q(\RAM[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3281_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net308),
    .Q(\RAM[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3282_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net592),
    .Q(\RAM[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3283_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net314),
    .Q(\RAM[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3284_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net326),
    .Q(\RAM[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3285_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net846),
    .Q(\RAM[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3286_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net934),
    .Q(\RAM[43][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3287_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net858),
    .Q(\RAM[43][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3288_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net510),
    .Q(\RAM[43][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3289_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net824),
    .Q(\RAM[43][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3290_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net658),
    .Q(\RAM[43][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3291_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net584),
    .Q(\RAM[43][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3292_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_0107_),
    .Q(net46));
 sky130_fd_sc_hd__dfxtp_1 _3293_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_0108_),
    .Q(net47));
 sky130_fd_sc_hd__dfxtp_1 _3294_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0109_),
    .Q(net48));
 sky130_fd_sc_hd__dfxtp_1 _3295_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net1222),
    .Q(net49));
 sky130_fd_sc_hd__dfxtp_1 _3296_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net1202),
    .Q(net50));
 sky130_fd_sc_hd__dfxtp_1 _3297_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net1214),
    .Q(net52));
 sky130_fd_sc_hd__dfxtp_1 _3298_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net616),
    .Q(\RAM[57][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3299_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net530),
    .Q(\RAM[57][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3300_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net682),
    .Q(\RAM[57][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3301_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net838),
    .Q(\RAM[57][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3302_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net756),
    .Q(\RAM[57][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3303_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net812),
    .Q(\RAM[57][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3304_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(net310),
    .Q(\RAM[48][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3305_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net234),
    .Q(\RAM[48][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3306_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(net230),
    .Q(\RAM[48][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3307_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(net252),
    .Q(\RAM[48][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3308_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net268),
    .Q(\RAM[48][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3309_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(net220),
    .Q(\RAM[48][5] ));
 sky130_fd_sc_hd__dfxtp_2 _3310_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_0021_),
    .Q(net53));
 sky130_fd_sc_hd__dfxtp_1 _3311_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(net1111),
    .Q(\instr_cycle[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3312_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_0023_),
    .Q(\instr_cycle[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3313_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(net1220),
    .Q(net64));
 sky130_fd_sc_hd__dfxtp_1 _3314_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(net1019),
    .Q(net65));
 sky130_fd_sc_hd__dfxtp_1 _3315_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(net1021),
    .Q(net66));
 sky130_fd_sc_hd__dfxtp_1 _3316_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net802),
    .Q(\RAM[46][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3317_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net594),
    .Q(\RAM[46][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3318_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net924),
    .Q(\RAM[46][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3319_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net484),
    .Q(\RAM[46][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3320_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net590),
    .Q(\RAM[46][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3321_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net922),
    .Q(\RAM[46][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3322_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net962),
    .Q(\RAM[59][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3323_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0135_),
    .Q(\RAM[59][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3324_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(_0136_),
    .Q(\RAM[59][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3325_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(_0137_),
    .Q(\RAM[59][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3326_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(_0138_),
    .Q(\RAM[59][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3327_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_0139_),
    .Q(\RAM[59][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3328_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0140_),
    .Q(net55));
 sky130_fd_sc_hd__dfxtp_1 _3329_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0141_),
    .Q(net56));
 sky130_fd_sc_hd__dfxtp_1 _3330_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0142_),
    .Q(net57));
 sky130_fd_sc_hd__dfxtp_1 _3331_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0143_),
    .Q(net58));
 sky130_fd_sc_hd__dfxtp_1 _3332_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0144_),
    .Q(net59));
 sky130_fd_sc_hd__dfxtp_1 _3333_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0145_),
    .Q(net60));
 sky130_fd_sc_hd__dfxtp_1 _3334_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net844),
    .Q(\RAM[47][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3335_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net502),
    .Q(\RAM[47][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3336_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net956),
    .Q(\RAM[47][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3337_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net470),
    .Q(\RAM[47][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3338_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net672),
    .Q(\RAM[47][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3339_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net854),
    .Q(\RAM[47][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3340_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net376),
    .Q(\RAM[56][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3341_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net216),
    .Q(\RAM[56][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3342_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net312),
    .Q(\RAM[56][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3343_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net294),
    .Q(\RAM[56][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3344_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net266),
    .Q(\RAM[56][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3345_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net236),
    .Q(\RAM[56][5] ));
 sky130_fd_sc_hd__dfxtp_2 _3346_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_0000_),
    .Q(\MAR[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3347_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(net1217),
    .Q(\MAR[1] ));
 sky130_fd_sc_hd__dfxtp_2 _3348_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_0002_),
    .Q(\MAR[2] ));
 sky130_fd_sc_hd__dfxtp_2 _3349_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0003_),
    .Q(\MAR[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3350_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(_0004_),
    .Q(\MAR[4] ));
 sky130_fd_sc_hd__dfxtp_2 _3351_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(net1200),
    .Q(net61));
 sky130_fd_sc_hd__dfxtp_1 _3352_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net926),
    .Q(\RAM[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3353_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net642),
    .Q(\RAM[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3354_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net914),
    .Q(\RAM[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3355_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net814),
    .Q(\RAM[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3356_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net688),
    .Q(\RAM[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3357_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net680),
    .Q(\RAM[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3358_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net930),
    .Q(\RAM[42][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3359_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net932),
    .Q(\RAM[42][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3360_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net542),
    .Q(\RAM[42][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3361_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net968),
    .Q(\RAM[42][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3362_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net742),
    .Q(\RAM[42][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3363_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net472),
    .Q(\RAM[42][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3364_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net952),
    .Q(\RAM[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3365_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net818),
    .Q(\RAM[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3366_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net654),
    .Q(\RAM[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3367_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net724),
    .Q(\RAM[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3368_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net648),
    .Q(\RAM[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3369_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net656),
    .Q(\RAM[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3370_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net716),
    .Q(\RAM[41][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3371_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net578),
    .Q(\RAM[41][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3372_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net832),
    .Q(\RAM[41][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3373_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net874),
    .Q(\RAM[41][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3374_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net552),
    .Q(\RAM[41][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3375_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net900),
    .Q(\RAM[41][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3376_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net306),
    .Q(\RAM[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3377_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net804),
    .Q(\RAM[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3378_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net764),
    .Q(\RAM[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3379_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net888),
    .Q(\RAM[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3380_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net534),
    .Q(\RAM[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3381_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net834),
    .Q(\RAM[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3382_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net348),
    .Q(\RAM[40][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3383_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net282),
    .Q(\RAM[40][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3384_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net828),
    .Q(\RAM[40][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3385_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net912),
    .Q(\RAM[40][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3386_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net296),
    .Q(\RAM[40][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3387_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net396),
    .Q(\RAM[40][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3388_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net322),
    .Q(\RAM[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3389_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net496),
    .Q(\RAM[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3390_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net262),
    .Q(\RAM[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3391_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net456),
    .Q(\RAM[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3392_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net488),
    .Q(\RAM[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3393_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net336),
    .Q(\RAM[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3394_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net920),
    .Q(\RAM[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3395_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net526),
    .Q(\RAM[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3396_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net940),
    .Q(\RAM[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3397_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net808),
    .Q(\RAM[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3398_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net524),
    .Q(\RAM[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3399_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net752),
    .Q(\RAM[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3400_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net1120),
    .Q(net69));
 sky130_fd_sc_hd__dfxtp_1 _3401_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_0207_),
    .Q(net41));
 sky130_fd_sc_hd__dfxtp_1 _3402_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_0208_),
    .Q(net42));
 sky130_fd_sc_hd__dfxtp_1 _3403_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net1060),
    .Q(net43));
 sky130_fd_sc_hd__dfxtp_1 _3404_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_0210_),
    .Q(net44));
 sky130_fd_sc_hd__dfxtp_1 _3405_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_0211_),
    .Q(net45));
 sky130_fd_sc_hd__dfxtp_1 _3406_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net754),
    .Q(\RAM[38][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3407_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net960),
    .Q(\RAM[38][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3408_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net896),
    .Q(\RAM[38][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3409_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net816),
    .Q(\RAM[38][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3410_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net728),
    .Q(\RAM[38][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3411_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net898),
    .Q(\RAM[38][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3412_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net188),
    .Q(\RAM[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3413_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net212),
    .Q(\RAM[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3414_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net184),
    .Q(\RAM[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3415_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net494),
    .Q(\RAM[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3416_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net214),
    .Q(\RAM[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3417_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net284),
    .Q(\RAM[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3418_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net460),
    .Q(\RAM[37][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3419_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net512),
    .Q(\RAM[37][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3420_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net872),
    .Q(\RAM[37][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3421_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net916),
    .Q(\RAM[37][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3422_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net978),
    .Q(\RAM[37][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3423_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net794),
    .Q(\RAM[37][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3424_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net446),
    .Q(\RAM[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3425_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net412),
    .Q(\RAM[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3426_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net410),
    .Q(\RAM[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3427_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net766),
    .Q(\RAM[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3428_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net710),
    .Q(\RAM[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3429_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net430),
    .Q(\RAM[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3430_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net486),
    .Q(\RAM[36][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3431_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net384),
    .Q(\RAM[36][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3432_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net350),
    .Q(\RAM[36][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3433_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net318),
    .Q(\RAM[36][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3434_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net650),
    .Q(\RAM[36][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3435_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net532),
    .Q(\RAM[36][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3436_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net560),
    .Q(\RAM[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3437_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net232),
    .Q(\RAM[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3438_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net248),
    .Q(\RAM[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3439_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net432),
    .Q(\RAM[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3440_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net240),
    .Q(\RAM[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3441_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net208),
    .Q(\RAM[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3442_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(net404),
    .Q(\RAM[61][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3443_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(net628),
    .Q(\RAM[61][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3444_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net860),
    .Q(\RAM[61][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3445_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net620),
    .Q(\RAM[61][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3446_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net508),
    .Q(\RAM[61][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3447_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net866),
    .Q(\RAM[61][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3448_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net1002),
    .Q(\imm_buff[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3449_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net1012),
    .Q(\imm_buff[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3450_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net776),
    .Q(\RAM[35][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3451_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net782),
    .Q(\RAM[35][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3452_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net660),
    .Q(\RAM[35][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3453_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net454),
    .Q(\RAM[35][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3454_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net666),
    .Q(\RAM[35][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3455_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net842),
    .Q(\RAM[35][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3456_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net372),
    .Q(\RAM[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3457_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net694),
    .Q(\RAM[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3458_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net466),
    .Q(\RAM[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3459_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net300),
    .Q(\RAM[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3460_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net190),
    .Q(\RAM[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3461_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net462),
    .Q(\RAM[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3462_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net434),
    .Q(\RAM[34][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3463_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net328),
    .Q(\RAM[34][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3464_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net390),
    .Q(\RAM[34][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3465_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net664),
    .Q(\RAM[34][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3466_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net280),
    .Q(\RAM[34][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3467_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net708),
    .Q(\RAM[34][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3468_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net704),
    .Q(\RAM[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3469_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net316),
    .Q(\RAM[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3470_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net360),
    .Q(\RAM[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3471_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net256),
    .Q(\RAM[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3472_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net474),
    .Q(\RAM[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3473_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net504),
    .Q(\RAM[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3474_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net196),
    .Q(\RAM[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3475_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net276),
    .Q(\RAM[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3476_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net424),
    .Q(\RAM[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3477_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net700),
    .Q(\RAM[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3478_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net452),
    .Q(\RAM[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3479_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net468),
    .Q(\RAM[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3480_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net338),
    .Q(\RAM[33][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3481_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net246),
    .Q(\RAM[33][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3482_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net392),
    .Q(\RAM[33][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3483_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net444),
    .Q(\RAM[33][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3484_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net274),
    .Q(\RAM[33][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3485_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net194),
    .Q(\RAM[33][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3486_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net820),
    .Q(\RAM[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3487_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net906),
    .Q(\RAM[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3488_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net830),
    .Q(\RAM[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3489_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net618),
    .Q(\RAM[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3490_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net908),
    .Q(\RAM[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3491_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net848),
    .Q(\RAM[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3492_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net198),
    .Q(\RAM[32][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3493_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net380),
    .Q(\RAM[32][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3494_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net298),
    .Q(\RAM[32][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3495_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net192),
    .Q(\RAM[32][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3496_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net398),
    .Q(\RAM[32][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3497_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net500),
    .Q(\RAM[32][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3498_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net362),
    .Q(\RAM[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3499_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net320),
    .Q(\RAM[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3500_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net414),
    .Q(\RAM[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3501_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net288),
    .Q(\RAM[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3502_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net422),
    .Q(\RAM[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3503_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net604),
    .Q(\RAM[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3504_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net892),
    .Q(\RAM[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3505_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net822),
    .Q(\RAM[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3506_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net806),
    .Q(\RAM[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3507_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net606),
    .Q(\RAM[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3508_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net632),
    .Q(\RAM[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3509_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net880),
    .Q(\RAM[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3510_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net624),
    .Q(\RAM[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3511_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net358),
    .Q(\RAM[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3512_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net726),
    .Q(\RAM[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3513_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net402),
    .Q(\RAM[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3514_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net400),
    .Q(\RAM[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3515_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net608),
    .Q(\RAM[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3516_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net902),
    .Q(\RAM[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3517_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net894),
    .Q(\RAM[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3518_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net540),
    .Q(\RAM[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3519_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net686),
    .Q(\RAM[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3520_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net520),
    .Q(\RAM[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3521_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net622),
    .Q(\RAM[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3522_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net406),
    .Q(\RAM[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3523_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net550),
    .Q(\RAM[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3524_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net948),
    .Q(\RAM[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3525_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net976),
    .Q(\RAM[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3526_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net970),
    .Q(\RAM[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3527_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net936),
    .Q(\RAM[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3528_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net272),
    .Q(\RAM[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3529_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net290),
    .Q(\RAM[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3530_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net370),
    .Q(\RAM[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3531_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net222),
    .Q(\RAM[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3532_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net352),
    .Q(\RAM[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3533_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net450),
    .Q(\RAM[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3534_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net438),
    .Q(\RAM[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3535_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net574),
    .Q(\RAM[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3536_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net790),
    .Q(\RAM[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3537_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net712),
    .Q(\RAM[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3538_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net736),
    .Q(\RAM[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3539_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net792),
    .Q(\RAM[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3540_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net850),
    .Q(\RAM[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3541_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net644),
    .Q(\RAM[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3542_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net684),
    .Q(\RAM[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3543_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net662),
    .Q(\RAM[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3544_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net862),
    .Q(\RAM[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3545_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net610),
    .Q(\RAM[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3546_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net226),
    .Q(\RAM[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3547_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net334),
    .Q(\RAM[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3548_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net286),
    .Q(\RAM[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3549_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net670),
    .Q(\RAM[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3550_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net186),
    .Q(\RAM[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3551_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net250),
    .Q(\RAM[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3552_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net958),
    .Q(\RAM[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3553_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net882),
    .Q(\RAM[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3554_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net910),
    .Q(\RAM[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3555_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net890),
    .Q(\RAM[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3556_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net760),
    .Q(\RAM[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3557_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net740),
    .Q(\RAM[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3558_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net242),
    .Q(\RAM[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3559_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net758),
    .Q(\RAM[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3560_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net440),
    .Q(\RAM[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3561_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net206),
    .Q(\RAM[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3562_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net388),
    .Q(\RAM[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3563_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net546),
    .Q(\RAM[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3564_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net810),
    .Q(\RAM[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3565_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net974),
    .Q(\RAM[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3566_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net426),
    .Q(\RAM[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3567_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net840),
    .Q(\RAM[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3568_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net778),
    .Q(\RAM[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3569_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net690),
    .Q(\RAM[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3570_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net228),
    .Q(\RAM[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3571_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net798),
    .Q(\RAM[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3572_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net598),
    .Q(\RAM[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3573_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net784),
    .Q(\RAM[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3574_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net330),
    .Q(\RAM[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3575_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net478),
    .Q(\RAM[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3576_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(net630),
    .Q(\RAM[62][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3577_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(net516),
    .Q(\RAM[62][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3578_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net536),
    .Q(\RAM[62][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3579_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(net634),
    .Q(\RAM[62][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3580_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net562),
    .Q(\RAM[62][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3581_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net576),
    .Q(\RAM[62][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3582_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net612),
    .Q(\RAM[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3583_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net548),
    .Q(\RAM[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3584_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net292),
    .Q(\RAM[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3585_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net482),
    .Q(\RAM[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3586_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net572),
    .Q(\RAM[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3587_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net480),
    .Q(\RAM[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3588_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net416),
    .Q(\RAM[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3589_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net332),
    .Q(\RAM[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3590_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net382),
    .Q(\RAM[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3591_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net566),
    .Q(\RAM[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3592_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net342),
    .Q(\RAM[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3593_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net394),
    .Q(\RAM[1][5] ));
 sky130_fd_sc_hd__dfxtp_2 _3594_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(net1087),
    .Q(\A[0] ));
 sky130_fd_sc_hd__dfxtp_2 _3595_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(net1097),
    .Q(\A[1] ));
 sky130_fd_sc_hd__dfxtp_4 _3596_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net1102),
    .Q(\A[2] ));
 sky130_fd_sc_hd__dfxtp_2 _3597_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net1072),
    .Q(\A[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3598_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net1083),
    .Q(\A[4] ));
 sky130_fd_sc_hd__dfxtp_2 _3599_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(net1113),
    .Q(\A[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3600_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(net1157),
    .Q(\B[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3601_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net1122),
    .Q(\B[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3602_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net1029),
    .Q(\B[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3603_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net1129),
    .Q(\B[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3604_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net1031),
    .Q(\B[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3605_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(net1104),
    .Q(\B[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3606_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_0006_),
    .Q(\P[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3607_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(_0007_),
    .Q(\P[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3608_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_0008_),
    .Q(\P[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3609_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(_0009_),
    .Q(\P[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3610_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0010_),
    .Q(\P[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3611_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(net1187),
    .Q(\P[5] ));
 sky130_fd_sc_hd__dfxtp_4 _3612_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(_0412_),
    .Q(net51));
 sky130_fd_sc_hd__dfxtp_4 _3613_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(net1230),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_1 _3614_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net1054),
    .Q(\PC[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3615_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_0415_),
    .Q(\PC[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3616_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(net1027),
    .Q(\PC[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3617_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net1023),
    .Q(\PC[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3618_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net1177),
    .Q(\PC[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3619_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net1033),
    .Q(\PC[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3620_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net1085),
    .Q(\PC[6] ));
 sky130_fd_sc_hd__dfxtp_2 _3621_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0421_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_2 _3622_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_0422_),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_2 _3623_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_0423_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_1 _3624_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0424_),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_1 _3625_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0425_),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_2 _3626_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_0012_),
    .Q(\insin[0] ));
 sky130_fd_sc_hd__dfxtp_2 _3627_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(_0013_),
    .Q(\insin[1] ));
 sky130_fd_sc_hd__dfxtp_2 _3628_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(net1162),
    .Q(\insin[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3629_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(net1152),
    .Q(\insin[3] ));
 sky130_fd_sc_hd__dfxtp_4 _3630_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(net1185),
    .Q(\insin[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3631_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(net1081),
    .Q(\insin[5] ));
 sky130_fd_sc_hd__dfxtp_2 _3632_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(net1040),
    .Q(net54));
 sky130_fd_sc_hd__dfxtp_1 _3633_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(net602),
    .Q(\imm_buff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3634_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(net796),
    .Q(\imm_buff[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3635_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net994),
    .Q(\imm_buff[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3636_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net1006),
    .Q(\imm_buff[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3637_ (.CLK(clknet_leaf_54_wb_clk_i),
    .D(net428),
    .Q(\last_PC[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3638_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(net218),
    .Q(\last_PC[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3639_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(net774),
    .Q(\last_PC[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3640_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net750),
    .Q(\last_PC[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3641_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net568),
    .Q(\last_PC[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3642_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net676),
    .Q(\last_PC[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3643_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(net378),
    .Q(\last_PC[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3644_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net476),
    .Q(\last_PC[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3645_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(net492),
    .Q(\last_PC[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3646_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(net588),
    .Q(\last_PC[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3647_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net626),
    .Q(\last_PC[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3648_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net528),
    .Q(\last_PC[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3649_ (.CLK(clknet_leaf_56_wb_clk_i),
    .D(net972),
    .Q(\last_flags[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3650_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(net998),
    .Q(\last_flags[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3651_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(net586),
    .Q(\last_A[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3652_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(net762),
    .Q(\last_A[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3653_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net886),
    .Q(\last_A[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3654_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net748),
    .Q(\last_A[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3655_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net744),
    .Q(\last_A[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3656_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(net938),
    .Q(\last_A[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3657_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(net800),
    .Q(\last_B[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3658_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net826),
    .Q(\last_B[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3659_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net506),
    .Q(\last_B[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3660_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net786),
    .Q(\last_B[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3661_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net514),
    .Q(\last_B[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3662_ (.CLK(clknet_leaf_57_wb_clk_i),
    .D(net258),
    .Q(\last_B[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3663_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(net698),
    .Q(\last_MAR[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3664_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(net668),
    .Q(\last_MAR[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3665_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net768),
    .Q(\last_MAR[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3666_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(net614),
    .Q(\last_MAR[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3667_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(net596),
    .Q(\last_MAR[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3668_ (.CLK(clknet_leaf_53_wb_clk_i),
    .D(net652),
    .Q(\last_MAR[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3669_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(net418),
    .Q(\last_P[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3670_ (.CLK(clknet_leaf_55_wb_clk_i),
    .D(net984),
    .Q(\last_P[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3671_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net564),
    .Q(\last_P[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3672_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net464),
    .Q(\last_P[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3673_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net946),
    .Q(\last_P[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3674_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net554),
    .Q(\last_P[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3675_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(net980),
    .Q(needs_irupt));
 sky130_fd_sc_hd__dfxtp_2 _3676_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(net1118),
    .Q(net62));
 sky130_fd_sc_hd__dfxtp_2 _3677_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0471_),
    .Q(\ROM_spi_cycle[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3678_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net1233),
    .Q(\ROM_spi_cycle[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3679_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net1100),
    .Q(\ROM_spi_cycle[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3680_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net1109),
    .Q(\ROM_spi_cycle[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3681_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net1225),
    .Q(\ROM_spi_cycle[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3682_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net1165),
    .Q(\startup_cycle[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3683_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net1008),
    .Q(\startup_cycle[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3684_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net1125),
    .Q(\startup_cycle[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3685_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net1235),
    .Q(\startup_cycle[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3686_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(net1089),
    .Q(\startup_cycle[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3687_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(net1210),
    .Q(\startup_cycle[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3688_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(net1091),
    .Q(\startup_cycle[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3689_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_0483_),
    .Q(last_inter));
 sky130_fd_sc_hd__dfxtp_1 _3690_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net1025),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_1 _3691_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_0485_),
    .Q(net68));
 sky130_fd_sc_hd__dfxtp_1 _3692_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(_0486_),
    .Q(net63));
 sky130_fd_sc_hd__dfxtp_1 _3693_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_0487_),
    .Q(ROM_OEB));
 sky130_fd_sc_hd__dfxtp_1 _3694_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_0488_),
    .Q(ROM_spi_mode));
 sky130_fd_sc_hd__dfxtp_1 _3695_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(_0489_),
    .Q(\ROM_spi_dat_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3696_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net982),
    .Q(\ROM_spi_dat_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3697_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net1004),
    .Q(\ROM_spi_dat_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3698_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net996),
    .Q(\ROM_spi_dat_out[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3699_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net1000),
    .Q(\ROM_spi_dat_out[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3700_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net988),
    .Q(\ROM_spi_dat_out[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3701_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net990),
    .Q(\ROM_spi_dat_out[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3702_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net992),
    .Q(\ROM_spi_dat_out[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3703_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net1077),
    .Q(\ROM_addr_buff[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3704_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net1132),
    .Q(\ROM_addr_buff[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3705_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net1136),
    .Q(\ROM_addr_buff[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3706_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net1145),
    .Q(\ROM_addr_buff[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3707_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net1139),
    .Q(\ROM_addr_buff[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3708_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net1037),
    .Q(\ROM_addr_buff[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3709_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net1093),
    .Q(\ROM_addr_buff[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3710_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net1155),
    .Q(\ROM_addr_buff[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3711_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net1181),
    .Q(\ROM_addr_buff[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3712_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net1194),
    .Q(\ROM_addr_buff[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3713_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net1068),
    .Q(\ROM_addr_buff[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3714_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_0508_),
    .Q(\ROM_addr_buff[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3715_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(net1143),
    .Q(\last_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _3716_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net1115),
    .Q(\last_addr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _3717_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net1057),
    .Q(\last_addr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _3718_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net1043),
    .Q(\last_addr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _3719_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(net1106),
    .Q(\last_addr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _3720_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(net1049),
    .Q(\last_addr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _3721_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(net1052),
    .Q(\last_addr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _3722_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(net1075),
    .Q(\last_addr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _3723_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(net1065),
    .Q(\last_addr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _3724_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(net1046),
    .Q(\last_addr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _3725_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net1017),
    .Q(\last_addr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _3726_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net1127),
    .Q(\last_addr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _3727_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(_0521_),
    .Q(spi_clkdiv));
 sky130_fd_sc_hd__dfxtp_1 _3728_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net210),
    .Q(\RAM[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3729_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net302),
    .Q(\RAM[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3730_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net346),
    .Q(\RAM[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3731_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net278),
    .Q(\RAM[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3732_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net260),
    .Q(\RAM[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3733_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net238),
    .Q(\RAM[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3734_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net720),
    .Q(\RAM[44][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3735_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net408),
    .Q(\RAM[44][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3736_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net706),
    .Q(\RAM[44][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3737_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net366),
    .Q(\RAM[44][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3738_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net870),
    .Q(\RAM[44][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3739_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net702),
    .Q(\RAM[44][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3740_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net448),
    .Q(\RAM[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3741_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net304),
    .Q(\RAM[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3742_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net856),
    .Q(\RAM[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3743_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net600),
    .Q(\RAM[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3744_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net772),
    .Q(\RAM[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3745_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net522),
    .Q(\RAM[9][5] ));
 sky130_fd_sc_hd__buf_1 _3767_ (.A(net38),
    .X(net35));
 sky130_fd_sc_hd__buf_1 _3768_ (.A(net38),
    .X(net37));
 sky130_fd_sc_hd__buf_1 _3769_ (.A(net19),
    .X(net39));
 sky130_fd_sc_hd__buf_1 _3770_ (.A(net21),
    .X(net20));
 sky130_fd_sc_hd__buf_1 _3771_ (.A(net23),
    .X(net22));
 sky130_fd_sc_hd__buf_1 _3772_ (.A(net25),
    .X(net24));
 sky130_fd_sc_hd__buf_1 _3773_ (.A(net27),
    .X(net26));
 sky130_fd_sc_hd__buf_1 _3774_ (.A(net29),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_4__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_5__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_6__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_3_7__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.A(clknet_3_4__leaf_wb_clk_i),
    .X(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.A(clknet_3_4__leaf_wb_clk_i),
    .X(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.A(clknet_3_5__leaf_wb_clk_i),
    .X(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.A(clknet_3_4__leaf_wb_clk_i),
    .X(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.A(clknet_3_7__leaf_wb_clk_i),
    .X(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.A(clknet_3_7__leaf_wb_clk_i),
    .X(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.A(clknet_3_7__leaf_wb_clk_i),
    .X(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.A(clknet_3_7__leaf_wb_clk_i),
    .X(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.A(clknet_3_7__leaf_wb_clk_i),
    .X(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.A(clknet_3_7__leaf_wb_clk_i),
    .X(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.A(clknet_3_7__leaf_wb_clk_i),
    .X(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.A(clknet_3_1__leaf_wb_clk_i),
    .X(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.A(clknet_3_7__leaf_wb_clk_i),
    .X(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.A(clknet_3_6__leaf_wb_clk_i),
    .X(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.A(clknet_3_3__leaf_wb_clk_i),
    .X(clknet_leaf_37_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.A(clknet_3_3__leaf_wb_clk_i),
    .X(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.A(clknet_3_3__leaf_wb_clk_i),
    .X(clknet_leaf_39_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.A(clknet_3_1__leaf_wb_clk_i),
    .X(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.A(clknet_3_3__leaf_wb_clk_i),
    .X(clknet_leaf_40_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.A(clknet_3_3__leaf_wb_clk_i),
    .X(clknet_leaf_41_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.A(clknet_3_3__leaf_wb_clk_i),
    .X(clknet_leaf_42_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.A(clknet_3_2__leaf_wb_clk_i),
    .X(clknet_leaf_43_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.A(clknet_3_2__leaf_wb_clk_i),
    .X(clknet_leaf_44_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.A(clknet_3_2__leaf_wb_clk_i),
    .X(clknet_leaf_45_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.A(clknet_3_2__leaf_wb_clk_i),
    .X(clknet_leaf_46_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.A(clknet_3_2__leaf_wb_clk_i),
    .X(clknet_leaf_47_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.A(clknet_3_2__leaf_wb_clk_i),
    .X(clknet_leaf_48_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.A(clknet_3_2__leaf_wb_clk_i),
    .X(clknet_leaf_49_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.A(clknet_3_1__leaf_wb_clk_i),
    .X(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.A(clknet_3_3__leaf_wb_clk_i),
    .X(clknet_leaf_50_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.A(clknet_3_3__leaf_wb_clk_i),
    .X(clknet_leaf_51_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.A(clknet_3_1__leaf_wb_clk_i),
    .X(clknet_leaf_52_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.A(clknet_3_1__leaf_wb_clk_i),
    .X(clknet_leaf_53_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_54_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_55_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_56_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_wb_clk_i (.A(clknet_3_0__leaf_wb_clk_i),
    .X(clknet_leaf_57_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.A(clknet_3_1__leaf_wb_clk_i),
    .X(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.A(clknet_3_4__leaf_wb_clk_i),
    .X(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.A(clknet_3_4__leaf_wb_clk_i),
    .X(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.A(clknet_3_4__leaf_wb_clk_i),
    .X(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.A(clknet_3_4__leaf_wb_clk_i),
    .X(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 fanout102 (.A(_0605_),
    .X(net102));
 sky130_fd_sc_hd__buf_6 fanout103 (.A(_0694_),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_8 fanout104 (.A(_0693_),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_8 fanout105 (.A(_0643_),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_8 fanout106 (.A(_0565_),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_4 fanout107 (.A(_0565_),
    .X(net107));
 sky130_fd_sc_hd__buf_4 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__buf_4 fanout110 (.A(net111),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_8 fanout111 (.A(_0560_),
    .X(net111));
 sky130_fd_sc_hd__buf_4 fanout112 (.A(net113),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_8 fanout113 (.A(_0559_),
    .X(net113));
 sky130_fd_sc_hd__buf_4 fanout114 (.A(_0551_),
    .X(net114));
 sky130_fd_sc_hd__buf_4 fanout115 (.A(_0551_),
    .X(net115));
 sky130_fd_sc_hd__buf_8 fanout116 (.A(net1199),
    .X(net116));
 sky130_fd_sc_hd__buf_4 fanout117 (.A(net118),
    .X(net117));
 sky130_fd_sc_hd__buf_4 fanout118 (.A(net1249),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_8 fanout119 (.A(net1211),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_4 fanout120 (.A(\MAR[3] ),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_8 fanout121 (.A(\MAR[3] ),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_4 fanout122 (.A(\MAR[3] ),
    .X(net122));
 sky130_fd_sc_hd__buf_6 fanout123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__buf_8 fanout124 (.A(\MAR[2] ),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_8 fanout125 (.A(net132),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_4 fanout126 (.A(net132),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_8 fanout127 (.A(net132),
    .X(net127));
 sky130_fd_sc_hd__buf_4 fanout128 (.A(net132),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_8 fanout129 (.A(net132),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_8 fanout130 (.A(net131),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_8 fanout131 (.A(net132),
    .X(net131));
 sky130_fd_sc_hd__buf_4 fanout132 (.A(net1216),
    .X(net132));
 sky130_fd_sc_hd__buf_8 fanout133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_8 fanout134 (.A(net1240),
    .X(net134));
 sky130_fd_sc_hd__buf_8 fanout135 (.A(\MAR[0] ),
    .X(net135));
 sky130_fd_sc_hd__buf_4 fanout136 (.A(\MAR[0] ),
    .X(net136));
 sky130_fd_sc_hd__buf_6 fanout137 (.A(net139),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_8 fanout138 (.A(net139),
    .X(net138));
 sky130_fd_sc_hd__buf_4 fanout139 (.A(\MAR[0] ),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_8 fanout140 (.A(net143),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_8 fanout141 (.A(net143),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_4 fanout142 (.A(net143),
    .X(net142));
 sky130_fd_sc_hd__buf_4 fanout143 (.A(\MAR[0] ),
    .X(net143));
 sky130_fd_sc_hd__buf_4 fanout144 (.A(net1166),
    .X(net144));
 sky130_fd_sc_hd__buf_2 fanout145 (.A(net1166),
    .X(net145));
 sky130_fd_sc_hd__buf_6 fanout146 (.A(net1170),
    .X(net146));
 sky130_fd_sc_hd__buf_4 fanout147 (.A(net148),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_4 fanout148 (.A(_0555_),
    .X(net148));
 sky130_fd_sc_hd__buf_4 fanout149 (.A(net150),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_8 fanout150 (.A(net151),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_4 fanout151 (.A(net18),
    .X(net151));
 sky130_fd_sc_hd__buf_4 fanout152 (.A(net157),
    .X(net152));
 sky130_fd_sc_hd__buf_4 fanout153 (.A(net157),
    .X(net153));
 sky130_fd_sc_hd__buf_4 fanout154 (.A(net157),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_2 fanout155 (.A(net157),
    .X(net155));
 sky130_fd_sc_hd__buf_4 fanout156 (.A(net157),
    .X(net156));
 sky130_fd_sc_hd__buf_4 fanout157 (.A(net18),
    .X(net157));
 sky130_fd_sc_hd__buf_4 fanout70 (.A(_1402_),
    .X(net70));
 sky130_fd_sc_hd__buf_4 fanout71 (.A(net72),
    .X(net71));
 sky130_fd_sc_hd__buf_4 fanout72 (.A(_1003_),
    .X(net72));
 sky130_fd_sc_hd__buf_4 fanout73 (.A(net74),
    .X(net73));
 sky130_fd_sc_hd__buf_4 fanout74 (.A(_1003_),
    .X(net74));
 sky130_fd_sc_hd__buf_4 fanout75 (.A(net76),
    .X(net75));
 sky130_fd_sc_hd__buf_4 fanout76 (.A(_1002_),
    .X(net76));
 sky130_fd_sc_hd__buf_4 fanout77 (.A(net78),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_8 fanout78 (.A(_1002_),
    .X(net78));
 sky130_fd_sc_hd__buf_4 fanout79 (.A(net80),
    .X(net79));
 sky130_fd_sc_hd__buf_4 fanout80 (.A(_1001_),
    .X(net80));
 sky130_fd_sc_hd__buf_4 fanout81 (.A(net82),
    .X(net81));
 sky130_fd_sc_hd__buf_4 fanout82 (.A(_1001_),
    .X(net82));
 sky130_fd_sc_hd__buf_4 fanout83 (.A(net85),
    .X(net83));
 sky130_fd_sc_hd__buf_2 fanout84 (.A(net85),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_4 fanout85 (.A(_1000_),
    .X(net85));
 sky130_fd_sc_hd__buf_4 fanout86 (.A(net87),
    .X(net86));
 sky130_fd_sc_hd__buf_4 fanout87 (.A(_1000_),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_4 fanout88 (.A(_0999_),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_4 fanout89 (.A(_0999_),
    .X(net89));
 sky130_fd_sc_hd__buf_4 fanout90 (.A(_0999_),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_4 fanout91 (.A(_0999_),
    .X(net91));
 sky130_fd_sc_hd__buf_4 fanout92 (.A(net93),
    .X(net92));
 sky130_fd_sc_hd__buf_4 fanout93 (.A(_0998_),
    .X(net93));
 sky130_fd_sc_hd__buf_4 fanout94 (.A(_0998_),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_4 fanout95 (.A(_0998_),
    .X(net95));
 sky130_fd_sc_hd__buf_6 fanout96 (.A(_0993_),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_8 fanout97 (.A(net99),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_4 fanout98 (.A(net99),
    .X(net98));
 sky130_fd_sc_hd__buf_6 fanout99 (.A(_1463_),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\RAM[49][4] ),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0218_),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_0525_),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_2 hold1000 (.A(\mem_cycle[3] ),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1001 (.A(_0045_),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1002 (.A(\ROM_addr_buff[8] ),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1003 (.A(_0505_),
    .X(net1181));
 sky130_fd_sc_hd__buf_2 hold1004 (.A(\mem_cycle[0] ),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1005 (.A(_0042_),
    .X(net1183));
 sky130_fd_sc_hd__clkbuf_2 hold1006 (.A(\insin[4] ),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1007 (.A(_0016_),
    .X(net1185));
 sky130_fd_sc_hd__buf_1 hold1008 (.A(\P[5] ),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1009 (.A(_0011_),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\RAM[34][4] ),
    .X(net279));
 sky130_fd_sc_hd__buf_2 hold1010 (.A(\mem_cycle[1] ),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1011 (.A(_1060_),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1012 (.A(_0043_),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1013 (.A(ROM_OEB),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1014 (.A(_1546_),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1015 (.A(\ROM_addr_buff[9] ),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1016 (.A(_0506_),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1017 (.A(\mem_cycle[1] ),
    .X(net1195));
 sky130_fd_sc_hd__buf_1 hold1018 (.A(_0574_),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1019 (.A(\P[1] ),
    .X(net1197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_0272_),
    .X(net280));
 sky130_fd_sc_hd__buf_1 hold1020 (.A(net34),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1021 (.A(net61),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1022 (.A(_0005_),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1023 (.A(net50),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1024 (.A(_0111_),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1025 (.A(net68),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1026 (.A(_1533_),
    .X(net1204));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1027 (.A(\mem_cycle[2] ),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1028 (.A(_1061_),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1029 (.A(_0044_),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\RAM[40][1] ),
    .X(net281));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold1030 (.A(\startup_cycle[5] ),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1031 (.A(_1504_),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1032 (.A(_0481_),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1033 (.A(\MAR[3] ),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1034 (.A(net48),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1035 (.A(net52),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1036 (.A(_0112_),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1037 (.A(net47),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1038 (.A(\MAR[1] ),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1039 (.A(_0001_),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_0189_),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1040 (.A(net64),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1041 (.A(_1126_),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1042 (.A(_0125_),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1043 (.A(net49),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1044 (.A(_0110_),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1045 (.A(\insin[0] ),
    .X(net1223));
 sky130_fd_sc_hd__buf_1 hold1046 (.A(\ROM_spi_cycle[4] ),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1047 (.A(_0475_),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1048 (.A(\insin[1] ),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1049 (.A(net46),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\RAM[6][5] ),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1050 (.A(net40),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1051 (.A(_1394_),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1052 (.A(_0413_),
    .X(net1230));
 sky130_fd_sc_hd__buf_1 hold1053 (.A(\ROM_spi_cycle[1] ),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1054 (.A(_1488_),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1055 (.A(_0472_),
    .X(net1233));
 sky130_fd_sc_hd__buf_1 hold1056 (.A(\startup_cycle[3] ),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1057 (.A(_0479_),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1058 (.A(net32),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1059 (.A(_1450_),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_0223_),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1060 (.A(\ROM_spi_cycle[0] ),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1061 (.A(\insin[3] ),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1062 (.A(\MAR[0] ),
    .X(net1240));
 sky130_fd_sc_hd__buf_1 hold1063 (.A(\P[4] ),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1064 (.A(\mem_cycle[2] ),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1065 (.A(\P[3] ),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1066 (.A(_1448_),
    .X(net1244));
 sky130_fd_sc_hd__buf_1 hold1067 (.A(net31),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1068 (.A(_1443_),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1069 (.A(\P[0] ),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\RAM[16][2] ),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1070 (.A(\P[2] ),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1071 (.A(\MAR[4] ),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1072 (.A(\B[1] ),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1073 (.A(\B[0] ),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1074 (.A(\PC[2] ),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1075 (.A(\PC[0] ),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1076 (.A(\B[3] ),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1077 (.A(\B[5] ),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1078 (.A(\B[4] ),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1079 (.A(\PC[5] ),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_0354_),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1080 (.A(\PC[3] ),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1081 (.A(\B[2] ),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1082 (.A(\PC[6] ),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1083 (.A(\PC[1] ),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1084 (.A(\PC[4] ),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1085 (.A(net31),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1086 (.A(\A[3] ),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1087 (.A(\instr_cycle[1] ),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\RAM[12][3] ),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\RAM[0][4] ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_0307_),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\RAM[2][1] ),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_0335_),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\RAM[25][2] ),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_0390_),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\RAM[56][3] ),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_0155_),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\RAM[40][4] ),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_0192_),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\RAM[32][2] ),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0266_),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_0300_),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\RAM[0][3] ),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_0265_),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\RAM[4][1] ),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_0523_),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\RAM[9][1] ),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(_0535_),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\RAM[23][0] ),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(_0182_),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\RAM[20][1] ),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\RAM[32][3] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_0096_),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\RAM[48][0] ),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_0119_),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\RAM[56][2] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(_0154_),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\RAM[20][3] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_0098_),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\RAM[10][1] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_0275_),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\RAM[36][3] ),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0301_),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(_0239_),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\RAM[12][1] ),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_0305_),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\RAM[24][0] ),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_0194_),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\RAM[52][0] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_0047_),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\RAM[20][4] ),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_0099_),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\RAM[34][1] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\RAM[33][5] ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(_0269_),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\RAM[18][4] ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_0380_),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\RAM[1][1] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(_0395_),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\RAM[16][1] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_0353_),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\RAM[24][5] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_0199_),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\RAM[33][0] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_0291_),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(_0286_),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\RAM[54][2] ),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_0073_),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\RAM[1][4] ),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_0398_),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\RAM[50][1] ),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_0025_),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\RAM[4][2] ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(_0524_),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\RAM[40][0] ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\RAM[5][0] ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_0188_),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\RAM[36][2] ),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_0238_),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\RAM[2][4] ),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(_0338_),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\RAM[52][2] ),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(_0049_),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\RAM[54][4] ),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_0075_),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\RAM[13][1] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_0280_),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(_0317_),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\RAM[10][2] ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(_0276_),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\RAM[12][0] ),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(_0304_),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\RAM[20][0] ),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(_0095_),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\RAM[44][3] ),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(_0531_),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\RAM[45][3] ),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\RAM[32][0] ),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(_0033_),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\RAM[2][2] ),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(_0336_),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\RAM[0][0] ),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(_0262_),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\RAM[54][0] ),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(_0071_),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\RAM[56][0] ),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(_0152_),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\last_PC[6] ),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0093_),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_0298_),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(_0437_),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\RAM[32][1] ),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_0299_),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\RAM[1][2] ),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(_0396_),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\RAM[36][1] ),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(_0237_),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\RAM[52][4] ),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_0051_),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\RAM[17][4] ),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\RAM[49][3] ),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_0368_),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\RAM[34][2] ),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(_0270_),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\RAM[33][2] ),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(_0288_),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\RAM[1][5] ),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(_0399_),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\RAM[40][5] ),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(_0193_),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\RAM[32][4] ),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0092_),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(_0302_),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\RAM[13][4] ),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(_0320_),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\RAM[13][3] ),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(_0319_),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\RAM[61][0] ),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(_0248_),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\RAM[14][0] ),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(_0328_),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\RAM[44][1] ),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\RAM[52][1] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(_0529_),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\RAM[7][2] ),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_0232_),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\RAM[7][1] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(_0231_),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\RAM[12][2] ),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(_0306_),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\RAM[1][0] ),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(_0394_),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\last_P[0] ),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_0048_),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(_0463_),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\RAM[52][3] ),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(_0050_),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\RAM[12][4] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(_0308_),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\RAM[5][2] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(_0282_),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\RAM[26][2] ),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(_0372_),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\last_PC[0] ),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\RAM[50][5] ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(_0431_),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\RAM[7][5] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(_0235_),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\RAM[8][3] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(_0245_),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\RAM[34][0] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(_0268_),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\RAM[29][2] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(_0067_),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\RAM[15][0] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_0029_),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(_0340_),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\RAM[17][2] ),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(_0366_),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\RAM[49][0] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(_0089_),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\RAM[33][3] ),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(_0289_),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\RAM[7][0] ),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(_0230_),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\RAM[9][0] ),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\RAM[17][3] ),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(_0534_),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\RAM[2][5] ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(_0339_),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\RAM[5][4] ),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(_0284_),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\RAM[35][3] ),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(_0259_),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\RAM[24][3] ),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_0197_),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\RAM[54][1] ),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0367_),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(_0072_),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\RAM[37][0] ),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(_0224_),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\RAM[0][5] ),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(_0267_),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\last_P[3] ),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(_0466_),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\RAM[0][2] ),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(_0264_),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\RAM[5][5] ),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\RAM[8][5] ),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(_0285_),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\RAM[47][3] ),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(_0149_),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\RAM[42][5] ),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(_0169_),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\RAM[10][4] ),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(_0278_),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\last_PC[7] ),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(_0438_),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\RAM[18][5] ),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\RAM[52][5] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0247_),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(_0381_),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\RAM[25][5] ),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(_0393_),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\RAM[25][3] ),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(_0391_),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\RAM[46][3] ),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(_0131_),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\RAM[36][0] ),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(_0236_),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\RAM[24][4] ),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\RAM[4][0] ),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(_0198_),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\RAM[50][4] ),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(_0028_),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\last_PC[8] ),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(_0439_),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\RAM[6][3] ),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(_0221_),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\RAM[24][1] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(_0195_),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\RAM[54][5] ),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0522_),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(_0076_),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\RAM[32][5] ),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(_0303_),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\RAM[47][1] ),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(_0147_),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\RAM[10][5] ),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(_0279_),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\last_B[2] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(_0453_),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\RAM[61][4] ),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\RAM[6][1] ),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(_0252_),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\RAM[43][2] ),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(_0103_),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\RAM[37][1] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(_0225_),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\last_B[4] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(_0455_),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\RAM[62][1] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(_0383_),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\RAM[39][4] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0219_),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(_0081_),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\RAM[30][4] ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(_0326_),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\RAM[9][5] ),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(_0539_),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\RAM[3][4] ),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(_0204_),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\RAM[3][1] ),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(_0201_),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\last_PC[11] ),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\RAM[6][4] ),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(_0442_),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\RAM[57][1] ),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(_0114_),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\RAM[36][5] ),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(_0241_),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\RAM[23][4] ),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(_0186_),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\RAM[62][2] ),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(_0384_),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\RAM[45][1] ),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_0222_),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(_0031_),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\RAM[30][2] ),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(_0324_),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\RAM[42][2] ),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(_0166_),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\RAM[51][1] ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(_0037_),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\RAM[17][5] ),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(_0369_),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\RAM[25][1] ),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\RAM[56][1] ),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(_0389_),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\RAM[14][1] ),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(_0329_),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\RAM[41][4] ),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(_0180_),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\last_P[5] ),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(_0468_),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\RAM[39][1] ),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(_0078_),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\RAM[51][4] ),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_0153_),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(_0040_),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\RAM[8][0] ),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(_0242_),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\RAM[62][4] ),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(_0386_),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\last_P[2] ),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(_0465_),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\RAM[1][3] ),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(_0397_),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\last_PC[4] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\last_PC[1] ),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(_0435_),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\RAM[50][0] ),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(_0024_),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\RAM[25][4] ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(_0392_),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\RAM[15][1] ),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(_0341_),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\RAM[62][5] ),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(_0387_),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\RAM[41][1] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0052_),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_0432_),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(_0177_),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\RAM[45][0] ),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(_0030_),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\RAM[54][3] ),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(_0074_),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\RAM[43][5] ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(_0106_),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\last_A[0] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(_0445_),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\last_PC[9] ),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\RAM[48][5] ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(_0440_),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\RAM[46][4] ),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(_0132_),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\RAM[20][2] ),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(_0097_),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\RAM[46][1] ),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(_0129_),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\last_MAR[4] ),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(_0461_),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\RAM[18][2] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0124_),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(_0378_),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\RAM[9][3] ),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(_0537_),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\imm_buff[0] ),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(_0427_),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\RAM[12][5] ),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(_0309_),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\RAM[31][3] ),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(_0313_),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\RAM[13][5] ),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\RAM[2][3] ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(_0321_),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\RAM[28][5] ),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(_0351_),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\RAM[25][0] ),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(_0388_),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\last_MAR[3] ),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(_0460_),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\RAM[57][0] ),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(_0113_),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\RAM[11][3] ),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_0337_),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(_0295_),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\RAM[61][3] ),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(_0251_),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\RAM[30][5] ),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(_0327_),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\RAM[13][0] ),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(_0316_),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\last_PC[10] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(_0441_),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\RAM[61][1] ),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\RAM[49][2] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(_0249_),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\RAM[62][0] ),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(_0382_),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\RAM[31][4] ),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(_0314_),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\RAM[62][3] ),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(_0385_),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\RAM[53][4] ),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(_0063_),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\RAM[29][0] ),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_0091_),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(_0065_),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\RAM[19][2] ),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(_0055_),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\RAM[21][1] ),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(_0159_),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\RAM[28][1] ),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(_0347_),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\RAM[51][5] ),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(_0041_),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\RAM[22][4] ),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\RAM[16][0] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(_0174_),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\RAM[36][4] ),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(_0240_),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\last_MAR[5] ),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(_0462_),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\RAM[22][2] ),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(_0172_),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\RAM[22][5] ),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(_0175_),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\RAM[43][4] ),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_0352_),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(_0105_),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\RAM[35][2] ),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(_0258_),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\RAM[28][3] ),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(_0349_),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\RAM[34][3] ),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(_0271_),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\RAM[35][4] ),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(_0260_),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\last_MAR[1] ),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\RAM[18][0] ),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(_0458_),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\RAM[16][3] ),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(_0355_),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\RAM[47][4] ),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(_0150_),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\RAM[19][5] ),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(_0058_),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\last_PC[5] ),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(_0436_),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\RAM[39][2] ),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\RAM[6][2] ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_0376_),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(_0079_),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\RAM[21][5] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(_0163_),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\RAM[57][2] ),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(_0115_),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\RAM[28][2] ),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(_0348_),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\RAM[30][3] ),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(_0325_),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\RAM[21][4] ),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\RAM[48][2] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(_0162_),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\RAM[26][5] ),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(_0375_),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\RAM[39][3] ),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(_0080_),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\RAM[0][1] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(_0263_),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\RAM[39][0] ),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(_0077_),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\last_MAR[0] ),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_0121_),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(_0457_),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\RAM[5][3] ),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(_0283_),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\RAM[44][5] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(_0533_),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\RAM[10][0] ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(_0274_),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\RAM[44][2] ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(_0530_),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\RAM[34][5] ),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\RAM[8][1] ),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(_0273_),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\RAM[7][4] ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(_0234_),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\RAM[15][3] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(_0343_),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\RAM[19][4] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(_0057_),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\RAM[41][0] ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(_0176_),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\RAM[19][3] ),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_0243_),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(_0056_),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\RAM[44][0] ),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(_0528_),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\RAM[55][2] ),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(_0085_),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\RAM[22][3] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(_0173_),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\RAM[13][2] ),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(_0318_),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(\RAM[38][4] ),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\RAM[48][1] ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(_0216_),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\RAM[55][1] ),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(_0084_),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(\RAM[29][1] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(_0066_),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(\RAM[29][4] ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(_0069_),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\RAM[15][4] ),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(_0344_),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(\RAM[55][5] ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_0120_),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(_0088_),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\RAM[27][5] ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(_0363_),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(\RAM[42][4] ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(_0168_),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\last_A[4] ),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(_0449_),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\RAM[29][5] ),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(_0070_),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\last_A[3] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\RAM[56][5] ),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(_0448_),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\last_PC[3] ),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(_0434_),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\RAM[3][5] ),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(_0205_),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\RAM[38][0] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(_0212_),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\RAM[57][4] ),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(_0117_),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\RAM[17][1] ),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_0157_),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(_0365_),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\RAM[27][4] ),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(_0362_),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\last_A[1] ),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(_0446_),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\RAM[23][2] ),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(_0184_),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\RAM[7][3] ),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(_0233_),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(\last_MAR[2] ),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\RAM[4][5] ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(_0459_),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(\RAM[55][0] ),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(_0083_),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(\RAM[9][4] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(_0538_),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\last_PC[2] ),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(_0433_),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(\RAM[35][0] ),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(_0256_),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\RAM[26][4] ),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0220_),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_0527_),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(_0374_),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\RAM[19][0] ),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(_0053_),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\RAM[35][1] ),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(_0257_),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\RAM[18][3] ),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(_0379_),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\last_B[3] ),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(_0454_),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(\RAM[45][5] ),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\RAM[8][4] ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(_0035_),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\RAM[15][2] ),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(_0342_),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\RAM[15][5] ),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(_0345_),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\RAM[37][5] ),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(_0229_),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\imm_buff[1] ),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(_0428_),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\RAM[18][1] ),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_0246_),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(_0377_),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\last_B[0] ),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(_0451_),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\RAM[46][0] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(_0128_),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\RAM[23][1] ),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(_0183_),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\RAM[31][2] ),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(_0312_),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\RAM[3][3] ),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\RAM[17][0] ),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(_0203_),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\RAM[26][0] ),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(_0370_),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\RAM[57][5] ),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(_0118_),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(\RAM[21][3] ),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(_0161_),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\RAM[38][3] ),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(_0215_),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\RAM[22][1] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_0364_),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(_0171_),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\RAM[11][0] ),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(_0292_),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\RAM[31][1] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(_0311_),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\RAM[43][3] ),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(_0104_),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\last_B[1] ),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(_0452_),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\RAM[40][2] ),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\RAM[49][5] ),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(_0190_),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\RAM[11][2] ),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(_0294_),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(\RAM[41][2] ),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(_0178_),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\RAM[23][5] ),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(_0187_),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\RAM[29][3] ),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(_0068_),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(\RAM[57][3] ),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_0094_),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(_0116_),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(\RAM[26][3] ),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(_0373_),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\RAM[35][5] ),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(_0261_),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(\RAM[47][0] ),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(_0146_),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(\RAM[20][5] ),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(_0100_),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(\RAM[11][5] ),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\RAM[33][1] ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(_0297_),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(\RAM[28][0] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(_0346_),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(\RAM[51][0] ),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(_0036_),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(\RAM[47][5] ),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(_0151_),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(\RAM[9][2] ),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(_0536_),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(\RAM[43][1] ),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_0287_),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(_0102_),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(\RAM[61][2] ),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(_0250_),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(\RAM[28][4] ),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(_0350_),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(\RAM[51][2] ),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(_0038_),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(\RAM[61][5] ),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(_0253_),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(\RAM[39][5] ),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\RAM[8][2] ),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(_0082_),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(\RAM[44][4] ),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(_0532_),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(\RAM[37][2] ),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(_0226_),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(\RAM[41][3] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(_0179_),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(\RAM[53][1] ),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(_0060_),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(\RAM[55][4] ),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\RAM[16][4] ),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_0244_),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(_0087_),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(\RAM[31][5] ),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(_0315_),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(\RAM[27][1] ),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(_0359_),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(\RAM[51][3] ),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(_0039_),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(\last_A[2] ),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(_0447_),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(\RAM[23][3] ),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\RAM[16][5] ),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(_0185_),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(\RAM[27][3] ),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(_0361_),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(\RAM[31][0] ),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(_0310_),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(\RAM[30][1] ),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(_0323_),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(\RAM[38][2] ),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(_0214_),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(\RAM[38][5] ),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_0357_),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(_0217_),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(\RAM[41][5] ),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(_0181_),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(\RAM[30][0] ),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(_0322_),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(\RAM[45][2] ),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(_0032_),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(\RAM[11][1] ),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(_0293_),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(\RAM[11][4] ),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\RAM[48][3] ),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(_0296_),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(\RAM[27][2] ),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(_0360_),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(\RAM[40][3] ),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(_0191_),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(\RAM[21][2] ),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(_0160_),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(\RAM[37][3] ),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(_0227_),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(\RAM[19][1] ),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_0122_),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(_0054_),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(\RAM[3][0] ),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(_0200_),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(\RAM[46][5] ),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(_0133_),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(\RAM[46][2] ),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(_0130_),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(\RAM[21][0] ),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(_0158_),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(\RAM[53][3] ),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\RAM[49][1] ),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(_0062_),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(\RAM[42][0] ),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(_0164_),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(\RAM[42][1] ),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(_0165_),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(\RAM[43][0] ),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(_0101_),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(\RAM[14][5] ),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(_0333_),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(\last_A[5] ),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_0090_),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(_0450_),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(\RAM[3][2] ),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(_0202_),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(\RAM[45][4] ),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(_0034_),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(\RAM[53][2] ),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(_0061_),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(\last_P[4] ),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(_0467_),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(\RAM[14][2] ),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\RAM[10][3] ),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(_0330_),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(\RAM[55][3] ),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(_0086_),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(\RAM[22][0] ),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(_0170_),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(\RAM[53][5] ),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(_0064_),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(\RAM[47][2] ),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(_0148_),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(\RAM[27][0] ),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_0277_),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(_0358_),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(\RAM[38][1] ),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(_0213_),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(\RAM[59][0] ),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(_0134_),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(\ROM_spi_dat_out[0] ),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(_1551_),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(\RAM[53][0] ),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(_0059_),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(\RAM[42][3] ),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\last_B[5] ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(_0167_),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(\RAM[14][4] ),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(_0332_),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(\last_flags[0] ),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(_0443_),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(\RAM[26][1] ),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(_0371_),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(\RAM[14][3] ),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(_0331_),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(\RAM[37][4] ),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0356_),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_0456_),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(_0228_),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(needs_irupt),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(_0469_),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(\ROM_spi_dat_out[1] ),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(_0490_),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(\last_P[1] ),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(_0464_),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(ROM_spi_mode),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(_1547_),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(\ROM_spi_dat_out[5] ),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\RAM[4][4] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(_0494_),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(\ROM_spi_dat_out[6] ),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(_0495_),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(\ROM_spi_dat_out[7] ),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(_0496_),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(\imm_buff[2] ),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(_0429_),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(\ROM_spi_dat_out[3] ),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(_0492_),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(\last_flags[1] ),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0526_),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(_0444_),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(\ROM_spi_dat_out[4] ),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(_0493_),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(\imm_buff[4] ),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(_0254_),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(\ROM_spi_dat_out[2] ),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(_0491_),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(\imm_buff[3] ),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(_0430_),
    .X(net1006));
 sky130_fd_sc_hd__buf_2 hold829 (.A(\startup_cycle[1] ),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\RAM[24][2] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(_0477_),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(spi_clkdiv),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(_1595_),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(\imm_buff[5] ),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(_0255_),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(\ROM_dest[1] ),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(_0626_),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(_0019_),
    .X(net1015));
 sky130_fd_sc_hd__clkbuf_2 hold838 (.A(\ROM_addr_buff[10] ),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(_0519_),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0196_),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(net65),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(_0126_),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(net66),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(_0127_),
    .X(net1021));
 sky130_fd_sc_hd__buf_1 hold844 (.A(\PC[3] ),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(_0417_),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(net67),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(_0484_),
    .X(net1025));
 sky130_fd_sc_hd__buf_1 hold848 (.A(\PC[2] ),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(_0416_),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\RAM[50][3] ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(\B[2] ),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(_0408_),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(\B[4] ),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(_0410_),
    .X(net1031));
 sky130_fd_sc_hd__buf_1 hold854 (.A(\PC[5] ),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(_0419_),
    .X(net1033));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold856 (.A(\ROM_dest[0] ),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(_0018_),
    .X(net1035));
 sky130_fd_sc_hd__buf_1 hold858 (.A(\ROM_addr_buff[5] ),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(_0502_),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_0027_),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_2 hold860 (.A(net54),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(_1459_),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(_0426_),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(\last_addr[3] ),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(_1586_),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(_0512_),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(\last_addr[9] ),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(_1592_),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(_0518_),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(\last_addr[5] ),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\RAM[56][4] ),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(_1588_),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(_0514_),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(\last_addr[6] ),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(_1589_),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(_0515_),
    .X(net1052));
 sky130_fd_sc_hd__clkbuf_2 hold875 (.A(\PC[0] ),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(_0414_),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(\last_addr[2] ),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(_1585_),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(_0511_),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(_0156_),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(\RAM[59][2] ),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(net43),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(_0209_),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(\RAM[59][3] ),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(_1141_),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(\last_addr[8] ),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(_1591_),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(_0517_),
    .X(net1065));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold888 (.A(net33),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(_1579_),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\RAM[48][4] ),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(_0507_),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(\RAM[59][1] ),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(_1139_),
    .X(net1070));
 sky130_fd_sc_hd__clkbuf_2 hold893 (.A(\A[3] ),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(_0403_),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(\RAM[59][4] ),
    .X(net1073));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold896 (.A(\ROM_addr_buff[7] ),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(_0516_),
    .X(net1075));
 sky130_fd_sc_hd__buf_1 hold898 (.A(\ROM_addr_buff[0] ),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(_0497_),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\RAM[6][0] ),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_0123_),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(\RAM[59][5] ),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(_1143_),
    .X(net1079));
 sky130_fd_sc_hd__clkbuf_2 hold902 (.A(\insin[5] ),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(_0017_),
    .X(net1081));
 sky130_fd_sc_hd__clkbuf_2 hold904 (.A(\A[4] ),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(_0404_),
    .X(net1083));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold906 (.A(\PC[6] ),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(_0420_),
    .X(net1085));
 sky130_fd_sc_hd__buf_2 hold908 (.A(\A[0] ),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(_0400_),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\RAM[50][2] ),
    .X(net269));
 sky130_fd_sc_hd__buf_2 hold910 (.A(\startup_cycle[4] ),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(_0480_),
    .X(net1089));
 sky130_fd_sc_hd__clkbuf_2 hold912 (.A(\startup_cycle[6] ),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(_0482_),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(\ROM_addr_buff[6] ),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(_0503_),
    .X(net1093));
 sky130_fd_sc_hd__clkbuf_2 hold916 (.A(\ROM_dest[2] ),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(_0020_),
    .X(net1095));
 sky130_fd_sc_hd__clkbuf_2 hold918 (.A(\A[1] ),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(_0401_),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_0026_),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(\ROM_spi_cycle[2] ),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(_1489_),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(_0473_),
    .X(net1100));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold923 (.A(\A[2] ),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(_0402_),
    .X(net1102));
 sky130_fd_sc_hd__buf_1 hold925 (.A(\B[5] ),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(_0411_),
    .X(net1104));
 sky130_fd_sc_hd__buf_1 hold927 (.A(\ROM_addr_buff[4] ),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(_0513_),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(\ROM_spi_cycle[3] ),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\RAM[2][0] ),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(_1492_),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(_0474_),
    .X(net1109));
 sky130_fd_sc_hd__clkbuf_2 hold932 (.A(net1266),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(_0022_),
    .X(net1111));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold934 (.A(\A[5] ),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(_0405_),
    .X(net1113));
 sky130_fd_sc_hd__buf_1 hold936 (.A(\ROM_addr_buff[1] ),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(_0510_),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(net62),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(_1465_),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_0334_),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(_0470_),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(net69),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(_0206_),
    .X(net1120));
 sky130_fd_sc_hd__buf_1 hold943 (.A(\B[1] ),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(_0407_),
    .X(net1122));
 sky130_fd_sc_hd__clkbuf_2 hold945 (.A(\startup_cycle[2] ),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(_1499_),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(_0478_),
    .X(net1125));
 sky130_fd_sc_hd__buf_1 hold948 (.A(\ROM_addr_buff[11] ),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(_0520_),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\RAM[33][4] ),
    .X(net273));
 sky130_fd_sc_hd__buf_1 hold950 (.A(\B[3] ),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(_0409_),
    .X(net1129));
 sky130_fd_sc_hd__buf_1 hold952 (.A(\PC[1] ),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(_1570_),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(_0498_),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(net45),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(net58),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(\ROM_addr_buff[2] ),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(_0499_),
    .X(net1136));
 sky130_fd_sc_hd__buf_1 hold959 (.A(\PC[4] ),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_0290_),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(_1573_),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(_0501_),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(net59),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(\last_addr[0] ),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(_1583_),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(_0509_),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold966 (.A(\ROM_addr_buff[3] ),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(_0500_),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(net41),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(net63),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\RAM[5][1] ),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(_1541_),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(net44),
    .X(net1149));
 sky130_fd_sc_hd__clkbuf_2 hold972 (.A(\insin[3] ),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(_0976_),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(_0015_),
    .X(net1152));
 sky130_fd_sc_hd__buf_1 hold975 (.A(net30),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold976 (.A(_1576_),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold977 (.A(_0504_),
    .X(net1155));
 sky130_fd_sc_hd__buf_1 hold978 (.A(\B[0] ),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold979 (.A(_0406_),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_0281_),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold980 (.A(net42),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold981 (.A(net57),
    .X(net1159));
 sky130_fd_sc_hd__clkbuf_2 hold982 (.A(\insin[2] ),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold983 (.A(_0975_),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold984 (.A(_0014_),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold985 (.A(net55),
    .X(net1163));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold986 (.A(\startup_cycle[0] ),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold987 (.A(_0476_),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold988 (.A(\instr_cycle[2] ),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold989 (.A(_1411_),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\RAM[4][3] ),
    .X(net277));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold990 (.A(\mem_cycle[4] ),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold991 (.A(_0046_),
    .X(net1169));
 sky130_fd_sc_hd__clkbuf_4 hold992 (.A(net53),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold993 (.A(_1438_),
    .X(net1171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold994 (.A(net56),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold995 (.A(net60),
    .X(net1173));
 sky130_fd_sc_hd__buf_1 hold996 (.A(net51),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold997 (.A(_1399_),
    .X(net1175));
 sky130_fd_sc_hd__buf_1 hold998 (.A(_1401_),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold999 (.A(_0418_),
    .X(net1177));
 sky130_fd_sc_hd__buf_1 input1 (.A(io_in[10]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(io_in[19]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(io_in[20]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(io_in[29]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(io_in[3]),
    .X(net13));
 sky130_fd_sc_hd__buf_4 input14 (.A(io_in[4]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input15 (.A(io_in[5]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input16 (.A(io_in[6]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(io_in[9]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(rst_n),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input2 (.A(io_in[11]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(io_in[12]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(io_in[13]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(io_in[14]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(io_in[15]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(io_in[16]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(io_in[17]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(io_in[18]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 max_cap1 (.A(_1083_),
    .X(net1265));
 sky130_fd_sc_hd__buf_4 max_cap100 (.A(_0992_),
    .X(net100));
 sky130_fd_sc_hd__buf_4 max_cap101 (.A(_0992_),
    .X(net101));
 sky130_fd_sc_hd__buf_12 output19 (.A(net19),
    .X(io_oeb[10]));
 sky130_fd_sc_hd__buf_12 output20 (.A(net20),
    .X(io_oeb[11]));
 sky130_fd_sc_hd__buf_12 output21 (.A(net21),
    .X(io_oeb[12]));
 sky130_fd_sc_hd__buf_12 output22 (.A(net22),
    .X(io_oeb[13]));
 sky130_fd_sc_hd__buf_12 output23 (.A(net23),
    .X(io_oeb[14]));
 sky130_fd_sc_hd__buf_12 output24 (.A(net24),
    .X(io_oeb[15]));
 sky130_fd_sc_hd__buf_12 output25 (.A(net25),
    .X(io_oeb[16]));
 sky130_fd_sc_hd__buf_12 output26 (.A(net26),
    .X(io_oeb[17]));
 sky130_fd_sc_hd__buf_12 output27 (.A(net27),
    .X(io_oeb[18]));
 sky130_fd_sc_hd__buf_12 output28 (.A(net28),
    .X(io_oeb[19]));
 sky130_fd_sc_hd__buf_12 output29 (.A(net29),
    .X(io_oeb[20]));
 sky130_fd_sc_hd__buf_12 output30 (.A(net30),
    .X(io_oeb[31]));
 sky130_fd_sc_hd__buf_12 output31 (.A(net31),
    .X(io_oeb[32]));
 sky130_fd_sc_hd__buf_12 output32 (.A(net32),
    .X(io_oeb[33]));
 sky130_fd_sc_hd__buf_12 output33 (.A(net33),
    .X(io_oeb[34]));
 sky130_fd_sc_hd__buf_12 output34 (.A(net34),
    .X(io_oeb[35]));
 sky130_fd_sc_hd__buf_12 output35 (.A(net35),
    .X(io_oeb[3]));
 sky130_fd_sc_hd__buf_12 output36 (.A(net36),
    .X(io_oeb[4]));
 sky130_fd_sc_hd__buf_12 output37 (.A(net37),
    .X(io_oeb[5]));
 sky130_fd_sc_hd__buf_12 output38 (.A(net38),
    .X(io_oeb[6]));
 sky130_fd_sc_hd__buf_12 output39 (.A(net39),
    .X(io_oeb[9]));
 sky130_fd_sc_hd__buf_12 output40 (.A(net40),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_12 output41 (.A(net41),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_12 output42 (.A(net42),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_12 output43 (.A(net43),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_12 output44 (.A(net44),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_12 output45 (.A(net45),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_12 output46 (.A(net46),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_12 output47 (.A(net47),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_12 output48 (.A(net48),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_12 output49 (.A(net49),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_12 output50 (.A(net50),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_12 output51 (.A(net51),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_12 output52 (.A(net52),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_12 output53 (.A(net53),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_12 output54 (.A(net54),
    .X(io_out[22]));
 sky130_fd_sc_hd__buf_12 output55 (.A(net55),
    .X(io_out[23]));
 sky130_fd_sc_hd__buf_12 output56 (.A(net56),
    .X(io_out[24]));
 sky130_fd_sc_hd__buf_12 output57 (.A(net57),
    .X(io_out[25]));
 sky130_fd_sc_hd__buf_12 output58 (.A(net58),
    .X(io_out[26]));
 sky130_fd_sc_hd__buf_12 output59 (.A(net59),
    .X(io_out[27]));
 sky130_fd_sc_hd__buf_12 output60 (.A(net60),
    .X(io_out[28]));
 sky130_fd_sc_hd__buf_12 output61 (.A(net116),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_12 output62 (.A(net62),
    .X(io_out[30]));
 sky130_fd_sc_hd__buf_12 output63 (.A(net63),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_12 output64 (.A(net64),
    .X(io_out[4]));
 sky130_fd_sc_hd__buf_12 output65 (.A(net65),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_12 output66 (.A(net66),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_12 output67 (.A(net67),
    .X(io_out[7]));
 sky130_fd_sc_hd__buf_12 output68 (.A(net68),
    .X(io_out[8]));
 sky130_fd_sc_hd__buf_12 output69 (.A(net69),
    .X(io_out[9]));
 sky130_fd_sc_hd__conb_1 scrapcpu_158 (.LO(net158));
 sky130_fd_sc_hd__conb_1 scrapcpu_159 (.LO(net159));
 sky130_fd_sc_hd__conb_1 scrapcpu_160 (.LO(net160));
 sky130_fd_sc_hd__conb_1 scrapcpu_161 (.LO(net161));
 sky130_fd_sc_hd__conb_1 scrapcpu_162 (.LO(net162));
 sky130_fd_sc_hd__conb_1 scrapcpu_163 (.LO(net163));
 sky130_fd_sc_hd__conb_1 scrapcpu_164 (.LO(net164));
 sky130_fd_sc_hd__conb_1 scrapcpu_165 (.LO(net165));
 sky130_fd_sc_hd__conb_1 scrapcpu_166 (.LO(net166));
 sky130_fd_sc_hd__conb_1 scrapcpu_167 (.LO(net167));
 sky130_fd_sc_hd__conb_1 scrapcpu_168 (.LO(net168));
 sky130_fd_sc_hd__conb_1 scrapcpu_169 (.LO(net169));
 sky130_fd_sc_hd__conb_1 scrapcpu_170 (.LO(net170));
 sky130_fd_sc_hd__conb_1 scrapcpu_171 (.LO(net171));
 sky130_fd_sc_hd__conb_1 scrapcpu_172 (.LO(net172));
 sky130_fd_sc_hd__conb_1 scrapcpu_173 (.LO(net173));
 sky130_fd_sc_hd__conb_1 scrapcpu_174 (.LO(net174));
 sky130_fd_sc_hd__conb_1 scrapcpu_175 (.LO(net175));
 sky130_fd_sc_hd__conb_1 scrapcpu_176 (.LO(net176));
 sky130_fd_sc_hd__conb_1 scrapcpu_177 (.LO(net177));
 sky130_fd_sc_hd__conb_1 scrapcpu_178 (.HI(net178));
 sky130_fd_sc_hd__buf_1 wire109 (.A(_0564_),
    .X(net109));
 assign io_oeb[0] = net158;
 assign io_oeb[1] = net159;
 assign io_oeb[21] = net163;
 assign io_oeb[22] = net164;
 assign io_oeb[23] = net165;
 assign io_oeb[24] = net166;
 assign io_oeb[25] = net167;
 assign io_oeb[26] = net168;
 assign io_oeb[27] = net169;
 assign io_oeb[28] = net170;
 assign io_oeb[29] = net178;
 assign io_oeb[2] = net160;
 assign io_oeb[30] = net171;
 assign io_oeb[7] = net161;
 assign io_oeb[8] = net162;
 assign io_out[29] = net172;
 assign io_out[31] = net173;
 assign io_out[32] = net174;
 assign io_out[33] = net175;
 assign io_out[34] = net176;
 assign io_out[35] = net177;
endmodule

